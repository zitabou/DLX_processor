
module hardwired_CU ( clk, rst, opcode, func, RF1, RF2, EN1, S1, S2, ALU3, 
        ALU2, ALU1, ALU0, SN, LnS, Wrd, BHU1, BHU0, EN3, S3, WF1, Ld );
  input [5:0] opcode;
  input [10:0] func;
  input clk, rst;
  output RF1, RF2, EN1, S1, S2, ALU3, ALU2, ALU1, ALU0, SN, LnS, Wrd, BHU1,
         BHU0, EN3, S3, WF1, Ld;
  wire   exe_type2, exe_type21, exe_type22, exe_type23, N190, n1, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n142, n143, n144, n145, n146;
  wire   [5:0] cw2;
  wire   [1:0] cw3;
  wire   [6:0] cw21;
  wire   [6:0] cw22;
  wire   [6:0] cw23;
  wire   [13:0] cw1;

  DFFR_X1 \cw2_reg[13]  ( .D(cw1[13]), .CK(clk), .RN(n4), .Q(S1) );
  DFFR_X1 \cw2_reg[12]  ( .D(cw1[12]), .CK(clk), .RN(n2), .Q(S2) );
  DFFR_X1 \cw2_reg[11]  ( .D(cw1[11]), .CK(clk), .RN(n2), .Q(ALU3) );
  DFFR_X1 \cw2_reg[10]  ( .D(cw1[10]), .CK(clk), .RN(n2), .Q(ALU2) );
  DFFR_X1 \cw2_reg[9]  ( .D(cw1[9]), .CK(clk), .RN(n2), .Q(ALU1) );
  DFFR_X1 \cw2_reg[8]  ( .D(cw1[8]), .CK(clk), .RN(n2), .Q(ALU0) );
  DFFR_X1 \cw2_reg[7]  ( .D(cw1[7]), .CK(clk), .RN(n2), .Q(SN) );
  DFFR_X1 \cw2_reg[6]  ( .D(cw1[6]), .CK(clk), .RN(n2), .Q(Ld) );
  DFFR_X1 \cw2_reg[5]  ( .D(cw1[5]), .CK(clk), .RN(n2), .Q(cw2[5]) );
  DFFR_X1 \cw2_reg[4]  ( .D(cw1[4]), .CK(clk), .RN(n2), .Q(cw2[4]) );
  DFFR_X1 \cw2_reg[3]  ( .D(cw1[3]), .CK(clk), .RN(n2), .Q(cw2[3]) );
  DFFR_X1 \cw2_reg[2]  ( .D(cw1[2]), .CK(clk), .RN(n3), .Q(cw2[2]) );
  DFFR_X1 \cw2_reg[1]  ( .D(cw1[1]), .CK(clk), .RN(n3), .Q(cw2[1]) );
  DFFR_X1 \cw2_reg[0]  ( .D(cw1[0]), .CK(clk), .RN(n3), .Q(cw2[0]) );
  DFFR_X1 \cw21_reg[6]  ( .D(Ld), .CK(clk), .RN(n3), .Q(cw21[6]) );
  DFFR_X1 \cw21_reg[5]  ( .D(cw2[5]), .CK(clk), .RN(n3), .Q(cw21[5]) );
  DFFR_X1 \cw21_reg[4]  ( .D(cw2[4]), .CK(clk), .RN(n3), .Q(cw21[4]) );
  DFFR_X1 \cw21_reg[3]  ( .D(cw2[3]), .CK(clk), .RN(n3), .Q(cw21[3]) );
  DFFR_X1 \cw21_reg[2]  ( .D(cw2[2]), .CK(clk), .RN(n3), .Q(cw21[2]) );
  DFFR_X1 \cw21_reg[1]  ( .D(cw2[1]), .CK(clk), .RN(n3), .Q(cw21[1]) );
  DFFR_X1 \cw21_reg[0]  ( .D(cw2[0]), .CK(clk), .RN(n3), .Q(cw21[0]) );
  DFFR_X1 \cw22_reg[6]  ( .D(cw21[6]), .CK(clk), .RN(n3), .Q(cw22[6]) );
  DFFR_X1 \cw22_reg[5]  ( .D(cw21[5]), .CK(clk), .RN(n4), .Q(cw22[5]) );
  DFFR_X1 \cw22_reg[4]  ( .D(cw21[4]), .CK(clk), .RN(n4), .Q(cw22[4]) );
  DFFR_X1 \cw22_reg[3]  ( .D(cw21[3]), .CK(clk), .RN(n4), .Q(cw22[3]) );
  DFFR_X1 \cw22_reg[2]  ( .D(cw21[2]), .CK(clk), .RN(n4), .Q(cw22[2]) );
  DFFR_X1 \cw22_reg[1]  ( .D(cw21[1]), .CK(clk), .RN(n4), .Q(cw22[1]) );
  DFFR_X1 \cw22_reg[0]  ( .D(cw21[0]), .CK(clk), .RN(n4), .Q(cw22[0]) );
  DFFR_X1 \cw23_reg[6]  ( .D(cw22[6]), .CK(clk), .RN(n4), .Q(cw23[6]) );
  DFFR_X1 \cw23_reg[5]  ( .D(cw22[5]), .CK(clk), .RN(n4), .Q(cw23[5]) );
  DFFR_X1 \cw23_reg[4]  ( .D(cw22[4]), .CK(clk), .RN(n4), .Q(cw23[4]) );
  DFFR_X1 \cw23_reg[3]  ( .D(cw22[3]), .CK(clk), .RN(n4), .Q(cw23[3]) );
  DFFR_X1 \cw23_reg[2]  ( .D(cw22[2]), .CK(clk), .RN(n5), .Q(cw23[2]) );
  DFFR_X1 \cw23_reg[1]  ( .D(cw22[1]), .CK(clk), .RN(n5), .Q(cw23[1]) );
  DFFR_X1 \cw23_reg[0]  ( .D(cw22[0]), .CK(clk), .RN(n5), .Q(cw23[0]) );
  DFFR_X1 exe_type2_reg ( .D(N190), .CK(clk), .RN(n5), .Q(exe_type2) );
  DFFR_X1 exe_type21_reg ( .D(exe_type2), .CK(clk), .RN(n5), .Q(exe_type21) );
  DFFR_X1 exe_type22_reg ( .D(exe_type21), .CK(clk), .RN(n5), .Q(exe_type22)
         );
  DFFR_X1 exe_type23_reg ( .D(exe_type22), .CK(clk), .RN(n5), .Q(exe_type23), 
        .QN(n1) );
  SDFFR_X1 \cw3_reg[6]  ( .D(cw23[6]), .SI(Ld), .SE(n1), .CK(clk), .RN(n5), 
        .Q(LnS) );
  SDFFR_X1 \cw3_reg[5]  ( .D(cw2[5]), .SI(cw23[5]), .SE(exe_type23), .CK(clk), 
        .RN(n5), .Q(Wrd) );
  SDFFR_X1 \cw3_reg[4]  ( .D(cw2[4]), .SI(cw23[4]), .SE(exe_type23), .CK(clk), 
        .RN(n5), .Q(BHU1) );
  SDFFR_X1 \cw3_reg[3]  ( .D(cw2[3]), .SI(cw23[3]), .SE(exe_type23), .CK(clk), 
        .RN(n6), .Q(BHU0) );
  SDFFR_X1 \cw3_reg[2]  ( .D(cw2[2]), .SI(cw23[2]), .SE(exe_type23), .CK(clk), 
        .RN(n6), .Q(EN3) );
  SDFFR_X1 \cw3_reg[1]  ( .D(cw2[1]), .SI(cw23[1]), .SE(exe_type23), .CK(clk), 
        .RN(n6), .Q(cw3[1]) );
  DFFR_X1 \cw4_reg[1]  ( .D(cw3[1]), .CK(clk), .RN(n5), .Q(S3) );
  SDFFR_X1 \cw3_reg[0]  ( .D(cw2[0]), .SI(cw23[0]), .SE(exe_type23), .CK(clk), 
        .RN(n6), .Q(cw3[0]) );
  DFFR_X1 \cw4_reg[0]  ( .D(cw3[0]), .CK(clk), .RN(n2), .Q(WF1) );
  NAND3_X1 U147 ( .A1(n23), .A2(n19), .A3(opcode[4]), .ZN(n52) );
  OAI33_X1 U148 ( .A1(n46), .A2(n77), .A3(n36), .B1(n78), .B2(n30), .B3(n79), 
        .ZN(n76) );
  NAND3_X1 U149 ( .A1(opcode[5]), .A2(opcode[1]), .A3(n115), .ZN(n114) );
  NAND3_X1 U150 ( .A1(n20), .A2(n13), .A3(n24), .ZN(n124) );
  NAND3_X1 U151 ( .A1(func[0]), .A2(n36), .A3(func[1]), .ZN(n119) );
  NAND3_X1 U152 ( .A1(n128), .A2(n143), .A3(func[5]), .ZN(n46) );
  NAND3_X1 U153 ( .A1(n30), .A2(n36), .A3(func[1]), .ZN(n98) );
  NAND3_X1 U154 ( .A1(func[3]), .A2(n128), .A3(func[5]), .ZN(n118) );
  NAND3_X1 U155 ( .A1(n30), .A2(n34), .A3(func[2]), .ZN(n47) );
  NAND3_X1 U156 ( .A1(n75), .A2(n48), .A3(n94), .ZN(n125) );
  NAND3_X1 U157 ( .A1(n143), .A2(n146), .A3(n128), .ZN(n78) );
  NAND3_X1 U158 ( .A1(opcode[3]), .A2(n19), .A3(opcode[1]), .ZN(n68) );
  NAND3_X1 U159 ( .A1(n22), .A2(opcode[5]), .A3(n90), .ZN(n138) );
  NAND3_X1 U160 ( .A1(n27), .A2(n19), .A3(n8), .ZN(n140) );
  NOR2_X1 U3 ( .A1(n144), .A2(n142), .ZN(n45) );
  INV_X1 U4 ( .A(n78), .ZN(n37) );
  NAND2_X1 U5 ( .A1(n37), .A2(n35), .ZN(n94) );
  INV_X1 U6 ( .A(n73), .ZN(n33) );
  INV_X1 U7 ( .A(n99), .ZN(n28) );
  OAI22_X1 U8 ( .A1(n78), .A2(n47), .B1(n45), .B2(n98), .ZN(n70) );
  NOR3_X1 U9 ( .A1(n77), .A2(n116), .A3(n36), .ZN(n74) );
  AOI21_X1 U10 ( .B1(n45), .B2(n78), .A(n119), .ZN(n127) );
  AOI21_X1 U11 ( .B1(n45), .B2(n46), .A(n47), .ZN(n42) );
  NOR3_X1 U12 ( .A1(n102), .A2(n26), .A3(n103), .ZN(cw1[4]) );
  NOR2_X1 U13 ( .A1(n118), .A2(n77), .ZN(n73) );
  NAND2_X1 U14 ( .A1(n80), .A2(n47), .ZN(n99) );
  NAND4_X1 U15 ( .A1(n117), .A2(n33), .A3(n75), .A4(n48), .ZN(n93) );
  OAI21_X1 U16 ( .B1(n97), .B2(n99), .A(n144), .ZN(n117) );
  NOR2_X1 U17 ( .A1(n100), .A2(n101), .ZN(cw1[5]) );
  INV_X1 U18 ( .A(n85), .ZN(n24) );
  INV_X1 U19 ( .A(n103), .ZN(n8) );
  INV_X1 U20 ( .A(n90), .ZN(n14) );
  INV_X1 U21 ( .A(n98), .ZN(n29) );
  INV_X1 U22 ( .A(n118), .ZN(n144) );
  INV_X1 U23 ( .A(n134), .ZN(n21) );
  INV_X1 U24 ( .A(n79), .ZN(n35) );
  INV_X1 U25 ( .A(n68), .ZN(n16) );
  INV_X1 U26 ( .A(n102), .ZN(n17) );
  INV_X1 U27 ( .A(n116), .ZN(n142) );
  AND2_X1 U28 ( .A1(n98), .A2(n119), .ZN(n80) );
  OR2_X1 U29 ( .A1(n8), .A2(n57), .ZN(n54) );
  NOR2_X1 U30 ( .A1(n97), .A2(n29), .ZN(n96) );
  INV_X1 U31 ( .A(n48), .ZN(n32) );
  NAND2_X1 U32 ( .A1(n109), .A2(n139), .ZN(EN1) );
  OAI21_X1 U33 ( .B1(n18), .B2(n137), .A(n26), .ZN(n139) );
  INV_X1 U34 ( .A(n101), .ZN(n18) );
  NAND2_X1 U35 ( .A1(n41), .A2(n135), .ZN(RF2) );
  OR3_X1 U36 ( .A1(n104), .A2(n25), .A3(n100), .ZN(n135) );
  NAND2_X1 U37 ( .A1(n109), .A2(n7), .ZN(RF1) );
  NOR2_X1 U38 ( .A1(n134), .A2(n13), .ZN(n141) );
  NOR4_X1 U39 ( .A1(n145), .A2(n143), .A3(n130), .A4(func[6]), .ZN(n129) );
  INV_X1 U40 ( .A(func[4]), .ZN(n145) );
  INV_X1 U41 ( .A(n67), .ZN(n12) );
  NOR3_X1 U42 ( .A1(func[4]), .A2(func[6]), .A3(n130), .ZN(n128) );
  AOI211_X1 U43 ( .C1(n13), .C2(n27), .A(n19), .B(n23), .ZN(n111) );
  OAI211_X1 U44 ( .C1(n81), .C2(n41), .A(n58), .B(n82), .ZN(cw1[7]) );
  NOR3_X1 U45 ( .A1(n92), .A2(n43), .A3(n93), .ZN(n81) );
  OAI22_X1 U46 ( .A1(n28), .A2(n78), .B1(n96), .B2(n46), .ZN(n92) );
  NAND4_X1 U47 ( .A1(n17), .A2(n8), .A3(n27), .A4(n26), .ZN(n41) );
  NOR2_X1 U48 ( .A1(n19), .A2(n53), .ZN(n90) );
  NAND4_X1 U49 ( .A1(n35), .A2(n129), .A3(func[0]), .A4(n146), .ZN(n75) );
  INV_X1 U50 ( .A(n110), .ZN(n9) );
  OAI211_X1 U51 ( .C1(n25), .C2(n111), .A(n14), .B(n101), .ZN(n110) );
  NOR4_X1 U52 ( .A1(n20), .A2(n27), .A3(n26), .A4(n103), .ZN(cw1[3]) );
  NAND2_X1 U53 ( .A1(func[0]), .A2(n34), .ZN(n77) );
  OAI221_X1 U54 ( .B1(n13), .B2(n68), .C1(n121), .C2(n41), .A(n122), .ZN(
        cw1[10]) );
  NOR4_X1 U55 ( .A1(n125), .A2(n70), .A3(n126), .A4(n127), .ZN(n121) );
  AOI221_X1 U56 ( .B1(n90), .B2(n22), .C1(n15), .C2(n24), .A(n123), .ZN(n122)
         );
  NOR3_X1 U57 ( .A1(n46), .A2(func[0]), .A3(n79), .ZN(n126) );
  OAI221_X1 U58 ( .B1(n112), .B2(n13), .C1(n113), .C2(n41), .A(n114), .ZN(
        cw1[11]) );
  AOI211_X1 U59 ( .C1(n142), .C2(n99), .A(n93), .B(n74), .ZN(n113) );
  OAI221_X1 U60 ( .B1(n58), .B2(n27), .C1(n59), .C2(n41), .A(n60), .ZN(cw1[8])
         );
  NOR3_X1 U61 ( .A1(n69), .A2(n44), .A3(n70), .ZN(n59) );
  AOI221_X1 U62 ( .B1(n61), .B2(n26), .C1(n15), .C2(n62), .A(n63), .ZN(n60) );
  OAI21_X1 U63 ( .B1(n80), .B2(n46), .A(n33), .ZN(n69) );
  NOR2_X1 U64 ( .A1(n23), .A2(n27), .ZN(n57) );
  NAND2_X1 U65 ( .A1(n19), .A2(n25), .ZN(n102) );
  OAI21_X1 U66 ( .B1(n111), .B2(n25), .A(n140), .ZN(n137) );
  NAND2_X1 U67 ( .A1(n13), .A2(n23), .ZN(n103) );
  NAND2_X1 U68 ( .A1(func[1]), .A2(func[2]), .ZN(n79) );
  INV_X1 U69 ( .A(func[2]), .ZN(n36) );
  NAND2_X1 U70 ( .A1(n57), .A2(n19), .ZN(n101) );
  NAND2_X1 U71 ( .A1(n85), .A2(n19), .ZN(n104) );
  AOI21_X1 U72 ( .B1(n25), .B2(n65), .A(n19), .ZN(n120) );
  OAI21_X1 U73 ( .B1(n8), .B2(n19), .A(n53), .ZN(n49) );
  INV_X1 U74 ( .A(func[0]), .ZN(n30) );
  NAND2_X1 U75 ( .A1(n115), .A2(n23), .ZN(n67) );
  INV_X1 U76 ( .A(n66), .ZN(n20) );
  INV_X1 U77 ( .A(n136), .ZN(n7) );
  NAND2_X1 U78 ( .A1(func[5]), .A2(n129), .ZN(n116) );
  OAI21_X1 U79 ( .B1(n53), .B2(n85), .A(n10), .ZN(n84) );
  INV_X1 U80 ( .A(n86), .ZN(n10) );
  INV_X1 U81 ( .A(n107), .ZN(n15) );
  NAND2_X1 U82 ( .A1(n85), .A2(n66), .ZN(n50) );
  INV_X1 U83 ( .A(func[1]), .ZN(n34) );
  INV_X1 U84 ( .A(func[5]), .ZN(n146) );
  NAND2_X1 U85 ( .A1(n71), .A2(n72), .ZN(n44) );
  AOI211_X1 U86 ( .C1(n73), .C2(func[2]), .A(n74), .B(n31), .ZN(n72) );
  AOI21_X1 U87 ( .B1(n29), .B2(n37), .A(n76), .ZN(n71) );
  INV_X1 U88 ( .A(n75), .ZN(n31) );
  INV_X1 U89 ( .A(n65), .ZN(n22) );
  INV_X1 U90 ( .A(func[3]), .ZN(n143) );
  NAND2_X1 U91 ( .A1(n94), .A2(n95), .ZN(n43) );
  OR3_X1 U92 ( .A1(n77), .A2(func[2]), .A3(n78), .ZN(n95) );
  NAND2_X1 U93 ( .A1(n75), .A2(n138), .ZN(N190) );
  NOR3_X1 U94 ( .A1(func[1]), .A2(func[2]), .A3(func[0]), .ZN(n97) );
  NAND4_X1 U95 ( .A1(func[3]), .A2(n97), .A3(n128), .A4(n146), .ZN(n48) );
  NOR4_X1 U96 ( .A1(n32), .A2(n42), .A3(n43), .A4(n44), .ZN(n40) );
  AOI221_X1 U97 ( .B1(n20), .B2(opcode[4]), .C1(opcode[2]), .C2(n54), .A(n55), 
        .ZN(n38) );
  INV_X1 U98 ( .A(n132), .ZN(n11) );
  AOI21_X1 U99 ( .B1(n104), .B2(n105), .A(n100), .ZN(cw1[2]) );
  OAI21_X1 U100 ( .B1(n131), .B2(n26), .A(n7), .ZN(cw1[0]) );
  OAI21_X1 U101 ( .B1(n106), .B2(n107), .A(n7), .ZN(cw1[1]) );
  OR4_X1 U102 ( .A1(func[7]), .A2(func[10]), .A3(func[9]), .A4(func[8]), .ZN(
        n130) );
  NAND2_X1 U103 ( .A1(n52), .A2(n14), .ZN(n51) );
  NOR3_X1 U104 ( .A1(opcode[1]), .A2(opcode[5]), .A3(n25), .ZN(n89) );
  AOI211_X1 U105 ( .C1(opcode[1]), .C2(n90), .A(n12), .B(n137), .ZN(n108) );
  NOR3_X1 U106 ( .A1(opcode[1]), .A2(opcode[3]), .A3(n115), .ZN(n132) );
  AOI21_X1 U107 ( .B1(opcode[3]), .B2(opcode[1]), .A(n50), .ZN(n134) );
  NAND2_X1 U108 ( .A1(opcode[1]), .A2(n27), .ZN(n85) );
  INV_X1 U109 ( .A(opcode[1]), .ZN(n23) );
  AOI21_X1 U110 ( .B1(n23), .B2(n56), .A(opcode[3]), .ZN(n55) );
  AND3_X1 U111 ( .A1(n64), .A2(opcode[4]), .A3(opcode[3]), .ZN(n63) );
  OAI21_X1 U112 ( .B1(opcode[3]), .B2(n65), .A(n66), .ZN(n62) );
  OAI222_X1 U113 ( .A1(n66), .A2(n65), .B1(opcode[3]), .B2(n67), .C1(opcode[4]), .C2(n68), .ZN(n61) );
  AOI22_X1 U114 ( .A1(opcode[3]), .A2(n88), .B1(n57), .B2(n25), .ZN(n87) );
  NOR3_X1 U115 ( .A1(n100), .A2(opcode[3]), .A3(n64), .ZN(cw1[6]) );
  NAND2_X1 U116 ( .A1(opcode[3]), .A2(opcode[2]), .ZN(n66) );
  INV_X1 U117 ( .A(opcode[3]), .ZN(n25) );
  OAI222_X1 U118 ( .A1(opcode[5]), .A2(n38), .B1(n39), .B2(n26), .C1(n40), 
        .C2(n41), .ZN(cw1[9]) );
  AOI22_X1 U119 ( .A1(n83), .A2(n26), .B1(opcode[5]), .B2(n84), .ZN(n82) );
  NOR2_X1 U120 ( .A1(n23), .A2(opcode[5]), .ZN(n91) );
  OAI21_X1 U121 ( .B1(opcode[5]), .B2(n108), .A(n109), .ZN(cw1[13]) );
  OAI21_X1 U122 ( .B1(opcode[5]), .B2(n9), .A(n109), .ZN(cw1[12]) );
  AOI211_X1 U123 ( .C1(n120), .C2(opcode[5]), .A(n16), .B(n89), .ZN(n112) );
  AOI21_X1 U124 ( .B1(n14), .B2(n124), .A(opcode[5]), .ZN(n123) );
  NAND2_X1 U125 ( .A1(opcode[5]), .A2(opcode[4]), .ZN(n107) );
  NAND2_X1 U126 ( .A1(opcode[5]), .A2(n13), .ZN(n100) );
  AOI21_X1 U127 ( .B1(n101), .B2(n108), .A(opcode[5]), .ZN(n136) );
  OAI21_X1 U128 ( .B1(n141), .B2(n86), .A(opcode[5]), .ZN(n109) );
  INV_X1 U129 ( .A(opcode[5]), .ZN(n26) );
  AOI221_X1 U130 ( .B1(opcode[0]), .B2(n49), .C1(n50), .C2(n13), .A(n51), .ZN(
        n39) );
  OAI21_X1 U131 ( .B1(opcode[0]), .B2(opcode[4]), .A(n19), .ZN(n56) );
  NAND2_X1 U132 ( .A1(opcode[0]), .A2(n13), .ZN(n88) );
  NAND2_X1 U133 ( .A1(opcode[0]), .A2(n23), .ZN(n65) );
  NOR3_X1 U134 ( .A1(n13), .A2(opcode[0]), .A3(n19), .ZN(n115) );
  INV_X1 U135 ( .A(opcode[0]), .ZN(n27) );
  AOI22_X1 U136 ( .A1(opcode[4]), .A2(n89), .B1(n90), .B2(n91), .ZN(n58) );
  AOI211_X1 U137 ( .C1(opcode[4]), .C2(n21), .A(n132), .B(n133), .ZN(n131) );
  NOR3_X1 U138 ( .A1(n102), .A2(opcode[4]), .A3(n27), .ZN(n133) );
  NAND2_X1 U139 ( .A1(opcode[4]), .A2(n25), .ZN(n53) );
  OAI21_X1 U140 ( .B1(opcode[4]), .B2(n104), .A(n11), .ZN(n86) );
  INV_X1 U141 ( .A(opcode[4]), .ZN(n13) );
  OAI21_X1 U142 ( .B1(opcode[2]), .B2(n87), .A(n67), .ZN(n83) );
  NOR2_X1 U143 ( .A1(n85), .A2(opcode[2]), .ZN(n64) );
  NAND2_X1 U144 ( .A1(opcode[2]), .A2(n25), .ZN(n105) );
  AOI221_X1 U145 ( .B1(n17), .B2(n23), .C1(n22), .C2(opcode[2]), .A(n21), .ZN(
        n106) );
  INV_X1 U146 ( .A(opcode[2]), .ZN(n19) );
  CLKBUF_X1 U161 ( .A(rst), .Z(n2) );
  CLKBUF_X1 U162 ( .A(rst), .Z(n3) );
  CLKBUF_X1 U163 ( .A(rst), .Z(n4) );
  CLKBUF_X1 U164 ( .A(rst), .Z(n5) );
  CLKBUF_X1 U165 ( .A(rst), .Z(n6) );
endmodule


module MUX21_0 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n3, n1;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_593 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_592 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_591 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_590 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_589 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_588 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_587 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_586 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_585 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_584 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_583 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_582 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_581 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_580 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_579 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_578 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_577 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_576 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_575 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_574 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_573 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_572 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_571 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_570 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_569 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_568 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_567 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_566 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_565 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_564 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_563 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_GENERIC_NBIT32_0 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   n1, n2, n3;

  MUX21_0 MUXES_0 ( .A(A[0]), .B(B[0]), .S(n3), .Y(Y[0]) );
  MUX21_593 MUXES_1 ( .A(A[1]), .B(B[1]), .S(n1), .Y(Y[1]) );
  MUX21_592 MUXES_2 ( .A(A[2]), .B(B[2]), .S(n1), .Y(Y[2]) );
  MUX21_591 MUXES_3 ( .A(A[3]), .B(B[3]), .S(n1), .Y(Y[3]) );
  MUX21_590 MUXES_4 ( .A(A[4]), .B(B[4]), .S(n1), .Y(Y[4]) );
  MUX21_589 MUXES_5 ( .A(A[5]), .B(B[5]), .S(n1), .Y(Y[5]) );
  MUX21_588 MUXES_6 ( .A(A[6]), .B(B[6]), .S(n1), .Y(Y[6]) );
  MUX21_587 MUXES_7 ( .A(A[7]), .B(B[7]), .S(n1), .Y(Y[7]) );
  MUX21_586 MUXES_8 ( .A(A[8]), .B(B[8]), .S(n1), .Y(Y[8]) );
  MUX21_585 MUXES_9 ( .A(A[9]), .B(B[9]), .S(n1), .Y(Y[9]) );
  MUX21_584 MUXES_10 ( .A(A[10]), .B(B[10]), .S(n1), .Y(Y[10]) );
  MUX21_583 MUXES_11 ( .A(A[11]), .B(B[11]), .S(n1), .Y(Y[11]) );
  MUX21_582 MUXES_12 ( .A(A[12]), .B(B[12]), .S(n1), .Y(Y[12]) );
  MUX21_581 MUXES_13 ( .A(A[13]), .B(B[13]), .S(n2), .Y(Y[13]) );
  MUX21_580 MUXES_14 ( .A(A[14]), .B(B[14]), .S(n2), .Y(Y[14]) );
  MUX21_579 MUXES_15 ( .A(A[15]), .B(B[15]), .S(n2), .Y(Y[15]) );
  MUX21_578 MUXES_16 ( .A(A[16]), .B(B[16]), .S(n2), .Y(Y[16]) );
  MUX21_577 MUXES_17 ( .A(A[17]), .B(B[17]), .S(n2), .Y(Y[17]) );
  MUX21_576 MUXES_18 ( .A(A[18]), .B(B[18]), .S(n2), .Y(Y[18]) );
  MUX21_575 MUXES_19 ( .A(A[19]), .B(B[19]), .S(n2), .Y(Y[19]) );
  MUX21_574 MUXES_20 ( .A(A[20]), .B(B[20]), .S(n2), .Y(Y[20]) );
  MUX21_573 MUXES_21 ( .A(A[21]), .B(B[21]), .S(n2), .Y(Y[21]) );
  MUX21_572 MUXES_22 ( .A(A[22]), .B(B[22]), .S(n2), .Y(Y[22]) );
  MUX21_571 MUXES_23 ( .A(A[23]), .B(B[23]), .S(n2), .Y(Y[23]) );
  MUX21_570 MUXES_24 ( .A(A[24]), .B(B[24]), .S(n2), .Y(Y[24]) );
  MUX21_569 MUXES_25 ( .A(A[25]), .B(B[25]), .S(n3), .Y(Y[25]) );
  MUX21_568 MUXES_26 ( .A(A[26]), .B(B[26]), .S(n3), .Y(Y[26]) );
  MUX21_567 MUXES_27 ( .A(A[27]), .B(B[27]), .S(n3), .Y(Y[27]) );
  MUX21_566 MUXES_28 ( .A(A[28]), .B(B[28]), .S(n3), .Y(Y[28]) );
  MUX21_565 MUXES_29 ( .A(A[29]), .B(B[29]), .S(n3), .Y(Y[29]) );
  MUX21_564 MUXES_30 ( .A(A[30]), .B(B[30]), .S(n3), .Y(Y[30]) );
  MUX21_563 MUXES_31 ( .A(A[31]), .B(B[31]), .S(n3), .Y(Y[31]) );
  BUF_X1 U1 ( .A(SEL), .Z(n2) );
  BUF_X1 U2 ( .A(SEL), .Z(n1) );
  BUF_X1 U3 ( .A(SEL), .Z(n3) );
endmodule


module MUX21_530 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_529 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_528 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_527 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_526 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_525 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_524 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_523 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_522 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_521 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_520 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_519 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_518 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_517 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_516 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_515 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_514 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_513 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_512 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_511 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_510 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_509 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_508 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_507 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_506 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_505 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_504 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  AOI22_X1 U1 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_503 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_502 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_501 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_500 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_499 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_GENERIC_NBIT32_4 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   n1, n2;

  MUX21_530 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_529 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_528 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_527 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
  MUX21_526 MUXES_4 ( .A(A[4]), .B(B[4]), .S(SEL), .Y(Y[4]) );
  MUX21_525 MUXES_5 ( .A(A[5]), .B(B[5]), .S(n2), .Y(Y[5]) );
  MUX21_524 MUXES_6 ( .A(A[6]), .B(B[6]), .S(n1), .Y(Y[6]) );
  MUX21_523 MUXES_7 ( .A(A[7]), .B(B[7]), .S(n1), .Y(Y[7]) );
  MUX21_522 MUXES_8 ( .A(A[8]), .B(B[8]), .S(n1), .Y(Y[8]) );
  MUX21_521 MUXES_9 ( .A(A[9]), .B(B[9]), .S(n1), .Y(Y[9]) );
  MUX21_520 MUXES_10 ( .A(A[10]), .B(B[10]), .S(n2), .Y(Y[10]) );
  MUX21_519 MUXES_11 ( .A(A[11]), .B(B[11]), .S(n1), .Y(Y[11]) );
  MUX21_518 MUXES_12 ( .A(A[12]), .B(B[12]), .S(n1), .Y(Y[12]) );
  MUX21_517 MUXES_13 ( .A(A[13]), .B(B[13]), .S(n1), .Y(Y[13]) );
  MUX21_516 MUXES_14 ( .A(A[14]), .B(B[14]), .S(n1), .Y(Y[14]) );
  MUX21_515 MUXES_15 ( .A(A[15]), .B(B[15]), .S(n1), .Y(Y[15]) );
  MUX21_514 MUXES_16 ( .A(A[16]), .B(B[16]), .S(n1), .Y(Y[16]) );
  MUX21_513 MUXES_17 ( .A(A[17]), .B(B[17]), .S(n1), .Y(Y[17]) );
  MUX21_512 MUXES_18 ( .A(A[18]), .B(B[18]), .S(n1), .Y(Y[18]) );
  MUX21_511 MUXES_19 ( .A(A[19]), .B(B[19]), .S(n1), .Y(Y[19]) );
  MUX21_510 MUXES_20 ( .A(A[20]), .B(B[20]), .S(n1), .Y(Y[20]) );
  MUX21_509 MUXES_21 ( .A(A[21]), .B(B[21]), .S(n1), .Y(Y[21]) );
  MUX21_508 MUXES_22 ( .A(A[22]), .B(B[22]), .S(n1), .Y(Y[22]) );
  MUX21_507 MUXES_23 ( .A(A[23]), .B(B[23]), .S(n1), .Y(Y[23]) );
  MUX21_506 MUXES_24 ( .A(A[24]), .B(B[24]), .S(n2), .Y(Y[24]) );
  MUX21_505 MUXES_25 ( .A(A[25]), .B(B[25]), .S(n2), .Y(Y[25]) );
  MUX21_504 MUXES_26 ( .A(A[26]), .B(B[26]), .S(n2), .Y(Y[26]) );
  MUX21_503 MUXES_27 ( .A(A[27]), .B(B[27]), .S(n1), .Y(Y[27]) );
  MUX21_502 MUXES_28 ( .A(A[28]), .B(B[28]), .S(n2), .Y(Y[28]) );
  MUX21_501 MUXES_29 ( .A(A[29]), .B(B[29]), .S(n1), .Y(Y[29]) );
  MUX21_500 MUXES_30 ( .A(A[30]), .B(B[30]), .S(SEL), .Y(Y[30]) );
  MUX21_499 MUXES_31 ( .A(A[31]), .B(B[31]), .S(SEL), .Y(Y[31]) );
  BUF_X2 U1 ( .A(SEL), .Z(n1) );
  CLKBUF_X1 U2 ( .A(SEL), .Z(n2) );
endmodule


module FETCH_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   \A[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n57;
  assign SUM[1] = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  AND2_X1 U1 ( .A1(A[3]), .A2(A[2]), .ZN(n1) );
  AND2_X1 U2 ( .A1(A[10]), .A2(n12), .ZN(n2) );
  AND2_X1 U3 ( .A1(A[26]), .A2(n7), .ZN(n3) );
  AND2_X1 U4 ( .A1(A[6]), .A2(n27), .ZN(n4) );
  AND2_X1 U5 ( .A1(A[7]), .A2(n4), .ZN(n5) );
  AND2_X1 U6 ( .A1(A[24]), .A2(n25), .ZN(n6) );
  AND2_X1 U7 ( .A1(A[25]), .A2(n6), .ZN(n7) );
  AND2_X1 U8 ( .A1(A[27]), .A2(n3), .ZN(n8) );
  AND2_X1 U9 ( .A1(A[28]), .A2(n8), .ZN(n9) );
  AND2_X1 U10 ( .A1(A[29]), .A2(n9), .ZN(n10) );
  AND2_X1 U11 ( .A1(A[8]), .A2(n5), .ZN(n11) );
  AND2_X1 U12 ( .A1(A[9]), .A2(n11), .ZN(n12) );
  AND2_X1 U13 ( .A1(A[11]), .A2(n2), .ZN(n13) );
  AND2_X1 U14 ( .A1(A[12]), .A2(n13), .ZN(n14) );
  AND2_X1 U15 ( .A1(A[13]), .A2(n14), .ZN(n15) );
  AND2_X1 U16 ( .A1(A[14]), .A2(n15), .ZN(n16) );
  AND2_X1 U17 ( .A1(A[15]), .A2(n16), .ZN(n17) );
  AND2_X1 U18 ( .A1(A[16]), .A2(n17), .ZN(n18) );
  AND2_X1 U19 ( .A1(A[17]), .A2(n18), .ZN(n19) );
  AND2_X1 U20 ( .A1(A[18]), .A2(n19), .ZN(n20) );
  AND2_X1 U21 ( .A1(A[19]), .A2(n20), .ZN(n21) );
  AND2_X1 U22 ( .A1(A[20]), .A2(n21), .ZN(n22) );
  AND2_X1 U23 ( .A1(A[21]), .A2(n22), .ZN(n23) );
  AND2_X1 U24 ( .A1(A[22]), .A2(n23), .ZN(n24) );
  AND2_X1 U25 ( .A1(A[23]), .A2(n24), .ZN(n25) );
  AND2_X1 U26 ( .A1(A[4]), .A2(n1), .ZN(n26) );
  AND2_X1 U27 ( .A1(A[5]), .A2(n26), .ZN(n27) );
  NAND2_X1 U28 ( .A1(A[30]), .A2(n10), .ZN(n57) );
  XOR2_X1 U29 ( .A(A[26]), .B(n7), .Z(SUM[26]) );
  XOR2_X1 U30 ( .A(A[27]), .B(n3), .Z(SUM[27]) );
  XOR2_X1 U31 ( .A(A[30]), .B(n10), .Z(SUM[30]) );
  XOR2_X1 U32 ( .A(A[29]), .B(n9), .Z(SUM[29]) );
  XOR2_X1 U33 ( .A(A[28]), .B(n8), .Z(SUM[28]) );
  XOR2_X1 U34 ( .A(A[25]), .B(n6), .Z(SUM[25]) );
  XOR2_X1 U35 ( .A(A[24]), .B(n25), .Z(SUM[24]) );
  XOR2_X1 U36 ( .A(A[23]), .B(n24), .Z(SUM[23]) );
  XOR2_X1 U37 ( .A(A[22]), .B(n23), .Z(SUM[22]) );
  XOR2_X1 U38 ( .A(A[21]), .B(n22), .Z(SUM[21]) );
  XOR2_X1 U39 ( .A(A[20]), .B(n21), .Z(SUM[20]) );
  XNOR2_X1 U40 ( .A(A[31]), .B(n57), .ZN(SUM[31]) );
  XOR2_X1 U41 ( .A(A[10]), .B(n12), .Z(SUM[10]) );
  XOR2_X1 U42 ( .A(A[11]), .B(n2), .Z(SUM[11]) );
  XOR2_X1 U43 ( .A(A[19]), .B(n20), .Z(SUM[19]) );
  XOR2_X1 U44 ( .A(A[18]), .B(n19), .Z(SUM[18]) );
  XOR2_X1 U45 ( .A(A[17]), .B(n18), .Z(SUM[17]) );
  XOR2_X1 U46 ( .A(A[16]), .B(n17), .Z(SUM[16]) );
  XOR2_X1 U47 ( .A(A[15]), .B(n16), .Z(SUM[15]) );
  XOR2_X1 U48 ( .A(A[14]), .B(n15), .Z(SUM[14]) );
  XOR2_X1 U49 ( .A(A[13]), .B(n14), .Z(SUM[13]) );
  XOR2_X1 U50 ( .A(A[12]), .B(n13), .Z(SUM[12]) );
  XOR2_X1 U51 ( .A(A[9]), .B(n11), .Z(SUM[9]) );
  INV_X1 U52 ( .A(A[2]), .ZN(SUM[2]) );
  XOR2_X1 U53 ( .A(A[3]), .B(A[2]), .Z(SUM[3]) );
  XOR2_X1 U54 ( .A(A[4]), .B(n1), .Z(SUM[4]) );
  XOR2_X1 U55 ( .A(A[8]), .B(n5), .Z(SUM[8]) );
  XOR2_X1 U56 ( .A(A[7]), .B(n4), .Z(SUM[7]) );
  XOR2_X1 U57 ( .A(A[6]), .B(n27), .Z(SUM[6]) );
  XOR2_X1 U58 ( .A(A[5]), .B(n26), .Z(SUM[5]) );
endmodule


module FETCH ( PC, hazard_PC, PC_sel, IRAM_addr, NPC );
  input [31:0] PC;
  input [31:0] hazard_PC;
  output [31:0] IRAM_addr;
  output [31:0] NPC;
  input PC_sel;


  MUX21_GENERIC_NBIT32_4 MUX ( .A(PC), .B(hazard_PC), .SEL(PC_sel), .Y(
        IRAM_addr) );
  FETCH_DW01_add_0 add_37 ( .A(IRAM_addr), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b1, 1'b0, 1'b0}), .CI(1'b0), .SUM(NPC) );
endmodule


module MUX21_562 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_561 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_560 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_559 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_558 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_557 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_556 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_555 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_554 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_553 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_552 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_551 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_550 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_549 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_548 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_547 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_546 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_545 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_544 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_543 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_542 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_541 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_540 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_539 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_538 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_537 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_536 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_535 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_534 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_533 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_532 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  AOI22_X1 U1 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_531 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_GENERIC_NBIT32_5 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   n1, n2, n3;

  MUX21_562 MUXES_0 ( .A(A[0]), .B(B[0]), .S(n1), .Y(Y[0]) );
  MUX21_561 MUXES_1 ( .A(A[1]), .B(B[1]), .S(n1), .Y(Y[1]) );
  MUX21_560 MUXES_2 ( .A(A[2]), .B(B[2]), .S(n1), .Y(Y[2]) );
  MUX21_559 MUXES_3 ( .A(A[3]), .B(B[3]), .S(n1), .Y(Y[3]) );
  MUX21_558 MUXES_4 ( .A(A[4]), .B(B[4]), .S(n1), .Y(Y[4]) );
  MUX21_557 MUXES_5 ( .A(A[5]), .B(B[5]), .S(n1), .Y(Y[5]) );
  MUX21_556 MUXES_6 ( .A(A[6]), .B(B[6]), .S(n1), .Y(Y[6]) );
  MUX21_555 MUXES_7 ( .A(A[7]), .B(B[7]), .S(n1), .Y(Y[7]) );
  MUX21_554 MUXES_8 ( .A(A[8]), .B(B[8]), .S(n1), .Y(Y[8]) );
  MUX21_553 MUXES_9 ( .A(A[9]), .B(B[9]), .S(n1), .Y(Y[9]) );
  MUX21_552 MUXES_10 ( .A(A[10]), .B(B[10]), .S(n1), .Y(Y[10]) );
  MUX21_551 MUXES_11 ( .A(A[11]), .B(B[11]), .S(n1), .Y(Y[11]) );
  MUX21_550 MUXES_12 ( .A(A[12]), .B(B[12]), .S(n2), .Y(Y[12]) );
  MUX21_549 MUXES_13 ( .A(A[13]), .B(B[13]), .S(n2), .Y(Y[13]) );
  MUX21_548 MUXES_14 ( .A(A[14]), .B(B[14]), .S(n2), .Y(Y[14]) );
  MUX21_547 MUXES_15 ( .A(A[15]), .B(B[15]), .S(n2), .Y(Y[15]) );
  MUX21_546 MUXES_16 ( .A(A[16]), .B(B[16]), .S(n2), .Y(Y[16]) );
  MUX21_545 MUXES_17 ( .A(A[17]), .B(B[17]), .S(n2), .Y(Y[17]) );
  MUX21_544 MUXES_18 ( .A(A[18]), .B(B[18]), .S(n2), .Y(Y[18]) );
  MUX21_543 MUXES_19 ( .A(A[19]), .B(B[19]), .S(n2), .Y(Y[19]) );
  MUX21_542 MUXES_20 ( .A(A[20]), .B(B[20]), .S(n2), .Y(Y[20]) );
  MUX21_541 MUXES_21 ( .A(A[21]), .B(B[21]), .S(n2), .Y(Y[21]) );
  MUX21_540 MUXES_22 ( .A(A[22]), .B(B[22]), .S(n2), .Y(Y[22]) );
  MUX21_539 MUXES_23 ( .A(A[23]), .B(B[23]), .S(n2), .Y(Y[23]) );
  MUX21_538 MUXES_24 ( .A(A[24]), .B(B[24]), .S(n3), .Y(Y[24]) );
  MUX21_537 MUXES_25 ( .A(A[25]), .B(B[25]), .S(n3), .Y(Y[25]) );
  MUX21_536 MUXES_26 ( .A(A[26]), .B(B[26]), .S(n3), .Y(Y[26]) );
  MUX21_535 MUXES_27 ( .A(A[27]), .B(B[27]), .S(n3), .Y(Y[27]) );
  MUX21_534 MUXES_28 ( .A(A[28]), .B(B[28]), .S(n3), .Y(Y[28]) );
  MUX21_533 MUXES_29 ( .A(A[29]), .B(B[29]), .S(n3), .Y(Y[29]) );
  MUX21_532 MUXES_30 ( .A(A[30]), .B(B[30]), .S(n3), .Y(Y[30]) );
  MUX21_531 MUXES_31 ( .A(A[31]), .B(B[31]), .S(n3), .Y(Y[31]) );
  BUF_X1 U1 ( .A(SEL), .Z(n2) );
  BUF_X1 U2 ( .A(SEL), .Z(n1) );
  BUF_X1 U3 ( .A(SEL), .Z(n3) );
endmodule


module dec_logic_WORD_size32_NREG32 ( instr, NPC_in, opcode, RS1, RS2, RD, 
        FUNC, IMM, IMM26 );
  input [31:0] instr;
  input [31:0] NPC_in;
  output [5:0] opcode;
  output [4:0] RS1;
  output [4:0] RS2;
  output [4:0] RD;
  output [10:0] FUNC;
  output [15:0] IMM;
  output [25:0] IMM26;
  wire   \instr[31] , \instr[30] , \instr[29] , \instr[28] , \instr[27] ,
         \instr[26] , N246, N247, N248, N249, N250, N251, N252, N253, N254,
         N255, N256, N257, N258, N259, N260, N261, N262, N263, N264, N265,
         N266, N267, N268, N269, N270, N271, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n65,
         n66, n67, n68, n69, n70;
  assign opcode[5] = \instr[31] ;
  assign \instr[31]  = instr[31];
  assign opcode[4] = \instr[30] ;
  assign \instr[30]  = instr[30];
  assign opcode[3] = \instr[29] ;
  assign \instr[29]  = instr[29];
  assign opcode[2] = \instr[28] ;
  assign \instr[28]  = instr[28];
  assign opcode[1] = \instr[27] ;
  assign \instr[27]  = instr[27];
  assign opcode[0] = \instr[26] ;
  assign \instr[26]  = instr[26];

  DLL_X1 \IMM26_reg[25]  ( .D(N271), .GN(n4), .Q(IMM26[25]) );
  DLL_X1 \IMM26_reg[24]  ( .D(N270), .GN(n4), .Q(IMM26[24]) );
  DLL_X1 \IMM26_reg[23]  ( .D(N269), .GN(n4), .Q(IMM26[23]) );
  DLL_X1 \IMM26_reg[22]  ( .D(N268), .GN(n4), .Q(IMM26[22]) );
  DLL_X1 \IMM26_reg[21]  ( .D(N267), .GN(n4), .Q(IMM26[21]) );
  DLL_X1 \IMM26_reg[20]  ( .D(N266), .GN(n4), .Q(IMM26[20]) );
  DLL_X1 \IMM26_reg[19]  ( .D(N265), .GN(n4), .Q(IMM26[19]) );
  DLL_X1 \IMM26_reg[18]  ( .D(N264), .GN(n4), .Q(IMM26[18]) );
  DLL_X1 \IMM26_reg[17]  ( .D(N263), .GN(n4), .Q(IMM26[17]) );
  DLL_X1 \IMM26_reg[16]  ( .D(N262), .GN(n4), .Q(IMM26[16]) );
  DLL_X1 \IMM26_reg[15]  ( .D(N261), .GN(n5), .Q(IMM26[15]) );
  DLL_X1 \IMM26_reg[14]  ( .D(N260), .GN(n5), .Q(IMM26[14]) );
  DLL_X1 \IMM26_reg[13]  ( .D(N259), .GN(n5), .Q(IMM26[13]) );
  DLL_X1 \IMM26_reg[12]  ( .D(N258), .GN(n5), .Q(IMM26[12]) );
  DLL_X1 \IMM26_reg[11]  ( .D(N257), .GN(n5), .Q(IMM26[11]) );
  DLL_X1 \IMM26_reg[10]  ( .D(N256), .GN(n5), .Q(IMM26[10]) );
  DLL_X1 \IMM26_reg[9]  ( .D(N255), .GN(n5), .Q(IMM26[9]) );
  DLL_X1 \IMM26_reg[8]  ( .D(N254), .GN(n5), .Q(IMM26[8]) );
  DLL_X1 \IMM26_reg[7]  ( .D(N253), .GN(n5), .Q(IMM26[7]) );
  DLL_X1 \IMM26_reg[6]  ( .D(N252), .GN(n5), .Q(IMM26[6]) );
  DLL_X1 \IMM26_reg[5]  ( .D(N251), .GN(n6), .Q(IMM26[5]) );
  DLL_X1 \IMM26_reg[4]  ( .D(N250), .GN(n6), .Q(IMM26[4]) );
  DLL_X1 \IMM26_reg[3]  ( .D(N249), .GN(n6), .Q(IMM26[3]) );
  DLL_X1 \IMM26_reg[2]  ( .D(N248), .GN(n6), .Q(IMM26[2]) );
  DLL_X1 \IMM26_reg[1]  ( .D(N247), .GN(n6), .Q(IMM26[1]) );
  DLL_X1 \IMM26_reg[0]  ( .D(N246), .GN(n6), .Q(IMM26[0]) );
  NAND3_X1 U134 ( .A1(n39), .A2(n1), .A3(instr[15]), .ZN(n46) );
  AND2_X1 U3 ( .A1(n36), .A2(n41), .ZN(n33) );
  NOR2_X1 U4 ( .A1(n68), .A2(n32), .ZN(RS1[4]) );
  NOR2_X1 U5 ( .A1(n68), .A2(n28), .ZN(RS1[0]) );
  BUF_X1 U6 ( .A(n36), .Z(n2) );
  INV_X1 U7 ( .A(n34), .ZN(n68) );
  OR2_X1 U8 ( .A1(n45), .A2(n65), .ZN(n47) );
  NOR2_X1 U9 ( .A1(n68), .A2(n29), .ZN(RS1[1]) );
  NOR2_X1 U10 ( .A1(n68), .A2(n30), .ZN(RS1[2]) );
  NOR2_X1 U11 ( .A1(n68), .A2(n31), .ZN(RS1[3]) );
  INV_X1 U12 ( .A(n37), .ZN(n66) );
  NAND2_X1 U13 ( .A1(n39), .A2(n1), .ZN(n45) );
  INV_X1 U14 ( .A(n39), .ZN(n67) );
  OAI21_X1 U15 ( .B1(n1), .B2(n22), .A(n46), .ZN(N261) );
  OAI21_X1 U16 ( .B1(n1), .B2(n23), .A(n46), .ZN(N262) );
  OAI21_X1 U17 ( .B1(n1), .B2(n24), .A(n46), .ZN(N263) );
  OAI21_X1 U18 ( .B1(n1), .B2(n25), .A(n46), .ZN(N264) );
  OAI21_X1 U19 ( .B1(n1), .B2(n26), .A(n46), .ZN(N265) );
  OAI21_X1 U20 ( .B1(n1), .B2(n27), .A(n46), .ZN(N266) );
  OAI21_X1 U21 ( .B1(n1), .B2(n28), .A(n46), .ZN(N267) );
  OAI21_X1 U22 ( .B1(n1), .B2(n29), .A(n46), .ZN(N268) );
  OAI21_X1 U23 ( .B1(n1), .B2(n30), .A(n46), .ZN(N269) );
  OAI21_X1 U24 ( .B1(n1), .B2(n31), .A(n46), .ZN(N270) );
  OAI21_X1 U25 ( .B1(n1), .B2(n32), .A(n46), .ZN(N271) );
  BUF_X1 U26 ( .A(n44), .Z(n5) );
  BUF_X1 U27 ( .A(n44), .Z(n4) );
  NOR2_X1 U28 ( .A1(n67), .A2(n7), .ZN(N246) );
  NOR2_X1 U29 ( .A1(n67), .A2(n8), .ZN(N247) );
  NOR2_X1 U30 ( .A1(n67), .A2(n9), .ZN(N248) );
  NOR2_X1 U31 ( .A1(n67), .A2(n10), .ZN(N249) );
  NOR2_X1 U32 ( .A1(n67), .A2(n11), .ZN(N250) );
  NOR2_X1 U33 ( .A1(n67), .A2(n12), .ZN(N251) );
  NOR2_X1 U34 ( .A1(n67), .A2(n13), .ZN(N252) );
  NOR2_X1 U35 ( .A1(n67), .A2(n14), .ZN(N253) );
  NOR2_X1 U36 ( .A1(n67), .A2(n15), .ZN(N254) );
  NOR2_X1 U37 ( .A1(n67), .A2(n16), .ZN(N255) );
  NOR2_X1 U38 ( .A1(n67), .A2(n17), .ZN(N256) );
  NOR2_X1 U39 ( .A1(n67), .A2(n18), .ZN(N257) );
  NOR2_X1 U40 ( .A1(n67), .A2(n19), .ZN(N258) );
  NOR2_X1 U41 ( .A1(n67), .A2(n20), .ZN(N259) );
  NOR2_X1 U42 ( .A1(n67), .A2(n21), .ZN(N260) );
  BUF_X1 U43 ( .A(n44), .Z(n6) );
  NOR4_X1 U44 ( .A1(n69), .A2(\instr[28] ), .A3(\instr[29] ), .A4(\instr[31] ), 
        .ZN(n64) );
  INV_X1 U45 ( .A(instr[11]), .ZN(n18) );
  INV_X1 U46 ( .A(instr[12]), .ZN(n19) );
  INV_X1 U47 ( .A(instr[14]), .ZN(n21) );
  INV_X1 U48 ( .A(instr[13]), .ZN(n20) );
  INV_X1 U49 ( .A(instr[16]), .ZN(n23) );
  INV_X1 U50 ( .A(instr[17]), .ZN(n24) );
  INV_X1 U51 ( .A(instr[18]), .ZN(n25) );
  INV_X1 U52 ( .A(instr[19]), .ZN(n26) );
  INV_X1 U53 ( .A(instr[20]), .ZN(n27) );
  INV_X1 U54 ( .A(instr[25]), .ZN(n32) );
  INV_X1 U55 ( .A(instr[24]), .ZN(n31) );
  INV_X1 U56 ( .A(instr[23]), .ZN(n30) );
  INV_X1 U57 ( .A(instr[22]), .ZN(n29) );
  INV_X1 U58 ( .A(instr[21]), .ZN(n28) );
  INV_X1 U59 ( .A(instr[15]), .ZN(n22) );
  OAI21_X1 U60 ( .B1(n65), .B2(n46), .A(n57), .ZN(IMM[15]) );
  NAND2_X1 U61 ( .A1(NPC_in[15]), .A2(n66), .ZN(n57) );
  OAI21_X1 U62 ( .B1(n21), .B2(n47), .A(n58), .ZN(IMM[14]) );
  NAND2_X1 U63 ( .A1(NPC_in[14]), .A2(n66), .ZN(n58) );
  OAI21_X1 U64 ( .B1(n20), .B2(n47), .A(n59), .ZN(IMM[13]) );
  NAND2_X1 U65 ( .A1(NPC_in[13]), .A2(n66), .ZN(n59) );
  OAI21_X1 U66 ( .B1(n19), .B2(n47), .A(n60), .ZN(IMM[12]) );
  NAND2_X1 U67 ( .A1(NPC_in[12]), .A2(n66), .ZN(n60) );
  OAI21_X1 U68 ( .B1(n18), .B2(n47), .A(n61), .ZN(IMM[11]) );
  NAND2_X1 U69 ( .A1(NPC_in[11]), .A2(n66), .ZN(n61) );
  OAI21_X1 U70 ( .B1(n17), .B2(n47), .A(n62), .ZN(IMM[10]) );
  NAND2_X1 U71 ( .A1(NPC_in[10]), .A2(n66), .ZN(n62) );
  OAI21_X1 U72 ( .B1(n16), .B2(n47), .A(n48), .ZN(IMM[9]) );
  NAND2_X1 U73 ( .A1(NPC_in[9]), .A2(n66), .ZN(n48) );
  OAI21_X1 U74 ( .B1(n15), .B2(n47), .A(n49), .ZN(IMM[8]) );
  NAND2_X1 U75 ( .A1(NPC_in[8]), .A2(n66), .ZN(n49) );
  OAI21_X1 U76 ( .B1(n14), .B2(n47), .A(n50), .ZN(IMM[7]) );
  NAND2_X1 U77 ( .A1(NPC_in[7]), .A2(n66), .ZN(n50) );
  OAI21_X1 U78 ( .B1(n13), .B2(n47), .A(n51), .ZN(IMM[6]) );
  NAND2_X1 U79 ( .A1(NPC_in[6]), .A2(n66), .ZN(n51) );
  OAI21_X1 U80 ( .B1(n12), .B2(n47), .A(n52), .ZN(IMM[5]) );
  NAND2_X1 U81 ( .A1(NPC_in[5]), .A2(n66), .ZN(n52) );
  OAI21_X1 U82 ( .B1(n11), .B2(n47), .A(n53), .ZN(IMM[4]) );
  NAND2_X1 U83 ( .A1(NPC_in[4]), .A2(n66), .ZN(n53) );
  OAI21_X1 U84 ( .B1(n10), .B2(n47), .A(n54), .ZN(IMM[3]) );
  NAND2_X1 U85 ( .A1(NPC_in[3]), .A2(n66), .ZN(n54) );
  OAI21_X1 U86 ( .B1(n9), .B2(n47), .A(n55), .ZN(IMM[2]) );
  NAND2_X1 U87 ( .A1(NPC_in[2]), .A2(n66), .ZN(n55) );
  OAI21_X1 U88 ( .B1(n8), .B2(n47), .A(n56), .ZN(IMM[1]) );
  NAND2_X1 U89 ( .A1(NPC_in[1]), .A2(n66), .ZN(n56) );
  OAI21_X1 U90 ( .B1(n7), .B2(n47), .A(n63), .ZN(IMM[0]) );
  NAND2_X1 U91 ( .A1(NPC_in[0]), .A2(n66), .ZN(n63) );
  INV_X1 U92 ( .A(instr[8]), .ZN(n15) );
  INV_X1 U93 ( .A(instr[9]), .ZN(n16) );
  INV_X1 U94 ( .A(instr[10]), .ZN(n17) );
  INV_X1 U95 ( .A(instr[7]), .ZN(n14) );
  INV_X1 U96 ( .A(instr[3]), .ZN(n10) );
  INV_X1 U97 ( .A(instr[4]), .ZN(n11) );
  INV_X1 U98 ( .A(instr[6]), .ZN(n13) );
  INV_X1 U99 ( .A(instr[5]), .ZN(n12) );
  INV_X1 U100 ( .A(instr[1]), .ZN(n8) );
  INV_X1 U101 ( .A(instr[2]), .ZN(n9) );
  INV_X1 U102 ( .A(instr[0]), .ZN(n7) );
  NAND2_X1 U103 ( .A1(\instr[26] ), .A2(n64), .ZN(n37) );
  NOR2_X1 U104 ( .A1(n33), .A2(n27), .ZN(RS2[4]) );
  NOR2_X1 U105 ( .A1(n33), .A2(n25), .ZN(RS2[2]) );
  NOR2_X1 U106 ( .A1(n33), .A2(n23), .ZN(RS2[0]) );
  NOR2_X1 U107 ( .A1(n33), .A2(n24), .ZN(RS2[1]) );
  NOR2_X1 U108 ( .A1(n33), .A2(n26), .ZN(RS2[3]) );
  NAND4_X1 U109 ( .A1(\instr[31] ), .A2(\instr[29] ), .A3(n42), .A4(n70), .ZN(
        n41) );
  CLKBUF_X1 U110 ( .A(n34), .Z(n1) );
  NAND2_X1 U111 ( .A1(n64), .A2(n70), .ZN(n34) );
  NAND2_X1 U112 ( .A1(n3), .A2(n43), .ZN(n36) );
  BUF_X1 U113 ( .A(n40), .Z(n3) );
  NOR4_X1 U114 ( .A1(\instr[27] ), .A2(\instr[29] ), .A3(\instr[30] ), .A4(
        \instr[31] ), .ZN(n40) );
  NOR2_X1 U115 ( .A1(\instr[28] ), .A2(\instr[26] ), .ZN(n43) );
  OAI221_X1 U116 ( .B1(n26), .B2(n35), .C1(n2), .C2(n21), .A(n37), .ZN(RD[3])
         );
  OAI221_X1 U117 ( .B1(n27), .B2(n35), .C1(n2), .C2(n22), .A(n37), .ZN(RD[4])
         );
  OAI221_X1 U118 ( .B1(n25), .B2(n35), .C1(n2), .C2(n20), .A(n37), .ZN(RD[2])
         );
  INV_X1 U119 ( .A(\instr[27] ), .ZN(n69) );
  OAI22_X1 U120 ( .A1(\instr[28] ), .A2(\instr[27] ), .B1(n43), .B2(n69), .ZN(
        n42) );
  OAI221_X1 U121 ( .B1(n23), .B2(n35), .C1(n2), .C2(n18), .A(n37), .ZN(RD[0])
         );
  OAI221_X1 U122 ( .B1(n24), .B2(n35), .C1(n2), .C2(n19), .A(n37), .ZN(RD[1])
         );
  NAND4_X1 U123 ( .A1(n33), .A2(n38), .A3(n39), .A4(n34), .ZN(n35) );
  AOI21_X1 U124 ( .B1(n3), .B2(\instr[28] ), .A(n45), .ZN(n44) );
  INV_X1 U125 ( .A(n2), .ZN(n65) );
  NOR2_X1 U126 ( .A1(n2), .A2(n11), .ZN(FUNC[4]) );
  NOR2_X1 U127 ( .A1(n2), .A2(n13), .ZN(FUNC[6]) );
  NOR2_X1 U128 ( .A1(n2), .A2(n12), .ZN(FUNC[5]) );
  NOR2_X1 U129 ( .A1(n2), .A2(n8), .ZN(FUNC[1]) );
  NOR2_X1 U130 ( .A1(n2), .A2(n7), .ZN(FUNC[0]) );
  NOR2_X1 U131 ( .A1(n2), .A2(n10), .ZN(FUNC[3]) );
  NOR2_X1 U132 ( .A1(n2), .A2(n9), .ZN(FUNC[2]) );
  NOR2_X1 U133 ( .A1(n2), .A2(n14), .ZN(FUNC[7]) );
  NOR2_X1 U135 ( .A1(n2), .A2(n17), .ZN(FUNC[10]) );
  NOR2_X1 U136 ( .A1(n2), .A2(n16), .ZN(FUNC[9]) );
  NOR2_X1 U137 ( .A1(n2), .A2(n15), .ZN(FUNC[8]) );
  NAND2_X1 U138 ( .A1(\instr[28] ), .A2(n3), .ZN(n38) );
  NAND2_X1 U139 ( .A1(\instr[30] ), .A2(n64), .ZN(n39) );
  INV_X1 U140 ( .A(\instr[30] ), .ZN(n70) );
endmodule


module my_xor_0 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_255 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_254 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_253 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_252 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_251 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_250 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_249 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_248 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_247 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_246 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_245 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_244 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_243 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_242 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_241 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_240 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_239 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_238 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_237 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_236 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_235 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_234 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_233 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_232 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_231 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_230 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_229 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_228 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_227 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_226 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_225 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module pg_net_0 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_250 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_249 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_248 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_247 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_246 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_245 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_244 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_243 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_242 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_241 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_240 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_239 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_238 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_237 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_236 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_235 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_234 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_233 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_232 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_231 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_230 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_229 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_228 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_227 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_226 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_225 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_224 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_223 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_222 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_221 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_BLOCK_0 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n2;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n2), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n2) );
endmodule


module PG_BLOCK_242 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_241 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AOI21_X1 U1 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U2 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U3 ( .A(n3), .ZN(PG_G) );
endmodule


module PG_BLOCK_240 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_239 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_238 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_237 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_236 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_235 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_234 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_233 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_232 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_231 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_230 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_229 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_0 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n2) );
endmodule


module PG_BLOCK_228 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_227 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_226 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_225 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_224 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_223 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_222 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_68 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_221 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_220 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_219 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_67 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_218 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AND2_X1 U2 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_217 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_66 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_65 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_64 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_63 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_62 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_61 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_0 ( A, B, Cin, Co );
  input [31:0] A;
  input [31:0] B;
  output [7:0] Co;
  input Cin;
  wire   \g_vector[4][31] , \g_vector[4][27] , \g_vector[3][31] ,
         \g_vector[3][23] , \g_vector[3][15] , \g_vector[2][31] ,
         \g_vector[2][27] , \g_vector[2][23] , \g_vector[2][19] ,
         \g_vector[2][15] , \g_vector[2][11] , \g_vector[2][7] ,
         \g_vector[1][31] , \g_vector[1][29] , \g_vector[1][27] ,
         \g_vector[1][25] , \g_vector[1][23] , \g_vector[1][21] ,
         \g_vector[1][19] , \g_vector[1][17] , \g_vector[1][15] ,
         \g_vector[1][13] , \g_vector[1][11] , \g_vector[1][9] ,
         \g_vector[1][7] , \g_vector[1][5] , \g_vector[1][3] ,
         \g_vector[1][1] , \g_vector[0][31] , \g_vector[0][30] ,
         \g_vector[0][29] , \g_vector[0][28] , \g_vector[0][27] ,
         \g_vector[0][26] , \g_vector[0][25] , \g_vector[0][24] ,
         \g_vector[0][23] , \g_vector[0][22] , \g_vector[0][21] ,
         \g_vector[0][20] , \g_vector[0][19] , \g_vector[0][18] ,
         \g_vector[0][17] , \g_vector[0][16] , \g_vector[0][15] ,
         \g_vector[0][14] , \g_vector[0][13] , \g_vector[0][12] ,
         \g_vector[0][11] , \g_vector[0][10] , \g_vector[0][9] ,
         \g_vector[0][8] , \g_vector[0][7] , \g_vector[0][6] ,
         \g_vector[0][5] , \g_vector[0][4] , \g_vector[0][3] ,
         \g_vector[0][2] , \g_vector[0][1] , \g_vector[0][0] ,
         \p_vector[4][31] , \p_vector[4][27] , \p_vector[3][31] ,
         \p_vector[3][23] , \p_vector[3][15] , \p_vector[2][31] ,
         \p_vector[2][27] , \p_vector[2][23] , \p_vector[2][19] ,
         \p_vector[2][15] , \p_vector[2][11] , \p_vector[2][7] ,
         \p_vector[1][31] , \p_vector[1][29] , \p_vector[1][27] ,
         \p_vector[1][25] , \p_vector[1][23] , \p_vector[1][21] ,
         \p_vector[1][19] , \p_vector[1][17] , \p_vector[1][15] ,
         \p_vector[1][13] , \p_vector[1][11] , \p_vector[1][9] ,
         \p_vector[1][7] , \p_vector[1][5] , \p_vector[1][3] ,
         \p_vector[0][31] , \p_vector[0][30] , \p_vector[0][29] ,
         \p_vector[0][28] , \p_vector[0][27] , \p_vector[0][26] ,
         \p_vector[0][25] , \p_vector[0][24] , \p_vector[0][23] ,
         \p_vector[0][22] , \p_vector[0][21] , \p_vector[0][20] ,
         \p_vector[0][19] , \p_vector[0][18] , \p_vector[0][17] ,
         \p_vector[0][16] , \p_vector[0][15] , \p_vector[0][14] ,
         \p_vector[0][13] , \p_vector[0][12] , \p_vector[0][11] ,
         \p_vector[0][10] , \p_vector[0][9] , \p_vector[0][8] ,
         \p_vector[0][7] , \p_vector[0][6] , \p_vector[0][5] ,
         \p_vector[0][4] , \p_vector[0][3] , \p_vector[0][2] ,
         \p_vector[0][1] , n3, n1, n2;

  pg_net_0 pg_network_31 ( .a(A[31]), .b(B[31]), .p(\p_vector[0][31] ), .g(
        \g_vector[0][31] ) );
  pg_net_250 pg_network_30 ( .a(A[30]), .b(B[30]), .p(\p_vector[0][30] ), .g(
        \g_vector[0][30] ) );
  pg_net_249 pg_network_29 ( .a(A[29]), .b(B[29]), .p(\p_vector[0][29] ), .g(
        \g_vector[0][29] ) );
  pg_net_248 pg_network_28 ( .a(A[28]), .b(B[28]), .p(\p_vector[0][28] ), .g(
        \g_vector[0][28] ) );
  pg_net_247 pg_network_27 ( .a(A[27]), .b(B[27]), .p(\p_vector[0][27] ), .g(
        \g_vector[0][27] ) );
  pg_net_246 pg_network_26 ( .a(A[26]), .b(B[26]), .p(\p_vector[0][26] ), .g(
        \g_vector[0][26] ) );
  pg_net_245 pg_network_25 ( .a(A[25]), .b(B[25]), .p(\p_vector[0][25] ), .g(
        \g_vector[0][25] ) );
  pg_net_244 pg_network_24 ( .a(A[24]), .b(B[24]), .p(\p_vector[0][24] ), .g(
        \g_vector[0][24] ) );
  pg_net_243 pg_network_23 ( .a(A[23]), .b(B[23]), .p(\p_vector[0][23] ), .g(
        \g_vector[0][23] ) );
  pg_net_242 pg_network_22 ( .a(A[22]), .b(B[22]), .p(\p_vector[0][22] ), .g(
        \g_vector[0][22] ) );
  pg_net_241 pg_network_21 ( .a(A[21]), .b(B[21]), .p(\p_vector[0][21] ), .g(
        \g_vector[0][21] ) );
  pg_net_240 pg_network_20 ( .a(A[20]), .b(B[20]), .p(\p_vector[0][20] ), .g(
        \g_vector[0][20] ) );
  pg_net_239 pg_network_19 ( .a(A[19]), .b(B[19]), .p(\p_vector[0][19] ), .g(
        \g_vector[0][19] ) );
  pg_net_238 pg_network_18 ( .a(A[18]), .b(B[18]), .p(\p_vector[0][18] ), .g(
        \g_vector[0][18] ) );
  pg_net_237 pg_network_17 ( .a(A[17]), .b(B[17]), .p(\p_vector[0][17] ), .g(
        \g_vector[0][17] ) );
  pg_net_236 pg_network_16 ( .a(A[16]), .b(B[16]), .p(\p_vector[0][16] ), .g(
        \g_vector[0][16] ) );
  pg_net_235 pg_network_15 ( .a(A[15]), .b(B[15]), .p(\p_vector[0][15] ), .g(
        \g_vector[0][15] ) );
  pg_net_234 pg_network_14 ( .a(A[14]), .b(B[14]), .p(\p_vector[0][14] ), .g(
        \g_vector[0][14] ) );
  pg_net_233 pg_network_13 ( .a(A[13]), .b(B[13]), .p(\p_vector[0][13] ), .g(
        \g_vector[0][13] ) );
  pg_net_232 pg_network_12 ( .a(A[12]), .b(B[12]), .p(\p_vector[0][12] ), .g(
        \g_vector[0][12] ) );
  pg_net_231 pg_network_11 ( .a(A[11]), .b(B[11]), .p(\p_vector[0][11] ), .g(
        \g_vector[0][11] ) );
  pg_net_230 pg_network_10 ( .a(A[10]), .b(B[10]), .p(\p_vector[0][10] ), .g(
        \g_vector[0][10] ) );
  pg_net_229 pg_network_9 ( .a(A[9]), .b(B[9]), .p(\p_vector[0][9] ), .g(
        \g_vector[0][9] ) );
  pg_net_228 pg_network_8 ( .a(A[8]), .b(B[8]), .p(\p_vector[0][8] ), .g(
        \g_vector[0][8] ) );
  pg_net_227 pg_network_7 ( .a(A[7]), .b(B[7]), .p(\p_vector[0][7] ), .g(
        \g_vector[0][7] ) );
  pg_net_226 pg_network_6 ( .a(A[6]), .b(B[6]), .p(\p_vector[0][6] ), .g(
        \g_vector[0][6] ) );
  pg_net_225 pg_network_5 ( .a(A[5]), .b(B[5]), .p(\p_vector[0][5] ), .g(
        \g_vector[0][5] ) );
  pg_net_224 pg_network_4 ( .a(A[4]), .b(B[4]), .p(\p_vector[0][4] ), .g(
        \g_vector[0][4] ) );
  pg_net_223 pg_network_3 ( .a(A[3]), .b(B[3]), .p(\p_vector[0][3] ), .g(
        \g_vector[0][3] ) );
  pg_net_222 pg_network_2 ( .a(A[2]), .b(B[2]), .p(\p_vector[0][2] ), .g(
        \g_vector[0][2] ) );
  pg_net_221 pg_network_1 ( .a(A[1]), .b(B[1]), .p(\p_vector[0][1] ), .g(
        \g_vector[0][1] ) );
  PG_BLOCK_0 std_PG_1_31 ( .p2(\p_vector[0][31] ), .g2(\g_vector[0][31] ), 
        .p1(\p_vector[0][30] ), .g1(\g_vector[0][30] ), .PG_P(
        \p_vector[1][31] ), .PG_G(\g_vector[1][31] ) );
  PG_BLOCK_242 std_PG_1_29 ( .p2(\p_vector[0][29] ), .g2(\g_vector[0][29] ), 
        .p1(\p_vector[0][28] ), .g1(\g_vector[0][28] ), .PG_P(
        \p_vector[1][29] ), .PG_G(\g_vector[1][29] ) );
  PG_BLOCK_241 std_PG_1_27 ( .p2(\p_vector[0][27] ), .g2(\g_vector[0][27] ), 
        .p1(\p_vector[0][26] ), .g1(\g_vector[0][26] ), .PG_P(
        \p_vector[1][27] ), .PG_G(\g_vector[1][27] ) );
  PG_BLOCK_240 std_PG_1_25 ( .p2(\p_vector[0][25] ), .g2(\g_vector[0][25] ), 
        .p1(\p_vector[0][24] ), .g1(\g_vector[0][24] ), .PG_P(
        \p_vector[1][25] ), .PG_G(\g_vector[1][25] ) );
  PG_BLOCK_239 std_PG_1_23 ( .p2(\p_vector[0][23] ), .g2(\g_vector[0][23] ), 
        .p1(\p_vector[0][22] ), .g1(\g_vector[0][22] ), .PG_P(
        \p_vector[1][23] ), .PG_G(\g_vector[1][23] ) );
  PG_BLOCK_238 std_PG_1_21 ( .p2(\p_vector[0][21] ), .g2(\g_vector[0][21] ), 
        .p1(\p_vector[0][20] ), .g1(\g_vector[0][20] ), .PG_P(
        \p_vector[1][21] ), .PG_G(\g_vector[1][21] ) );
  PG_BLOCK_237 std_PG_1_19 ( .p2(\p_vector[0][19] ), .g2(\g_vector[0][19] ), 
        .p1(\p_vector[0][18] ), .g1(\g_vector[0][18] ), .PG_P(
        \p_vector[1][19] ), .PG_G(\g_vector[1][19] ) );
  PG_BLOCK_236 std_PG_1_17 ( .p2(\p_vector[0][17] ), .g2(\g_vector[0][17] ), 
        .p1(\p_vector[0][16] ), .g1(\g_vector[0][16] ), .PG_P(
        \p_vector[1][17] ), .PG_G(\g_vector[1][17] ) );
  PG_BLOCK_235 std_PG_1_15 ( .p2(\p_vector[0][15] ), .g2(\g_vector[0][15] ), 
        .p1(\p_vector[0][14] ), .g1(\g_vector[0][14] ), .PG_P(
        \p_vector[1][15] ), .PG_G(\g_vector[1][15] ) );
  PG_BLOCK_234 std_PG_1_13 ( .p2(\p_vector[0][13] ), .g2(\g_vector[0][13] ), 
        .p1(\p_vector[0][12] ), .g1(\g_vector[0][12] ), .PG_P(
        \p_vector[1][13] ), .PG_G(\g_vector[1][13] ) );
  PG_BLOCK_233 std_PG_1_11 ( .p2(\p_vector[0][11] ), .g2(\g_vector[0][11] ), 
        .p1(\p_vector[0][10] ), .g1(\g_vector[0][10] ), .PG_P(
        \p_vector[1][11] ), .PG_G(\g_vector[1][11] ) );
  PG_BLOCK_232 std_PG_1_9 ( .p2(\p_vector[0][9] ), .g2(\g_vector[0][9] ), .p1(
        \p_vector[0][8] ), .g1(\g_vector[0][8] ), .PG_P(\p_vector[1][9] ), 
        .PG_G(\g_vector[1][9] ) );
  PG_BLOCK_231 std_PG_1_7 ( .p2(\p_vector[0][7] ), .g2(\g_vector[0][7] ), .p1(
        \p_vector[0][6] ), .g1(\g_vector[0][6] ), .PG_P(\p_vector[1][7] ), 
        .PG_G(\g_vector[1][7] ) );
  PG_BLOCK_230 std_PG_1_5 ( .p2(\p_vector[0][5] ), .g2(\g_vector[0][5] ), .p1(
        \p_vector[0][4] ), .g1(\g_vector[0][4] ), .PG_P(\p_vector[1][5] ), 
        .PG_G(\g_vector[1][5] ) );
  PG_BLOCK_229 std_PG_1_3 ( .p2(\p_vector[0][3] ), .g2(\g_vector[0][3] ), .p1(
        \p_vector[0][2] ), .g1(\g_vector[0][2] ), .PG_P(\p_vector[1][3] ), 
        .PG_G(\g_vector[1][3] ) );
  G_BLOCK_0 std_G_1_1 ( .p2(\p_vector[0][1] ), .g2(\g_vector[0][1] ), .g1(
        \g_vector[0][0] ), .G(\g_vector[1][1] ) );
  PG_BLOCK_228 std_PG_2_31 ( .p2(\p_vector[1][31] ), .g2(\g_vector[1][31] ), 
        .p1(\p_vector[1][29] ), .g1(\g_vector[1][29] ), .PG_P(
        \p_vector[2][31] ), .PG_G(\g_vector[2][31] ) );
  PG_BLOCK_227 std_PG_2_27 ( .p2(\p_vector[1][27] ), .g2(\g_vector[1][27] ), 
        .p1(\p_vector[1][25] ), .g1(\g_vector[1][25] ), .PG_P(
        \p_vector[2][27] ), .PG_G(\g_vector[2][27] ) );
  PG_BLOCK_226 std_PG_2_23 ( .p2(\p_vector[1][23] ), .g2(\g_vector[1][23] ), 
        .p1(\p_vector[1][21] ), .g1(\g_vector[1][21] ), .PG_P(
        \p_vector[2][23] ), .PG_G(\g_vector[2][23] ) );
  PG_BLOCK_225 std_PG_2_19 ( .p2(\p_vector[1][19] ), .g2(\g_vector[1][19] ), 
        .p1(\p_vector[1][17] ), .g1(\g_vector[1][17] ), .PG_P(
        \p_vector[2][19] ), .PG_G(\g_vector[2][19] ) );
  PG_BLOCK_224 std_PG_2_15 ( .p2(\p_vector[1][15] ), .g2(\g_vector[1][15] ), 
        .p1(\p_vector[1][13] ), .g1(\g_vector[1][13] ), .PG_P(
        \p_vector[2][15] ), .PG_G(\g_vector[2][15] ) );
  PG_BLOCK_223 std_PG_2_11 ( .p2(\p_vector[1][11] ), .g2(\g_vector[1][11] ), 
        .p1(\p_vector[1][9] ), .g1(\g_vector[1][9] ), .PG_P(\p_vector[2][11] ), 
        .PG_G(\g_vector[2][11] ) );
  PG_BLOCK_222 std_PG_2_7 ( .p2(\p_vector[1][7] ), .g2(\g_vector[1][7] ), .p1(
        \p_vector[1][5] ), .g1(\g_vector[1][5] ), .PG_P(\p_vector[2][7] ), 
        .PG_G(\g_vector[2][7] ) );
  G_BLOCK_68 std_G_2_3 ( .p2(\p_vector[1][3] ), .g2(\g_vector[1][3] ), .g1(
        \g_vector[1][1] ), .G(Co[0]) );
  PG_BLOCK_221 std_PG_3_31 ( .p2(\p_vector[2][31] ), .g2(\g_vector[2][31] ), 
        .p1(\p_vector[2][27] ), .g1(\g_vector[2][27] ), .PG_P(
        \p_vector[3][31] ), .PG_G(\g_vector[3][31] ) );
  PG_BLOCK_220 std_PG_3_23 ( .p2(\p_vector[2][23] ), .g2(\g_vector[2][23] ), 
        .p1(\p_vector[2][19] ), .g1(\g_vector[2][19] ), .PG_P(
        \p_vector[3][23] ), .PG_G(\g_vector[3][23] ) );
  PG_BLOCK_219 std_PG_3_15 ( .p2(\p_vector[2][15] ), .g2(\g_vector[2][15] ), 
        .p1(\p_vector[2][11] ), .g1(\g_vector[2][11] ), .PG_P(
        \p_vector[3][15] ), .PG_G(\g_vector[3][15] ) );
  G_BLOCK_67 std_G_3_7 ( .p2(\p_vector[2][7] ), .g2(\g_vector[2][7] ), .g1(
        Co[0]), .G(Co[1]) );
  PG_BLOCK_218 std_PG_4_31 ( .p2(\p_vector[3][31] ), .g2(\g_vector[3][31] ), 
        .p1(\p_vector[3][23] ), .g1(\g_vector[3][23] ), .PG_P(
        \p_vector[4][31] ), .PG_G(\g_vector[4][31] ) );
  PG_BLOCK_217 add_PG_4_31_1 ( .p2(\p_vector[2][27] ), .g2(\g_vector[2][27] ), 
        .p1(\p_vector[3][23] ), .g1(\g_vector[3][23] ), .PG_P(
        \p_vector[4][27] ), .PG_G(\g_vector[4][27] ) );
  G_BLOCK_66 std_G_4_15 ( .p2(\p_vector[3][15] ), .g2(\g_vector[3][15] ), .g1(
        Co[1]), .G(Co[3]) );
  G_BLOCK_65 add_G_4_15_1 ( .p2(\p_vector[2][11] ), .g2(\g_vector[2][11] ), 
        .g1(Co[1]), .G(Co[2]) );
  G_BLOCK_64 std_G_5_31 ( .p2(\p_vector[4][31] ), .g2(\g_vector[4][31] ), .g1(
        Co[3]), .G(Co[7]) );
  G_BLOCK_63 add_G_5_31_1 ( .p2(\p_vector[4][27] ), .g2(\g_vector[4][27] ), 
        .g1(Co[3]), .G(Co[6]) );
  G_BLOCK_62 add_G_5_31_2 ( .p2(\p_vector[3][23] ), .g2(\g_vector[3][23] ), 
        .g1(Co[3]), .G(Co[5]) );
  G_BLOCK_61 add_G_5_31_3 ( .p2(\p_vector[2][19] ), .g2(\g_vector[2][19] ), 
        .g1(Co[3]), .G(Co[4]) );
  INV_X1 U1 ( .A(B[0]), .ZN(n2) );
  OAI21_X1 U2 ( .B1(n1), .B2(n2), .A(n3), .ZN(\g_vector[0][0] ) );
  OAI21_X1 U3 ( .B1(A[0]), .B2(B[0]), .A(Cin), .ZN(n3) );
  INV_X1 U4 ( .A(A[0]), .ZN(n1) );
endmodule


module FA_0 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_511 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_510 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_509 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_0 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_0 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_511 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_510 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_509 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_508 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_507 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_506 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_505 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_127 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_508 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_507 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_506 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_505 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_392 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_391 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_390 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_389 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_GENERIC_NBIT4_0 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_392 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_391 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_390 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_389 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_0 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_0 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_127 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_0 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module FA_504 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_503 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_502 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_501 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_126 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_504 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_503 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_502 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_501 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_500 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_499 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_498 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_497 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_125 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_500 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_499 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_498 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_497 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_388 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_387 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  AOI22_X1 U1 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U2 ( .A(S), .ZN(n2) );
  INV_X1 U3 ( .A(n4), .ZN(Y) );
endmodule


module MUX21_386 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  AOI22_X1 U1 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U2 ( .A(S), .ZN(n2) );
  INV_X1 U3 ( .A(n4), .ZN(Y) );
endmodule


module MUX21_385 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_GENERIC_NBIT4_63 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_388 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_387 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_386 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_385 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_63 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_126 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_125 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_63 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module FA_496 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_495 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_494 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_493 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_124 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_496 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_495 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_494 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_493 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_492 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_491 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_490 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_489 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_123 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_492 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_491 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_490 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_489 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_384 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_383 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_382 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_381 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_GENERIC_NBIT4_62 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_384 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_383 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_382 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_381 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_62 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_124 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_123 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_62 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module FA_488 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_487 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_486 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_485 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_122 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_488 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_487 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_486 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_485 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_484 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_483 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_482 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_481 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_121 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_484 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_483 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_482 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_481 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_380 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_379 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_378 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_377 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  AOI22_X1 U1 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U2 ( .A(S), .ZN(n2) );
  INV_X1 U3 ( .A(n4), .ZN(Y) );
endmodule


module MUX21_GENERIC_NBIT4_61 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_380 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_379 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_378 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_377 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_61 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_122 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_121 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_61 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module FA_480 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_479 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_478 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_477 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_120 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_480 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_479 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_478 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_477 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_476 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_475 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_474 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_473 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_119 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_476 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_475 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_474 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_473 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_376 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_375 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  AOI22_X1 U1 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U2 ( .A(S), .ZN(n2) );
  INV_X1 U3 ( .A(n4), .ZN(Y) );
endmodule


module MUX21_374 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  AOI22_X1 U1 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U2 ( .A(S), .ZN(n2) );
  INV_X1 U3 ( .A(n4), .ZN(Y) );
endmodule


module MUX21_373 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  AOI22_X1 U1 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U2 ( .A(S), .ZN(n2) );
  INV_X1 U3 ( .A(n4), .ZN(Y) );
endmodule


module MUX21_GENERIC_NBIT4_60 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_376 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_375 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_374 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_373 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_60 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_120 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_119 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_60 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module FA_472 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_471 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_470 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_469 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_118 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_472 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_471 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_470 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_469 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_468 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_467 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_466 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_465 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_117 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_468 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_467 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_466 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_465 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_372 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_371 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  AOI22_X1 U1 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U2 ( .A(S), .ZN(n2) );
  INV_X1 U3 ( .A(n4), .ZN(Y) );
endmodule


module MUX21_370 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  AOI22_X1 U1 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U2 ( .A(S), .ZN(n2) );
  INV_X1 U3 ( .A(n4), .ZN(Y) );
endmodule


module MUX21_369 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  AOI22_X1 U1 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U2 ( .A(S), .ZN(n2) );
  INV_X1 U3 ( .A(n4), .ZN(Y) );
endmodule


module MUX21_GENERIC_NBIT4_59 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_372 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_371 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_370 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_369 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_59 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_118 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_117 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_59 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module FA_464 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_463 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_462 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_461 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_116 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_464 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_463 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_462 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_461 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_460 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_459 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_458 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_457 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_115 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_460 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_459 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_458 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_457 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_368 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_367 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  AOI22_X1 U1 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U2 ( .A(S), .ZN(n2) );
  INV_X1 U3 ( .A(n4), .ZN(Y) );
endmodule


module MUX21_366 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  AOI22_X1 U1 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U2 ( .A(S), .ZN(n2) );
  INV_X1 U3 ( .A(n4), .ZN(Y) );
endmodule


module MUX21_365 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  AOI22_X1 U1 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U2 ( .A(S), .ZN(n2) );
  INV_X1 U3 ( .A(n4), .ZN(Y) );
endmodule


module MUX21_GENERIC_NBIT4_58 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_368 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_367 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_366 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_365 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_58 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_116 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_115 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_58 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module FA_456 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_455 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_454 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_453 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_114 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_456 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_455 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_454 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_453 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_452 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_451 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_450 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_449 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_113 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_452 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_451 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_450 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_449 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_364 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_363 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  AOI22_X1 U1 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U2 ( .A(S), .ZN(n2) );
  INV_X1 U3 ( .A(n4), .ZN(Y) );
endmodule


module MUX21_362 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  AOI22_X1 U1 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U2 ( .A(S), .ZN(n2) );
  INV_X1 U3 ( .A(n4), .ZN(Y) );
endmodule


module MUX21_361 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_GENERIC_NBIT4_57 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_364 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_363 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_362 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_361 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_57 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_114 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_113 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_57 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module sum_generator_n_bit32_n_CSB8_0 ( A, B, C_in, S );
  input [31:0] A;
  input [31:0] B;
  input [7:0] C_in;
  output [31:0] S;


  carry_select_block_n4_0 csb_0 ( .A(A[3:0]), .B(B[3:0]), .C_sel(C_in[0]), .S(
        S[3:0]) );
  carry_select_block_n4_63 csb_1 ( .A(A[7:4]), .B(B[7:4]), .C_sel(C_in[1]), 
        .S(S[7:4]) );
  carry_select_block_n4_62 csb_2 ( .A(A[11:8]), .B(B[11:8]), .C_sel(C_in[2]), 
        .S(S[11:8]) );
  carry_select_block_n4_61 csb_3 ( .A(A[15:12]), .B(B[15:12]), .C_sel(C_in[3]), 
        .S(S[15:12]) );
  carry_select_block_n4_60 csb_4 ( .A(A[19:16]), .B(B[19:16]), .C_sel(C_in[4]), 
        .S(S[19:16]) );
  carry_select_block_n4_59 csb_5 ( .A(A[23:20]), .B(B[23:20]), .C_sel(C_in[5]), 
        .S(S[23:20]) );
  carry_select_block_n4_58 csb_6 ( .A(A[27:24]), .B(B[27:24]), .C_sel(C_in[6]), 
        .S(S[27:24]) );
  carry_select_block_n4_57 csb_7 ( .A(A[31:28]), .B(B[31:28]), .C_sel(C_in[7]), 
        .S(S[31:28]) );
endmodule


module P4_ADDER_NBIT32_0 ( A, B, Cin, S, Cout, ovf );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Cin;
  output Cout, ovf;
  wire   n1, n2;
  wire   [31:0] xor_b;
  wire   [6:0] carry;

  XOR2_X1 U3 ( .A(xor_b[31]), .B(A[31]), .Z(n2) );
  my_xor_0 bc_xor_31 ( .A(B[31]), .B(Cin), .xor_out(xor_b[31]) );
  my_xor_255 bc_xor_30 ( .A(B[30]), .B(Cin), .xor_out(xor_b[30]) );
  my_xor_254 bc_xor_29 ( .A(B[29]), .B(Cin), .xor_out(xor_b[29]) );
  my_xor_253 bc_xor_28 ( .A(B[28]), .B(Cin), .xor_out(xor_b[28]) );
  my_xor_252 bc_xor_27 ( .A(B[27]), .B(Cin), .xor_out(xor_b[27]) );
  my_xor_251 bc_xor_26 ( .A(B[26]), .B(Cin), .xor_out(xor_b[26]) );
  my_xor_250 bc_xor_25 ( .A(B[25]), .B(Cin), .xor_out(xor_b[25]) );
  my_xor_249 bc_xor_24 ( .A(B[24]), .B(Cin), .xor_out(xor_b[24]) );
  my_xor_248 bc_xor_23 ( .A(B[23]), .B(Cin), .xor_out(xor_b[23]) );
  my_xor_247 bc_xor_22 ( .A(B[22]), .B(Cin), .xor_out(xor_b[22]) );
  my_xor_246 bc_xor_21 ( .A(B[21]), .B(Cin), .xor_out(xor_b[21]) );
  my_xor_245 bc_xor_20 ( .A(B[20]), .B(Cin), .xor_out(xor_b[20]) );
  my_xor_244 bc_xor_19 ( .A(B[19]), .B(Cin), .xor_out(xor_b[19]) );
  my_xor_243 bc_xor_18 ( .A(B[18]), .B(Cin), .xor_out(xor_b[18]) );
  my_xor_242 bc_xor_17 ( .A(B[17]), .B(Cin), .xor_out(xor_b[17]) );
  my_xor_241 bc_xor_16 ( .A(B[16]), .B(Cin), .xor_out(xor_b[16]) );
  my_xor_240 bc_xor_15 ( .A(B[15]), .B(Cin), .xor_out(xor_b[15]) );
  my_xor_239 bc_xor_14 ( .A(B[14]), .B(Cin), .xor_out(xor_b[14]) );
  my_xor_238 bc_xor_13 ( .A(B[13]), .B(Cin), .xor_out(xor_b[13]) );
  my_xor_237 bc_xor_12 ( .A(B[12]), .B(Cin), .xor_out(xor_b[12]) );
  my_xor_236 bc_xor_11 ( .A(B[11]), .B(Cin), .xor_out(xor_b[11]) );
  my_xor_235 bc_xor_10 ( .A(B[10]), .B(Cin), .xor_out(xor_b[10]) );
  my_xor_234 bc_xor_9 ( .A(B[9]), .B(Cin), .xor_out(xor_b[9]) );
  my_xor_233 bc_xor_8 ( .A(B[8]), .B(Cin), .xor_out(xor_b[8]) );
  my_xor_232 bc_xor_7 ( .A(B[7]), .B(Cin), .xor_out(xor_b[7]) );
  my_xor_231 bc_xor_6 ( .A(B[6]), .B(Cin), .xor_out(xor_b[6]) );
  my_xor_230 bc_xor_5 ( .A(B[5]), .B(Cin), .xor_out(xor_b[5]) );
  my_xor_229 bc_xor_4 ( .A(B[4]), .B(Cin), .xor_out(xor_b[4]) );
  my_xor_228 bc_xor_3 ( .A(B[3]), .B(Cin), .xor_out(xor_b[3]) );
  my_xor_227 bc_xor_2 ( .A(B[2]), .B(Cin), .xor_out(xor_b[2]) );
  my_xor_226 bc_xor_1 ( .A(B[1]), .B(Cin), .xor_out(xor_b[1]) );
  my_xor_225 bc_xor_0 ( .A(B[0]), .B(Cin), .xor_out(xor_b[0]) );
  CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_0 CG ( .A(A), .B(xor_b), .Cin(Cin), 
        .Co({Cout, carry}) );
  sum_generator_n_bit32_n_CSB8_0 SG ( .A(A), .B(xor_b), .C_in({carry, Cin}), 
        .S(S) );
  NOR2_X1 U1 ( .A1(n1), .A2(n2), .ZN(ovf) );
  XNOR2_X1 U2 ( .A(A[31]), .B(S[31]), .ZN(n1) );
endmodule


module jump_logic_WORD_size32_NREG32_reg_file_size32 ( opcode, RSA, WB_RD, 
        MEM_RD, Rega, ALU_out, MEM_out, Rega_new, mux_s, flag );
  input [5:0] opcode;
  input [4:0] RSA;
  input [4:0] WB_RD;
  input [4:0] MEM_RD;
  input [31:0] Rega;
  input [31:0] ALU_out;
  input [31:0] MEM_out;
  output [31:0] Rega_new;
  output mux_s, flag;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76;

  BUF_X1 U3 ( .A(n11), .Z(n1) );
  BUF_X1 U4 ( .A(n11), .Z(n2) );
  BUF_X1 U5 ( .A(n11), .Z(n3) );
  BUF_X1 U6 ( .A(n12), .Z(n5) );
  BUF_X1 U7 ( .A(n12), .Z(n4) );
  BUF_X1 U8 ( .A(n13), .Z(n8) );
  BUF_X1 U9 ( .A(n13), .Z(n7) );
  BUF_X1 U10 ( .A(n12), .Z(n6) );
  BUF_X1 U11 ( .A(n13), .Z(n9) );
  INV_X1 U12 ( .A(n10), .ZN(Rega_new[31]) );
  AOI222_X1 U13 ( .A1(ALU_out[31]), .A2(n1), .B1(MEM_out[31]), .B2(n6), .C1(
        Rega[31]), .C2(n9), .ZN(n10) );
  INV_X1 U14 ( .A(n14), .ZN(Rega_new[30]) );
  INV_X1 U15 ( .A(n15), .ZN(Rega_new[29]) );
  INV_X1 U16 ( .A(n16), .ZN(Rega_new[28]) );
  INV_X1 U17 ( .A(n17), .ZN(Rega_new[27]) );
  INV_X1 U18 ( .A(n18), .ZN(Rega_new[26]) );
  INV_X1 U19 ( .A(n19), .ZN(Rega_new[25]) );
  INV_X1 U20 ( .A(n20), .ZN(Rega_new[24]) );
  INV_X1 U21 ( .A(n21), .ZN(Rega_new[23]) );
  INV_X1 U22 ( .A(n22), .ZN(Rega_new[22]) );
  INV_X1 U23 ( .A(n23), .ZN(Rega_new[21]) );
  INV_X1 U24 ( .A(n24), .ZN(Rega_new[20]) );
  INV_X1 U25 ( .A(n25), .ZN(Rega_new[19]) );
  INV_X1 U26 ( .A(n26), .ZN(Rega_new[18]) );
  INV_X1 U27 ( .A(n27), .ZN(Rega_new[17]) );
  INV_X1 U28 ( .A(n28), .ZN(Rega_new[16]) );
  INV_X1 U29 ( .A(n29), .ZN(Rega_new[15]) );
  INV_X1 U30 ( .A(n30), .ZN(Rega_new[6]) );
  INV_X1 U31 ( .A(n31), .ZN(Rega_new[5]) );
  INV_X1 U32 ( .A(n32), .ZN(Rega_new[4]) );
  INV_X1 U33 ( .A(n33), .ZN(Rega_new[3]) );
  AND4_X1 U34 ( .A1(n34), .A2(n35), .A3(opcode[1]), .A4(opcode[4]), .ZN(mux_s)
         );
  OAI22_X1 U35 ( .A1(n36), .A2(n37), .B1(n38), .B2(n39), .ZN(flag) );
  INV_X1 U36 ( .A(n35), .ZN(n39) );
  AOI22_X1 U37 ( .A1(n40), .A2(n41), .B1(opcode[1]), .B2(n34), .ZN(n38) );
  AND2_X1 U38 ( .A1(n37), .A2(n36), .ZN(n40) );
  NAND3_X1 U39 ( .A1(n42), .A2(n35), .A3(n41), .ZN(n37) );
  NOR3_X1 U40 ( .A1(opcode[1]), .A2(opcode[4]), .A3(n34), .ZN(n41) );
  INV_X1 U41 ( .A(opcode[2]), .ZN(n34) );
  NOR2_X1 U42 ( .A1(opcode[5]), .A2(opcode[3]), .ZN(n35) );
  INV_X1 U43 ( .A(opcode[0]), .ZN(n42) );
  NAND4_X1 U44 ( .A1(n43), .A2(n44), .A3(n45), .A4(n46), .ZN(n36) );
  NOR4_X1 U45 ( .A1(n47), .A2(n48), .A3(n49), .A4(n50), .ZN(n46) );
  NAND4_X1 U46 ( .A1(n29), .A2(n28), .A3(n27), .A4(n26), .ZN(n50) );
  AOI222_X1 U47 ( .A1(ALU_out[18]), .A2(n1), .B1(MEM_out[18]), .B2(n6), .C1(
        Rega[18]), .C2(n9), .ZN(n26) );
  AOI222_X1 U48 ( .A1(ALU_out[17]), .A2(n1), .B1(MEM_out[17]), .B2(n6), .C1(
        Rega[17]), .C2(n9), .ZN(n27) );
  AOI222_X1 U49 ( .A1(ALU_out[16]), .A2(n1), .B1(MEM_out[16]), .B2(n6), .C1(
        Rega[16]), .C2(n9), .ZN(n28) );
  AOI222_X1 U50 ( .A1(ALU_out[15]), .A2(n1), .B1(MEM_out[15]), .B2(n6), .C1(
        Rega[15]), .C2(n9), .ZN(n29) );
  NAND4_X1 U51 ( .A1(n25), .A2(n24), .A3(n23), .A4(n22), .ZN(n49) );
  AOI222_X1 U52 ( .A1(ALU_out[22]), .A2(n1), .B1(MEM_out[22]), .B2(n6), .C1(
        Rega[22]), .C2(n9), .ZN(n22) );
  AOI222_X1 U53 ( .A1(ALU_out[21]), .A2(n1), .B1(MEM_out[21]), .B2(n6), .C1(
        Rega[21]), .C2(n9), .ZN(n23) );
  AOI222_X1 U54 ( .A1(ALU_out[20]), .A2(n1), .B1(MEM_out[20]), .B2(n6), .C1(
        Rega[20]), .C2(n9), .ZN(n24) );
  AOI222_X1 U55 ( .A1(ALU_out[19]), .A2(n1), .B1(MEM_out[19]), .B2(n6), .C1(
        Rega[19]), .C2(n9), .ZN(n25) );
  NAND4_X1 U56 ( .A1(n21), .A2(n20), .A3(n19), .A4(n18), .ZN(n48) );
  AOI222_X1 U57 ( .A1(ALU_out[26]), .A2(n1), .B1(MEM_out[26]), .B2(n6), .C1(
        Rega[26]), .C2(n9), .ZN(n18) );
  AOI222_X1 U58 ( .A1(ALU_out[25]), .A2(n1), .B1(MEM_out[25]), .B2(n5), .C1(
        Rega[25]), .C2(n8), .ZN(n19) );
  AOI222_X1 U59 ( .A1(ALU_out[24]), .A2(n2), .B1(MEM_out[24]), .B2(n5), .C1(
        Rega[24]), .C2(n8), .ZN(n20) );
  AOI222_X1 U60 ( .A1(ALU_out[23]), .A2(n2), .B1(MEM_out[23]), .B2(n5), .C1(
        Rega[23]), .C2(n8), .ZN(n21) );
  NAND4_X1 U61 ( .A1(n17), .A2(n16), .A3(n15), .A4(n14), .ZN(n47) );
  AOI222_X1 U62 ( .A1(ALU_out[30]), .A2(n2), .B1(MEM_out[30]), .B2(n5), .C1(
        Rega[30]), .C2(n8), .ZN(n14) );
  AOI222_X1 U63 ( .A1(ALU_out[29]), .A2(n2), .B1(MEM_out[29]), .B2(n5), .C1(
        Rega[29]), .C2(n8), .ZN(n15) );
  AOI222_X1 U64 ( .A1(ALU_out[28]), .A2(n2), .B1(MEM_out[28]), .B2(n5), .C1(
        Rega[28]), .C2(n8), .ZN(n16) );
  AOI222_X1 U65 ( .A1(ALU_out[27]), .A2(n2), .B1(MEM_out[27]), .B2(n5), .C1(
        Rega[27]), .C2(n8), .ZN(n17) );
  NOR4_X1 U66 ( .A1(n51), .A2(Rega_new[0]), .A3(Rega_new[2]), .A4(Rega_new[1]), 
        .ZN(n45) );
  INV_X1 U67 ( .A(n52), .ZN(Rega_new[1]) );
  AOI222_X1 U68 ( .A1(ALU_out[1]), .A2(n2), .B1(MEM_out[1]), .B2(n5), .C1(
        Rega[1]), .C2(n8), .ZN(n52) );
  INV_X1 U69 ( .A(n53), .ZN(Rega_new[2]) );
  AOI222_X1 U70 ( .A1(ALU_out[2]), .A2(n2), .B1(MEM_out[2]), .B2(n5), .C1(
        Rega[2]), .C2(n8), .ZN(n53) );
  INV_X1 U71 ( .A(n54), .ZN(Rega_new[0]) );
  AOI222_X1 U72 ( .A1(ALU_out[0]), .A2(n2), .B1(MEM_out[0]), .B2(n5), .C1(
        Rega[0]), .C2(n8), .ZN(n54) );
  NAND4_X1 U73 ( .A1(n33), .A2(n32), .A3(n31), .A4(n30), .ZN(n51) );
  AOI222_X1 U74 ( .A1(ALU_out[6]), .A2(n2), .B1(MEM_out[6]), .B2(n5), .C1(
        Rega[6]), .C2(n8), .ZN(n30) );
  AOI222_X1 U75 ( .A1(ALU_out[5]), .A2(n2), .B1(MEM_out[5]), .B2(n4), .C1(
        Rega[5]), .C2(n7), .ZN(n31) );
  AOI222_X1 U76 ( .A1(ALU_out[4]), .A2(n3), .B1(MEM_out[4]), .B2(n4), .C1(
        Rega[4]), .C2(n7), .ZN(n32) );
  AOI222_X1 U77 ( .A1(ALU_out[3]), .A2(n3), .B1(MEM_out[3]), .B2(n4), .C1(
        Rega[3]), .C2(n7), .ZN(n33) );
  NOR4_X1 U78 ( .A1(Rega_new[14]), .A2(Rega_new[13]), .A3(Rega_new[12]), .A4(
        Rega_new[11]), .ZN(n44) );
  INV_X1 U79 ( .A(n55), .ZN(Rega_new[11]) );
  AOI222_X1 U80 ( .A1(ALU_out[11]), .A2(n3), .B1(MEM_out[11]), .B2(n4), .C1(
        Rega[11]), .C2(n7), .ZN(n55) );
  INV_X1 U81 ( .A(n56), .ZN(Rega_new[12]) );
  AOI222_X1 U82 ( .A1(ALU_out[12]), .A2(n3), .B1(MEM_out[12]), .B2(n4), .C1(
        Rega[12]), .C2(n7), .ZN(n56) );
  INV_X1 U83 ( .A(n57), .ZN(Rega_new[13]) );
  AOI222_X1 U84 ( .A1(ALU_out[13]), .A2(n3), .B1(MEM_out[13]), .B2(n4), .C1(
        Rega[13]), .C2(n7), .ZN(n57) );
  INV_X1 U85 ( .A(n58), .ZN(Rega_new[14]) );
  AOI222_X1 U86 ( .A1(ALU_out[14]), .A2(n3), .B1(MEM_out[14]), .B2(n4), .C1(
        Rega[14]), .C2(n7), .ZN(n58) );
  NOR4_X1 U87 ( .A1(Rega_new[10]), .A2(Rega_new[9]), .A3(Rega_new[8]), .A4(
        Rega_new[7]), .ZN(n43) );
  INV_X1 U88 ( .A(n59), .ZN(Rega_new[7]) );
  AOI222_X1 U89 ( .A1(ALU_out[7]), .A2(n3), .B1(MEM_out[7]), .B2(n4), .C1(
        Rega[7]), .C2(n7), .ZN(n59) );
  INV_X1 U90 ( .A(n60), .ZN(Rega_new[8]) );
  AOI222_X1 U91 ( .A1(ALU_out[8]), .A2(n3), .B1(MEM_out[8]), .B2(n4), .C1(
        Rega[8]), .C2(n7), .ZN(n60) );
  INV_X1 U92 ( .A(n61), .ZN(Rega_new[9]) );
  AOI222_X1 U93 ( .A1(ALU_out[9]), .A2(n3), .B1(MEM_out[9]), .B2(n4), .C1(
        Rega[9]), .C2(n7), .ZN(n61) );
  INV_X1 U94 ( .A(n62), .ZN(Rega_new[10]) );
  AOI222_X1 U95 ( .A1(ALU_out[10]), .A2(n3), .B1(MEM_out[10]), .B2(n4), .C1(
        Rega[10]), .C2(n7), .ZN(n62) );
  AND2_X1 U96 ( .A1(n63), .A2(n64), .ZN(n13) );
  NOR2_X1 U97 ( .A1(n63), .A2(n3), .ZN(n12) );
  NAND4_X1 U98 ( .A1(n65), .A2(n66), .A3(n67), .A4(n68), .ZN(n63) );
  NOR2_X1 U99 ( .A1(n69), .A2(n70), .ZN(n68) );
  XOR2_X1 U100 ( .A(WB_RD[4]), .B(RSA[4]), .Z(n70) );
  XOR2_X1 U101 ( .A(WB_RD[2]), .B(RSA[2]), .Z(n69) );
  XNOR2_X1 U102 ( .A(RSA[0]), .B(WB_RD[0]), .ZN(n67) );
  XNOR2_X1 U103 ( .A(RSA[1]), .B(WB_RD[1]), .ZN(n66) );
  XNOR2_X1 U104 ( .A(RSA[3]), .B(WB_RD[3]), .ZN(n65) );
  INV_X1 U105 ( .A(n64), .ZN(n11) );
  NAND3_X1 U106 ( .A1(n71), .A2(n72), .A3(n73), .ZN(n64) );
  NOR3_X1 U107 ( .A1(n74), .A2(n75), .A3(n76), .ZN(n73) );
  XOR2_X1 U108 ( .A(RSA[3]), .B(MEM_RD[3]), .Z(n76) );
  XOR2_X1 U109 ( .A(RSA[1]), .B(MEM_RD[1]), .Z(n75) );
  XOR2_X1 U110 ( .A(RSA[0]), .B(MEM_RD[0]), .Z(n74) );
  XNOR2_X1 U111 ( .A(RSA[2]), .B(MEM_RD[2]), .ZN(n72) );
  XNOR2_X1 U112 ( .A(RSA[4]), .B(MEM_RD[4]), .ZN(n71) );
endmodule


module MUX21_498 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_497 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_496 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_495 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_494 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_493 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_492 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_491 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_490 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_489 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_488 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_487 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_486 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_485 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_484 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_483 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_482 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_481 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_480 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_479 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_478 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_477 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_476 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_475 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_474 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_473 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_472 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_471 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_470 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_469 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_468 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_467 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_GENERIC_NBIT32_3 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   n1, n2, n3;

  MUX21_498 MUXES_0 ( .A(A[0]), .B(B[0]), .S(n1), .Y(Y[0]) );
  MUX21_497 MUXES_1 ( .A(A[1]), .B(B[1]), .S(n1), .Y(Y[1]) );
  MUX21_496 MUXES_2 ( .A(A[2]), .B(B[2]), .S(n1), .Y(Y[2]) );
  MUX21_495 MUXES_3 ( .A(A[3]), .B(B[3]), .S(n1), .Y(Y[3]) );
  MUX21_494 MUXES_4 ( .A(A[4]), .B(B[4]), .S(n1), .Y(Y[4]) );
  MUX21_493 MUXES_5 ( .A(A[5]), .B(B[5]), .S(n1), .Y(Y[5]) );
  MUX21_492 MUXES_6 ( .A(A[6]), .B(B[6]), .S(n1), .Y(Y[6]) );
  MUX21_491 MUXES_7 ( .A(A[7]), .B(B[7]), .S(n1), .Y(Y[7]) );
  MUX21_490 MUXES_8 ( .A(A[8]), .B(B[8]), .S(n1), .Y(Y[8]) );
  MUX21_489 MUXES_9 ( .A(A[9]), .B(B[9]), .S(n1), .Y(Y[9]) );
  MUX21_488 MUXES_10 ( .A(A[10]), .B(B[10]), .S(n1), .Y(Y[10]) );
  MUX21_487 MUXES_11 ( .A(A[11]), .B(B[11]), .S(n1), .Y(Y[11]) );
  MUX21_486 MUXES_12 ( .A(A[12]), .B(B[12]), .S(n2), .Y(Y[12]) );
  MUX21_485 MUXES_13 ( .A(A[13]), .B(B[13]), .S(n2), .Y(Y[13]) );
  MUX21_484 MUXES_14 ( .A(A[14]), .B(B[14]), .S(n2), .Y(Y[14]) );
  MUX21_483 MUXES_15 ( .A(A[15]), .B(B[15]), .S(n2), .Y(Y[15]) );
  MUX21_482 MUXES_16 ( .A(A[16]), .B(B[16]), .S(n2), .Y(Y[16]) );
  MUX21_481 MUXES_17 ( .A(A[17]), .B(B[17]), .S(n2), .Y(Y[17]) );
  MUX21_480 MUXES_18 ( .A(A[18]), .B(B[18]), .S(n2), .Y(Y[18]) );
  MUX21_479 MUXES_19 ( .A(A[19]), .B(B[19]), .S(n2), .Y(Y[19]) );
  MUX21_478 MUXES_20 ( .A(A[20]), .B(B[20]), .S(n2), .Y(Y[20]) );
  MUX21_477 MUXES_21 ( .A(A[21]), .B(B[21]), .S(n2), .Y(Y[21]) );
  MUX21_476 MUXES_22 ( .A(A[22]), .B(B[22]), .S(n2), .Y(Y[22]) );
  MUX21_475 MUXES_23 ( .A(A[23]), .B(B[23]), .S(n2), .Y(Y[23]) );
  MUX21_474 MUXES_24 ( .A(A[24]), .B(B[24]), .S(n3), .Y(Y[24]) );
  MUX21_473 MUXES_25 ( .A(A[25]), .B(B[25]), .S(n3), .Y(Y[25]) );
  MUX21_472 MUXES_26 ( .A(A[26]), .B(B[26]), .S(n3), .Y(Y[26]) );
  MUX21_471 MUXES_27 ( .A(A[27]), .B(B[27]), .S(n3), .Y(Y[27]) );
  MUX21_470 MUXES_28 ( .A(A[28]), .B(B[28]), .S(n3), .Y(Y[28]) );
  MUX21_469 MUXES_29 ( .A(A[29]), .B(B[29]), .S(n3), .Y(Y[29]) );
  MUX21_468 MUXES_30 ( .A(A[30]), .B(B[30]), .S(n3), .Y(Y[30]) );
  MUX21_467 MUXES_31 ( .A(A[31]), .B(B[31]), .S(n3), .Y(Y[31]) );
  BUF_X1 U1 ( .A(SEL), .Z(n2) );
  BUF_X1 U2 ( .A(SEL), .Z(n1) );
  BUF_X1 U3 ( .A(SEL), .Z(n3) );
endmodule



    module stall_detection_unit_op_code_size6_func_size11_PC_reg_size32_reg_file_size32_DW01_sub_0 ( 
        A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   \A[0] , n1, n2, n3;
  wire   [32:0] carry;
  assign DIFF[1] = A[1];
  assign DIFF[0] = \A[0] ;
  assign \A[0]  = A[0];

  XNOR2_X1 U1 ( .A(A[10]), .B(carry[10]), .ZN(DIFF[10]) );
  XNOR2_X1 U2 ( .A(A[11]), .B(carry[11]), .ZN(DIFF[11]) );
  XNOR2_X1 U3 ( .A(A[13]), .B(carry[13]), .ZN(DIFF[13]) );
  XNOR2_X1 U4 ( .A(A[15]), .B(carry[15]), .ZN(DIFF[15]) );
  XNOR2_X1 U5 ( .A(A[16]), .B(carry[16]), .ZN(DIFF[16]) );
  XNOR2_X1 U6 ( .A(A[17]), .B(carry[17]), .ZN(DIFF[17]) );
  XNOR2_X1 U7 ( .A(A[18]), .B(carry[18]), .ZN(DIFF[18]) );
  XNOR2_X1 U8 ( .A(A[19]), .B(carry[19]), .ZN(DIFF[19]) );
  XNOR2_X1 U9 ( .A(A[5]), .B(carry[5]), .ZN(DIFF[5]) );
  XNOR2_X1 U10 ( .A(A[8]), .B(carry[8]), .ZN(DIFF[8]) );
  XNOR2_X1 U11 ( .A(A[9]), .B(carry[9]), .ZN(DIFF[9]) );
  XNOR2_X1 U12 ( .A(A[20]), .B(carry[20]), .ZN(DIFF[20]) );
  XNOR2_X1 U13 ( .A(A[21]), .B(carry[21]), .ZN(DIFF[21]) );
  XNOR2_X1 U14 ( .A(A[22]), .B(carry[22]), .ZN(DIFF[22]) );
  XNOR2_X1 U15 ( .A(A[23]), .B(carry[23]), .ZN(DIFF[23]) );
  XNOR2_X1 U16 ( .A(A[24]), .B(carry[24]), .ZN(DIFF[24]) );
  XNOR2_X1 U17 ( .A(A[25]), .B(carry[25]), .ZN(DIFF[25]) );
  XNOR2_X1 U18 ( .A(A[26]), .B(carry[26]), .ZN(DIFF[26]) );
  XNOR2_X1 U19 ( .A(A[27]), .B(carry[27]), .ZN(DIFF[27]) );
  XNOR2_X1 U20 ( .A(A[28]), .B(carry[28]), .ZN(DIFF[28]) );
  XNOR2_X1 U21 ( .A(A[29]), .B(carry[29]), .ZN(DIFF[29]) );
  XNOR2_X1 U22 ( .A(A[30]), .B(carry[30]), .ZN(DIFF[30]) );
  XNOR2_X1 U23 ( .A(A[7]), .B(carry[7]), .ZN(DIFF[7]) );
  XNOR2_X1 U24 ( .A(n3), .B(A[2]), .ZN(DIFF[2]) );
  XNOR2_X1 U25 ( .A(A[3]), .B(carry[3]), .ZN(DIFF[3]) );
  XNOR2_X1 U26 ( .A(A[4]), .B(carry[4]), .ZN(DIFF[4]) );
  XNOR2_X1 U27 ( .A(A[12]), .B(carry[12]), .ZN(DIFF[12]) );
  XNOR2_X1 U28 ( .A(A[14]), .B(carry[14]), .ZN(DIFF[14]) );
  XNOR2_X1 U29 ( .A(A[6]), .B(carry[6]), .ZN(DIFF[6]) );
  XNOR2_X1 U30 ( .A(A[31]), .B(carry[31]), .ZN(DIFF[31]) );
  NAND2_X1 U31 ( .A1(n1), .A2(n2), .ZN(carry[31]) );
  INV_X1 U32 ( .A(A[30]), .ZN(n1) );
  INV_X1 U33 ( .A(carry[30]), .ZN(n2) );
  OR2_X1 U34 ( .A1(n3), .A2(A[2]), .ZN(carry[3]) );
  OR2_X1 U35 ( .A1(A[3]), .A2(carry[3]), .ZN(carry[4]) );
  OR2_X1 U36 ( .A1(A[7]), .A2(carry[7]), .ZN(carry[8]) );
  OR2_X1 U37 ( .A1(A[8]), .A2(carry[8]), .ZN(carry[9]) );
  OR2_X1 U38 ( .A1(A[9]), .A2(carry[9]), .ZN(carry[10]) );
  OR2_X1 U39 ( .A1(A[10]), .A2(carry[10]), .ZN(carry[11]) );
  OR2_X1 U40 ( .A1(A[11]), .A2(carry[11]), .ZN(carry[12]) );
  OR2_X1 U41 ( .A1(A[12]), .A2(carry[12]), .ZN(carry[13]) );
  OR2_X1 U42 ( .A1(A[13]), .A2(carry[13]), .ZN(carry[14]) );
  OR2_X1 U43 ( .A1(A[14]), .A2(carry[14]), .ZN(carry[15]) );
  OR2_X1 U44 ( .A1(A[15]), .A2(carry[15]), .ZN(carry[16]) );
  OR2_X1 U45 ( .A1(A[16]), .A2(carry[16]), .ZN(carry[17]) );
  OR2_X1 U46 ( .A1(A[22]), .A2(carry[22]), .ZN(carry[23]) );
  OR2_X1 U47 ( .A1(A[23]), .A2(carry[23]), .ZN(carry[24]) );
  OR2_X1 U48 ( .A1(A[24]), .A2(carry[24]), .ZN(carry[25]) );
  OR2_X1 U49 ( .A1(A[25]), .A2(carry[25]), .ZN(carry[26]) );
  OR2_X1 U50 ( .A1(A[26]), .A2(carry[26]), .ZN(carry[27]) );
  OR2_X1 U51 ( .A1(A[27]), .A2(carry[27]), .ZN(carry[28]) );
  OR2_X1 U52 ( .A1(A[28]), .A2(carry[28]), .ZN(carry[29]) );
  OR2_X1 U53 ( .A1(A[29]), .A2(carry[29]), .ZN(carry[30]) );
  OR2_X1 U54 ( .A1(A[4]), .A2(carry[4]), .ZN(carry[5]) );
  OR2_X1 U55 ( .A1(A[5]), .A2(carry[5]), .ZN(carry[6]) );
  OR2_X1 U56 ( .A1(A[6]), .A2(carry[6]), .ZN(carry[7]) );
  INV_X1 U57 ( .A(B[2]), .ZN(n3) );
  OR2_X1 U58 ( .A1(A[17]), .A2(carry[17]), .ZN(carry[18]) );
  OR2_X1 U59 ( .A1(A[18]), .A2(carry[18]), .ZN(carry[19]) );
  OR2_X1 U60 ( .A1(A[19]), .A2(carry[19]), .ZN(carry[20]) );
  OR2_X1 U61 ( .A1(A[20]), .A2(carry[20]), .ZN(carry[21]) );
  OR2_X1 U62 ( .A1(A[21]), .A2(carry[21]), .ZN(carry[22]) );
endmodule



    module stall_detection_unit_op_code_size6_func_size11_PC_reg_size32_reg_file_size32_DW01_sub_1 ( 
        A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   \A[0] , n1, n2, n3;
  wire   [32:0] carry;
  assign DIFF[1] = A[1];
  assign DIFF[0] = \A[0] ;
  assign \A[0]  = A[0];

  INV_X1 U1 ( .A(B[2]), .ZN(n3) );
  INV_X1 U2 ( .A(carry[30]), .ZN(n2) );
  XNOR2_X1 U3 ( .A(A[8]), .B(carry[8]), .ZN(DIFF[8]) );
  XNOR2_X1 U4 ( .A(A[9]), .B(carry[9]), .ZN(DIFF[9]) );
  XNOR2_X1 U5 ( .A(A[10]), .B(carry[10]), .ZN(DIFF[10]) );
  XNOR2_X1 U6 ( .A(A[11]), .B(carry[11]), .ZN(DIFF[11]) );
  XNOR2_X1 U7 ( .A(A[12]), .B(carry[12]), .ZN(DIFF[12]) );
  XNOR2_X1 U8 ( .A(A[13]), .B(carry[13]), .ZN(DIFF[13]) );
  XNOR2_X1 U9 ( .A(A[14]), .B(carry[14]), .ZN(DIFF[14]) );
  XNOR2_X1 U10 ( .A(A[15]), .B(carry[15]), .ZN(DIFF[15]) );
  XNOR2_X1 U11 ( .A(A[3]), .B(carry[3]), .ZN(DIFF[3]) );
  XNOR2_X1 U12 ( .A(A[4]), .B(carry[4]), .ZN(DIFF[4]) );
  XNOR2_X1 U13 ( .A(A[5]), .B(carry[5]), .ZN(DIFF[5]) );
  XNOR2_X1 U14 ( .A(A[6]), .B(carry[6]), .ZN(DIFF[6]) );
  XNOR2_X1 U15 ( .A(A[7]), .B(carry[7]), .ZN(DIFF[7]) );
  XNOR2_X1 U16 ( .A(A[16]), .B(carry[16]), .ZN(DIFF[16]) );
  XNOR2_X1 U17 ( .A(A[17]), .B(carry[17]), .ZN(DIFF[17]) );
  XNOR2_X1 U18 ( .A(A[18]), .B(carry[18]), .ZN(DIFF[18]) );
  XNOR2_X1 U19 ( .A(A[19]), .B(carry[19]), .ZN(DIFF[19]) );
  XNOR2_X1 U20 ( .A(A[20]), .B(carry[20]), .ZN(DIFF[20]) );
  XNOR2_X1 U21 ( .A(A[21]), .B(carry[21]), .ZN(DIFF[21]) );
  XNOR2_X1 U22 ( .A(A[22]), .B(carry[22]), .ZN(DIFF[22]) );
  XNOR2_X1 U23 ( .A(A[23]), .B(carry[23]), .ZN(DIFF[23]) );
  XNOR2_X1 U24 ( .A(A[24]), .B(carry[24]), .ZN(DIFF[24]) );
  XNOR2_X1 U25 ( .A(A[25]), .B(carry[25]), .ZN(DIFF[25]) );
  XNOR2_X1 U26 ( .A(A[26]), .B(carry[26]), .ZN(DIFF[26]) );
  XNOR2_X1 U27 ( .A(A[27]), .B(carry[27]), .ZN(DIFF[27]) );
  XNOR2_X1 U28 ( .A(A[28]), .B(carry[28]), .ZN(DIFF[28]) );
  XNOR2_X1 U29 ( .A(A[29]), .B(carry[29]), .ZN(DIFF[29]) );
  XNOR2_X1 U30 ( .A(A[30]), .B(carry[30]), .ZN(DIFF[30]) );
  XNOR2_X1 U31 ( .A(n3), .B(A[2]), .ZN(DIFF[2]) );
  XNOR2_X1 U32 ( .A(A[31]), .B(carry[31]), .ZN(DIFF[31]) );
  NAND2_X1 U33 ( .A1(n1), .A2(n2), .ZN(carry[31]) );
  INV_X1 U34 ( .A(A[30]), .ZN(n1) );
  OR2_X1 U35 ( .A1(n3), .A2(A[2]), .ZN(carry[3]) );
  OR2_X1 U36 ( .A1(A[3]), .A2(carry[3]), .ZN(carry[4]) );
  OR2_X1 U37 ( .A1(A[4]), .A2(carry[4]), .ZN(carry[5]) );
  OR2_X1 U38 ( .A1(A[5]), .A2(carry[5]), .ZN(carry[6]) );
  OR2_X1 U39 ( .A1(A[6]), .A2(carry[6]), .ZN(carry[7]) );
  OR2_X1 U40 ( .A1(A[7]), .A2(carry[7]), .ZN(carry[8]) );
  OR2_X1 U41 ( .A1(A[8]), .A2(carry[8]), .ZN(carry[9]) );
  OR2_X1 U42 ( .A1(A[9]), .A2(carry[9]), .ZN(carry[10]) );
  OR2_X1 U43 ( .A1(A[10]), .A2(carry[10]), .ZN(carry[11]) );
  OR2_X1 U44 ( .A1(A[11]), .A2(carry[11]), .ZN(carry[12]) );
  OR2_X1 U45 ( .A1(A[12]), .A2(carry[12]), .ZN(carry[13]) );
  OR2_X1 U46 ( .A1(A[13]), .A2(carry[13]), .ZN(carry[14]) );
  OR2_X1 U47 ( .A1(A[14]), .A2(carry[14]), .ZN(carry[15]) );
  OR2_X1 U48 ( .A1(A[15]), .A2(carry[15]), .ZN(carry[16]) );
  OR2_X1 U49 ( .A1(A[16]), .A2(carry[16]), .ZN(carry[17]) );
  OR2_X1 U50 ( .A1(A[17]), .A2(carry[17]), .ZN(carry[18]) );
  OR2_X1 U51 ( .A1(A[18]), .A2(carry[18]), .ZN(carry[19]) );
  OR2_X1 U52 ( .A1(A[19]), .A2(carry[19]), .ZN(carry[20]) );
  OR2_X1 U53 ( .A1(A[20]), .A2(carry[20]), .ZN(carry[21]) );
  OR2_X1 U54 ( .A1(A[21]), .A2(carry[21]), .ZN(carry[22]) );
  OR2_X1 U55 ( .A1(A[22]), .A2(carry[22]), .ZN(carry[23]) );
  OR2_X1 U56 ( .A1(A[23]), .A2(carry[23]), .ZN(carry[24]) );
  OR2_X1 U57 ( .A1(A[24]), .A2(carry[24]), .ZN(carry[25]) );
  OR2_X1 U58 ( .A1(A[25]), .A2(carry[25]), .ZN(carry[26]) );
  OR2_X1 U59 ( .A1(A[26]), .A2(carry[26]), .ZN(carry[27]) );
  OR2_X1 U60 ( .A1(A[27]), .A2(carry[27]), .ZN(carry[28]) );
  OR2_X1 U61 ( .A1(A[28]), .A2(carry[28]), .ZN(carry[29]) );
  OR2_X1 U62 ( .A1(A[29]), .A2(carry[29]), .ZN(carry[30]) );
endmodule



    module stall_detection_unit_op_code_size6_func_size11_PC_reg_size32_reg_file_size32_DW01_sub_2 ( 
        A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   \A[0] , n1, n2, n3;
  wire   [32:0] carry;
  assign DIFF[1] = A[1];
  assign DIFF[0] = \A[0] ;
  assign \A[0]  = A[0];

  XNOR2_X1 U1 ( .A(A[10]), .B(carry[10]), .ZN(DIFF[10]) );
  XNOR2_X1 U2 ( .A(A[11]), .B(carry[11]), .ZN(DIFF[11]) );
  XNOR2_X1 U3 ( .A(A[13]), .B(carry[13]), .ZN(DIFF[13]) );
  XNOR2_X1 U4 ( .A(A[15]), .B(carry[15]), .ZN(DIFF[15]) );
  XNOR2_X1 U5 ( .A(A[16]), .B(carry[16]), .ZN(DIFF[16]) );
  XNOR2_X1 U6 ( .A(A[17]), .B(carry[17]), .ZN(DIFF[17]) );
  XNOR2_X1 U7 ( .A(A[18]), .B(carry[18]), .ZN(DIFF[18]) );
  XNOR2_X1 U8 ( .A(A[19]), .B(carry[19]), .ZN(DIFF[19]) );
  XNOR2_X1 U9 ( .A(A[5]), .B(carry[5]), .ZN(DIFF[5]) );
  XNOR2_X1 U10 ( .A(A[8]), .B(carry[8]), .ZN(DIFF[8]) );
  XNOR2_X1 U11 ( .A(A[9]), .B(carry[9]), .ZN(DIFF[9]) );
  XNOR2_X1 U12 ( .A(A[20]), .B(carry[20]), .ZN(DIFF[20]) );
  XNOR2_X1 U13 ( .A(A[21]), .B(carry[21]), .ZN(DIFF[21]) );
  XNOR2_X1 U14 ( .A(A[22]), .B(carry[22]), .ZN(DIFF[22]) );
  XNOR2_X1 U15 ( .A(A[23]), .B(carry[23]), .ZN(DIFF[23]) );
  XNOR2_X1 U16 ( .A(A[24]), .B(carry[24]), .ZN(DIFF[24]) );
  XNOR2_X1 U17 ( .A(A[25]), .B(carry[25]), .ZN(DIFF[25]) );
  XNOR2_X1 U18 ( .A(A[26]), .B(carry[26]), .ZN(DIFF[26]) );
  XNOR2_X1 U19 ( .A(A[27]), .B(carry[27]), .ZN(DIFF[27]) );
  XNOR2_X1 U20 ( .A(A[28]), .B(carry[28]), .ZN(DIFF[28]) );
  XNOR2_X1 U21 ( .A(A[29]), .B(carry[29]), .ZN(DIFF[29]) );
  XNOR2_X1 U22 ( .A(A[30]), .B(carry[30]), .ZN(DIFF[30]) );
  XNOR2_X1 U23 ( .A(A[7]), .B(carry[7]), .ZN(DIFF[7]) );
  XNOR2_X1 U24 ( .A(n3), .B(A[2]), .ZN(DIFF[2]) );
  XNOR2_X1 U25 ( .A(A[3]), .B(carry[3]), .ZN(DIFF[3]) );
  XNOR2_X1 U26 ( .A(A[4]), .B(carry[4]), .ZN(DIFF[4]) );
  XNOR2_X1 U27 ( .A(A[12]), .B(carry[12]), .ZN(DIFF[12]) );
  XNOR2_X1 U28 ( .A(A[14]), .B(carry[14]), .ZN(DIFF[14]) );
  XNOR2_X1 U29 ( .A(A[6]), .B(carry[6]), .ZN(DIFF[6]) );
  XNOR2_X1 U30 ( .A(A[31]), .B(carry[31]), .ZN(DIFF[31]) );
  NAND2_X1 U31 ( .A1(n1), .A2(n2), .ZN(carry[31]) );
  INV_X1 U32 ( .A(A[30]), .ZN(n1) );
  INV_X1 U33 ( .A(carry[30]), .ZN(n2) );
  OR2_X1 U34 ( .A1(n3), .A2(A[2]), .ZN(carry[3]) );
  OR2_X1 U35 ( .A1(A[3]), .A2(carry[3]), .ZN(carry[4]) );
  OR2_X1 U36 ( .A1(A[4]), .A2(carry[4]), .ZN(carry[5]) );
  OR2_X1 U37 ( .A1(A[5]), .A2(carry[5]), .ZN(carry[6]) );
  OR2_X1 U38 ( .A1(A[6]), .A2(carry[6]), .ZN(carry[7]) );
  OR2_X1 U39 ( .A1(A[7]), .A2(carry[7]), .ZN(carry[8]) );
  OR2_X1 U40 ( .A1(A[8]), .A2(carry[8]), .ZN(carry[9]) );
  OR2_X1 U41 ( .A1(A[9]), .A2(carry[9]), .ZN(carry[10]) );
  OR2_X1 U42 ( .A1(A[10]), .A2(carry[10]), .ZN(carry[11]) );
  OR2_X1 U43 ( .A1(A[11]), .A2(carry[11]), .ZN(carry[12]) );
  OR2_X1 U44 ( .A1(A[12]), .A2(carry[12]), .ZN(carry[13]) );
  OR2_X1 U45 ( .A1(A[13]), .A2(carry[13]), .ZN(carry[14]) );
  OR2_X1 U46 ( .A1(A[14]), .A2(carry[14]), .ZN(carry[15]) );
  OR2_X1 U47 ( .A1(A[15]), .A2(carry[15]), .ZN(carry[16]) );
  OR2_X1 U48 ( .A1(A[16]), .A2(carry[16]), .ZN(carry[17]) );
  OR2_X1 U49 ( .A1(A[17]), .A2(carry[17]), .ZN(carry[18]) );
  OR2_X1 U50 ( .A1(A[18]), .A2(carry[18]), .ZN(carry[19]) );
  OR2_X1 U51 ( .A1(A[19]), .A2(carry[19]), .ZN(carry[20]) );
  OR2_X1 U52 ( .A1(A[20]), .A2(carry[20]), .ZN(carry[21]) );
  OR2_X1 U53 ( .A1(A[21]), .A2(carry[21]), .ZN(carry[22]) );
  OR2_X1 U54 ( .A1(A[22]), .A2(carry[22]), .ZN(carry[23]) );
  OR2_X1 U55 ( .A1(A[23]), .A2(carry[23]), .ZN(carry[24]) );
  OR2_X1 U56 ( .A1(A[24]), .A2(carry[24]), .ZN(carry[25]) );
  OR2_X1 U57 ( .A1(A[25]), .A2(carry[25]), .ZN(carry[26]) );
  OR2_X1 U58 ( .A1(A[26]), .A2(carry[26]), .ZN(carry[27]) );
  OR2_X1 U59 ( .A1(A[27]), .A2(carry[27]), .ZN(carry[28]) );
  OR2_X1 U60 ( .A1(A[28]), .A2(carry[28]), .ZN(carry[29]) );
  OR2_X1 U61 ( .A1(A[29]), .A2(carry[29]), .ZN(carry[30]) );
  INV_X1 U62 ( .A(B[2]), .ZN(n3) );
endmodule



    module stall_detection_unit_op_code_size6_func_size11_PC_reg_size32_reg_file_size32_DW01_sub_3 ( 
        A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   \A[0] , n1, n2;
  wire   [32:0] carry;
  assign DIFF[1] = A[1];
  assign DIFF[0] = \A[0] ;
  assign \A[0]  = A[0];

  XNOR2_X1 U1 ( .A(A[10]), .B(carry[10]), .ZN(DIFF[10]) );
  XNOR2_X1 U2 ( .A(A[11]), .B(carry[11]), .ZN(DIFF[11]) );
  XNOR2_X1 U3 ( .A(A[13]), .B(carry[13]), .ZN(DIFF[13]) );
  XNOR2_X1 U4 ( .A(A[15]), .B(carry[15]), .ZN(DIFF[15]) );
  XNOR2_X1 U5 ( .A(A[16]), .B(carry[16]), .ZN(DIFF[16]) );
  XNOR2_X1 U6 ( .A(A[17]), .B(carry[17]), .ZN(DIFF[17]) );
  XNOR2_X1 U7 ( .A(A[18]), .B(carry[18]), .ZN(DIFF[18]) );
  XNOR2_X1 U8 ( .A(A[19]), .B(carry[19]), .ZN(DIFF[19]) );
  XNOR2_X1 U9 ( .A(A[5]), .B(carry[5]), .ZN(DIFF[5]) );
  XNOR2_X1 U10 ( .A(A[8]), .B(carry[8]), .ZN(DIFF[8]) );
  XNOR2_X1 U11 ( .A(A[9]), .B(carry[9]), .ZN(DIFF[9]) );
  XNOR2_X1 U12 ( .A(A[20]), .B(carry[20]), .ZN(DIFF[20]) );
  XNOR2_X1 U13 ( .A(A[21]), .B(carry[21]), .ZN(DIFF[21]) );
  XNOR2_X1 U14 ( .A(A[22]), .B(carry[22]), .ZN(DIFF[22]) );
  XNOR2_X1 U15 ( .A(A[23]), .B(carry[23]), .ZN(DIFF[23]) );
  XNOR2_X1 U16 ( .A(A[24]), .B(carry[24]), .ZN(DIFF[24]) );
  XNOR2_X1 U17 ( .A(A[25]), .B(carry[25]), .ZN(DIFF[25]) );
  XNOR2_X1 U18 ( .A(A[26]), .B(carry[26]), .ZN(DIFF[26]) );
  XNOR2_X1 U19 ( .A(A[27]), .B(carry[27]), .ZN(DIFF[27]) );
  XNOR2_X1 U20 ( .A(A[28]), .B(carry[28]), .ZN(DIFF[28]) );
  XNOR2_X1 U21 ( .A(A[29]), .B(carry[29]), .ZN(DIFF[29]) );
  XNOR2_X1 U22 ( .A(A[30]), .B(carry[30]), .ZN(DIFF[30]) );
  XNOR2_X1 U23 ( .A(A[7]), .B(carry[7]), .ZN(DIFF[7]) );
  INV_X1 U24 ( .A(A[2]), .ZN(DIFF[2]) );
  XNOR2_X1 U25 ( .A(A[3]), .B(A[2]), .ZN(DIFF[3]) );
  XNOR2_X1 U26 ( .A(A[4]), .B(carry[4]), .ZN(DIFF[4]) );
  XNOR2_X1 U27 ( .A(A[12]), .B(carry[12]), .ZN(DIFF[12]) );
  XNOR2_X1 U28 ( .A(A[14]), .B(carry[14]), .ZN(DIFF[14]) );
  XNOR2_X1 U29 ( .A(A[6]), .B(carry[6]), .ZN(DIFF[6]) );
  OR2_X1 U30 ( .A1(A[3]), .A2(A[2]), .ZN(carry[4]) );
  XNOR2_X1 U31 ( .A(A[31]), .B(carry[31]), .ZN(DIFF[31]) );
  NAND2_X1 U32 ( .A1(n1), .A2(n2), .ZN(carry[31]) );
  INV_X1 U33 ( .A(A[30]), .ZN(n1) );
  INV_X1 U34 ( .A(carry[30]), .ZN(n2) );
  OR2_X1 U35 ( .A1(A[4]), .A2(carry[4]), .ZN(carry[5]) );
  OR2_X1 U36 ( .A1(A[7]), .A2(carry[7]), .ZN(carry[8]) );
  OR2_X1 U37 ( .A1(A[8]), .A2(carry[8]), .ZN(carry[9]) );
  OR2_X1 U38 ( .A1(A[9]), .A2(carry[9]), .ZN(carry[10]) );
  OR2_X1 U39 ( .A1(A[10]), .A2(carry[10]), .ZN(carry[11]) );
  OR2_X1 U40 ( .A1(A[11]), .A2(carry[11]), .ZN(carry[12]) );
  OR2_X1 U41 ( .A1(A[12]), .A2(carry[12]), .ZN(carry[13]) );
  OR2_X1 U42 ( .A1(A[13]), .A2(carry[13]), .ZN(carry[14]) );
  OR2_X1 U43 ( .A1(A[14]), .A2(carry[14]), .ZN(carry[15]) );
  OR2_X1 U44 ( .A1(A[15]), .A2(carry[15]), .ZN(carry[16]) );
  OR2_X1 U45 ( .A1(A[16]), .A2(carry[16]), .ZN(carry[17]) );
  OR2_X1 U46 ( .A1(A[23]), .A2(carry[23]), .ZN(carry[24]) );
  OR2_X1 U47 ( .A1(A[24]), .A2(carry[24]), .ZN(carry[25]) );
  OR2_X1 U48 ( .A1(A[25]), .A2(carry[25]), .ZN(carry[26]) );
  OR2_X1 U49 ( .A1(A[26]), .A2(carry[26]), .ZN(carry[27]) );
  OR2_X1 U50 ( .A1(A[27]), .A2(carry[27]), .ZN(carry[28]) );
  OR2_X1 U51 ( .A1(A[28]), .A2(carry[28]), .ZN(carry[29]) );
  OR2_X1 U52 ( .A1(A[29]), .A2(carry[29]), .ZN(carry[30]) );
  OR2_X1 U53 ( .A1(A[5]), .A2(carry[5]), .ZN(carry[6]) );
  OR2_X1 U54 ( .A1(A[6]), .A2(carry[6]), .ZN(carry[7]) );
  OR2_X1 U55 ( .A1(A[17]), .A2(carry[17]), .ZN(carry[18]) );
  OR2_X1 U56 ( .A1(A[18]), .A2(carry[18]), .ZN(carry[19]) );
  OR2_X1 U57 ( .A1(A[19]), .A2(carry[19]), .ZN(carry[20]) );
  OR2_X1 U58 ( .A1(A[20]), .A2(carry[20]), .ZN(carry[21]) );
  OR2_X1 U59 ( .A1(A[21]), .A2(carry[21]), .ZN(carry[22]) );
  OR2_X1 U60 ( .A1(A[22]), .A2(carry[22]), .ZN(carry[23]) );
endmodule



    module stall_detection_unit_op_code_size6_func_size11_PC_reg_size32_reg_file_size32 ( 
        opcode, RSA, RSB, RD, FUNC, EXE_RD, NPC_in, Ld, RD_inmul, 
        flag_structHzd, flag_ismul, opcode_out, RD_out, FUNC_out, NPC_out, 
        PC_sel );
  input [5:0] opcode;
  input [4:0] RSA;
  input [4:0] RSB;
  input [4:0] RD;
  input [10:0] FUNC;
  input [4:0] EXE_RD;
  input [31:0] NPC_in;
  input [4:0] RD_inmul;
  output [5:0] opcode_out;
  output [4:0] RD_out;
  output [10:0] FUNC_out;
  output [31:0] NPC_out;
  input Ld, flag_structHzd, flag_ismul;
  output PC_sel;
  wire   n172, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N104, N105, N106, N107, N108, N109, N110,
         N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121,
         N122, N123, N124, N125, N126, N127, N128, N129, N130, N131, N132,
         N133, N134, N135, N141, N142, N143, N144, N145, N146, N147, N148,
         N149, N150, N151, N152, N153, N154, N155, N156, N157, N158, N159,
         N160, N161, N162, N163, N164, N165, N166, N167, N168, N169, N170,
         N171, N172, N265, N266, N267, N268, N269, N270, N271, N272, N273,
         N274, N275, N276, N277, N278, N279, N280, N281, N282, N283, N284,
         N285, N286, N287, N288, N289, N290, N291, N292, N293, N294, N295,
         N296, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n29, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171;
  assign FUNC_out[10] = FUNC[10];
  assign FUNC_out[9] = FUNC[9];
  assign FUNC_out[8] = FUNC[8];
  assign FUNC_out[7] = FUNC[7];
  assign FUNC_out[6] = FUNC[6];
  assign FUNC_out[5] = FUNC[5];
  assign FUNC_out[4] = FUNC[4];
  assign FUNC_out[3] = FUNC[3];
  assign FUNC_out[2] = FUNC[2];
  assign FUNC_out[1] = FUNC[1];
  assign FUNC_out[0] = FUNC[0];

  stall_detection_unit_op_code_size6_func_size11_PC_reg_size32_reg_file_size32_DW01_sub_0 sub_100_aco ( 
        .A(NPC_in), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, flag_structHzd, 1'b0, 
        1'b0}), .CI(1'b0), .DIFF({N296, N295, N294, N293, N292, N291, N290, 
        N289, N288, N287, N286, N285, N284, N283, N282, N281, N280, N279, N278, 
        N277, N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, 
        N265}) );
  stall_detection_unit_op_code_size6_func_size11_PC_reg_size32_reg_file_size32_DW01_sub_1 sub_73_aco ( 
        .A(NPC_in), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n171, 1'b0, 1'b0}), 
        .CI(1'b0), .DIFF({N135, N134, N133, N132, N131, N130, N129, N128, N127, 
        N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, 
        N114, N113, N112, N111, N110, N109, N108, N107, N106, N105, N104}) );
  stall_detection_unit_op_code_size6_func_size11_PC_reg_size32_reg_file_size32_DW01_sub_2 sub_60_aco ( 
        .A(NPC_in), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n170, 1'b0, 1'b0}), 
        .CI(1'b0), .DIFF({N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, 
        N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, 
        N41, N40, N39, N38, N37, N36, N35, N34}) );
  stall_detection_unit_op_code_size6_func_size11_PC_reg_size32_reg_file_size32_DW01_sub_3 r107 ( 
        .A(NPC_in), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0}), 
        .CI(1'b0), .DIFF({N172, N171, N170, N169, N168, N167, N166, N165, N164, 
        N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, 
        N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141}) );
  NOR2_X2 U6 ( .A1(PC_sel), .A2(n25), .ZN(opcode_out[3]) );
  NOR2_X2 U9 ( .A1(PC_sel), .A2(n22), .ZN(opcode_out[5]) );
  BUF_X1 U10 ( .A(n172), .Z(PC_sel) );
  BUF_X1 U11 ( .A(n16), .Z(n18) );
  BUF_X1 U12 ( .A(n19), .Z(n21) );
  BUF_X1 U13 ( .A(n57), .Z(n15) );
  BUF_X1 U14 ( .A(n4), .Z(n6) );
  BUF_X1 U15 ( .A(n4), .Z(n7) );
  BUF_X1 U16 ( .A(n5), .Z(n9) );
  BUF_X1 U17 ( .A(n57), .Z(n13) );
  BUF_X1 U18 ( .A(n5), .Z(n8) );
  BUF_X1 U20 ( .A(n57), .Z(n14) );
  BUF_X1 U21 ( .A(n42), .Z(n10) );
  BUF_X1 U22 ( .A(n42), .Z(n11) );
  BUF_X1 U23 ( .A(n41), .Z(n4) );
  BUF_X1 U24 ( .A(n41), .Z(n5) );
  BUF_X1 U25 ( .A(n42), .Z(n12) );
  NOR2_X1 U26 ( .A1(n23), .A2(n9), .ZN(n172) );
  BUF_X1 U27 ( .A(n58), .Z(n16) );
  CLKBUF_X1 U28 ( .A(n16), .Z(n17) );
  BUF_X1 U29 ( .A(n59), .Z(n19) );
  CLKBUF_X1 U30 ( .A(n19), .Z(n20) );
  OAI33_X1 U31 ( .A1(n155), .A2(n156), .A3(n157), .B1(n158), .B2(n159), .B3(
        n160), .ZN(n2) );
  CLKBUF_X1 U32 ( .A(n23), .Z(n3) );
  NAND2_X1 U33 ( .A1(n3), .A2(n24), .ZN(opcode_out[4]) );
  INV_X1 U34 ( .A(opcode[4]), .ZN(n24) );
  NAND2_X1 U35 ( .A1(n3), .A2(n29), .ZN(opcode_out[2]) );
  INV_X1 U36 ( .A(opcode[2]), .ZN(n29) );
  NOR2_X1 U37 ( .A1(PC_sel), .A2(n33), .ZN(opcode_out[1]) );
  NAND2_X1 U38 ( .A1(n3), .A2(n34), .ZN(opcode_out[0]) );
  INV_X1 U39 ( .A(opcode[0]), .ZN(n34) );
  NOR2_X1 U40 ( .A1(n35), .A2(n36), .ZN(RD_out[4]) );
  INV_X1 U41 ( .A(RD[4]), .ZN(n36) );
  NOR2_X1 U42 ( .A1(n35), .A2(n37), .ZN(RD_out[3]) );
  NOR2_X1 U43 ( .A1(n35), .A2(n38), .ZN(RD_out[2]) );
  INV_X1 U44 ( .A(RD[2]), .ZN(n38) );
  NOR2_X1 U45 ( .A1(n35), .A2(n39), .ZN(RD_out[1]) );
  NOR2_X1 U46 ( .A1(n35), .A2(n40), .ZN(RD_out[0]) );
  NOR3_X1 U47 ( .A1(n6), .A2(n10), .A3(n43), .ZN(n35) );
  INV_X1 U48 ( .A(n44), .ZN(n43) );
  MUX2_X1 U49 ( .A(n45), .B(n170), .S(Ld), .Z(n44) );
  AOI222_X1 U50 ( .A1(n171), .A2(n10), .B1(n45), .B2(n46), .C1(n170), .C2(Ld), 
        .ZN(n23) );
  INV_X1 U51 ( .A(n47), .ZN(n46) );
  OR2_X1 U52 ( .A1(flag_structHzd), .A2(n48), .ZN(n45) );
  NOR2_X1 U53 ( .A1(n49), .A2(n50), .ZN(n171) );
  AND4_X1 U54 ( .A1(n51), .A2(n52), .A3(n53), .A4(n54), .ZN(n50) );
  NOR2_X1 U55 ( .A1(RSA[1]), .A2(RSA[0]), .ZN(n54) );
  INV_X1 U56 ( .A(RSA[2]), .ZN(n53) );
  INV_X1 U57 ( .A(RSA[4]), .ZN(n52) );
  NAND2_X1 U58 ( .A1(n55), .A2(n56), .ZN(NPC_out[9]) );
  AOI222_X1 U59 ( .A1(N43), .A2(n15), .B1(N150), .B2(n18), .C1(N274), .C2(n21), 
        .ZN(n56) );
  AOI22_X1 U60 ( .A1(NPC_in[9]), .A2(n6), .B1(N113), .B2(n10), .ZN(n55) );
  NAND2_X1 U61 ( .A1(n60), .A2(n61), .ZN(NPC_out[8]) );
  AOI222_X1 U62 ( .A1(N42), .A2(n15), .B1(N149), .B2(n18), .C1(N273), .C2(n21), 
        .ZN(n61) );
  AOI22_X1 U63 ( .A1(NPC_in[8]), .A2(n6), .B1(N112), .B2(n10), .ZN(n60) );
  NAND2_X1 U64 ( .A1(n62), .A2(n63), .ZN(NPC_out[7]) );
  AOI222_X1 U65 ( .A1(N41), .A2(n15), .B1(N148), .B2(n18), .C1(N272), .C2(n21), 
        .ZN(n63) );
  AOI22_X1 U66 ( .A1(NPC_in[7]), .A2(n6), .B1(N111), .B2(n10), .ZN(n62) );
  NAND2_X1 U67 ( .A1(n64), .A2(n65), .ZN(NPC_out[6]) );
  AOI222_X1 U68 ( .A1(N40), .A2(n15), .B1(N147), .B2(n18), .C1(N271), .C2(n21), 
        .ZN(n65) );
  AOI22_X1 U69 ( .A1(NPC_in[6]), .A2(n6), .B1(N110), .B2(n10), .ZN(n64) );
  NAND2_X1 U70 ( .A1(n66), .A2(n67), .ZN(NPC_out[5]) );
  AOI222_X1 U71 ( .A1(N39), .A2(n15), .B1(N146), .B2(n17), .C1(N270), .C2(n20), 
        .ZN(n67) );
  AOI22_X1 U72 ( .A1(NPC_in[5]), .A2(n6), .B1(N109), .B2(n10), .ZN(n66) );
  NAND2_X1 U73 ( .A1(n68), .A2(n69), .ZN(NPC_out[4]) );
  AOI222_X1 U74 ( .A1(N38), .A2(n15), .B1(N145), .B2(n16), .C1(N269), .C2(n19), 
        .ZN(n69) );
  AOI22_X1 U75 ( .A1(NPC_in[4]), .A2(n6), .B1(N108), .B2(n10), .ZN(n68) );
  NAND2_X1 U76 ( .A1(n70), .A2(n71), .ZN(NPC_out[3]) );
  AOI222_X1 U77 ( .A1(N37), .A2(n15), .B1(N144), .B2(n58), .C1(N268), .C2(n59), 
        .ZN(n71) );
  AOI22_X1 U78 ( .A1(NPC_in[3]), .A2(n7), .B1(N107), .B2(n11), .ZN(n70) );
  NAND2_X1 U79 ( .A1(n72), .A2(n73), .ZN(NPC_out[31]) );
  AOI222_X1 U80 ( .A1(N65), .A2(n15), .B1(N172), .B2(n18), .C1(N296), .C2(n21), 
        .ZN(n73) );
  AOI22_X1 U81 ( .A1(NPC_in[31]), .A2(n6), .B1(N135), .B2(n10), .ZN(n72) );
  NAND2_X1 U82 ( .A1(n74), .A2(n75), .ZN(NPC_out[30]) );
  AOI222_X1 U83 ( .A1(N64), .A2(n15), .B1(N171), .B2(n18), .C1(N295), .C2(n21), 
        .ZN(n75) );
  AOI22_X1 U84 ( .A1(NPC_in[30]), .A2(n6), .B1(N134), .B2(n10), .ZN(n74) );
  NAND2_X1 U85 ( .A1(n76), .A2(n77), .ZN(NPC_out[2]) );
  AOI222_X1 U86 ( .A1(N36), .A2(n15), .B1(N143), .B2(n58), .C1(N267), .C2(n59), 
        .ZN(n77) );
  AOI22_X1 U87 ( .A1(NPC_in[2]), .A2(n6), .B1(N106), .B2(n11), .ZN(n76) );
  NAND2_X1 U88 ( .A1(n78), .A2(n79), .ZN(NPC_out[29]) );
  AOI222_X1 U89 ( .A1(N63), .A2(n14), .B1(N170), .B2(n18), .C1(N294), .C2(n21), 
        .ZN(n79) );
  AOI22_X1 U90 ( .A1(NPC_in[29]), .A2(n7), .B1(N133), .B2(n11), .ZN(n78) );
  NAND2_X1 U91 ( .A1(n80), .A2(n81), .ZN(NPC_out[28]) );
  AOI222_X1 U92 ( .A1(N62), .A2(n14), .B1(N169), .B2(n18), .C1(N293), .C2(n21), 
        .ZN(n81) );
  AOI22_X1 U93 ( .A1(NPC_in[28]), .A2(n7), .B1(N132), .B2(n11), .ZN(n80) );
  NAND2_X1 U94 ( .A1(n82), .A2(n83), .ZN(NPC_out[27]) );
  AOI222_X1 U95 ( .A1(N61), .A2(n14), .B1(N168), .B2(n18), .C1(N292), .C2(n21), 
        .ZN(n83) );
  AOI22_X1 U96 ( .A1(NPC_in[27]), .A2(n7), .B1(N131), .B2(n11), .ZN(n82) );
  NAND2_X1 U97 ( .A1(n84), .A2(n85), .ZN(NPC_out[26]) );
  AOI222_X1 U98 ( .A1(N60), .A2(n14), .B1(N167), .B2(n18), .C1(N291), .C2(n21), 
        .ZN(n85) );
  AOI22_X1 U99 ( .A1(NPC_in[26]), .A2(n7), .B1(N130), .B2(n11), .ZN(n84) );
  NAND2_X1 U100 ( .A1(n86), .A2(n87), .ZN(NPC_out[25]) );
  AOI222_X1 U101 ( .A1(N59), .A2(n14), .B1(N166), .B2(n18), .C1(N290), .C2(n21), .ZN(n87) );
  AOI22_X1 U102 ( .A1(NPC_in[25]), .A2(n7), .B1(N129), .B2(n11), .ZN(n86) );
  NAND2_X1 U103 ( .A1(n88), .A2(n89), .ZN(NPC_out[24]) );
  AOI222_X1 U104 ( .A1(N58), .A2(n14), .B1(N165), .B2(n18), .C1(N289), .C2(n21), .ZN(n89) );
  AOI22_X1 U105 ( .A1(NPC_in[24]), .A2(n7), .B1(N128), .B2(n11), .ZN(n88) );
  NAND2_X1 U106 ( .A1(n90), .A2(n91), .ZN(NPC_out[23]) );
  AOI222_X1 U107 ( .A1(N57), .A2(n14), .B1(N164), .B2(n18), .C1(N288), .C2(n21), .ZN(n91) );
  AOI22_X1 U108 ( .A1(NPC_in[23]), .A2(n7), .B1(N127), .B2(n11), .ZN(n90) );
  NAND2_X1 U109 ( .A1(n92), .A2(n93), .ZN(NPC_out[22]) );
  AOI222_X1 U110 ( .A1(N56), .A2(n14), .B1(N163), .B2(n18), .C1(N287), .C2(n21), .ZN(n93) );
  AOI22_X1 U111 ( .A1(NPC_in[22]), .A2(n7), .B1(N126), .B2(n11), .ZN(n92) );
  NAND2_X1 U112 ( .A1(n94), .A2(n95), .ZN(NPC_out[21]) );
  AOI222_X1 U113 ( .A1(N55), .A2(n14), .B1(N162), .B2(n18), .C1(N286), .C2(n21), .ZN(n95) );
  AOI22_X1 U114 ( .A1(NPC_in[21]), .A2(n7), .B1(N125), .B2(n11), .ZN(n94) );
  NAND2_X1 U115 ( .A1(n96), .A2(n97), .ZN(NPC_out[20]) );
  AOI222_X1 U116 ( .A1(N54), .A2(n14), .B1(N161), .B2(n18), .C1(N285), .C2(n21), .ZN(n97) );
  AOI22_X1 U117 ( .A1(NPC_in[20]), .A2(n7), .B1(N124), .B2(n12), .ZN(n96) );
  NAND2_X1 U118 ( .A1(n98), .A2(n99), .ZN(NPC_out[1]) );
  AOI222_X1 U119 ( .A1(N35), .A2(n14), .B1(N142), .B2(n18), .C1(N266), .C2(n21), .ZN(n99) );
  AOI22_X1 U120 ( .A1(NPC_in[1]), .A2(n8), .B1(N105), .B2(n12), .ZN(n98) );
  NAND2_X1 U121 ( .A1(n100), .A2(n101), .ZN(NPC_out[19]) );
  AOI222_X1 U122 ( .A1(N53), .A2(n13), .B1(N160), .B2(n17), .C1(N284), .C2(n20), .ZN(n101) );
  AOI22_X1 U123 ( .A1(NPC_in[19]), .A2(n8), .B1(N123), .B2(n12), .ZN(n100) );
  NAND2_X1 U124 ( .A1(n102), .A2(n103), .ZN(NPC_out[18]) );
  AOI222_X1 U125 ( .A1(N52), .A2(n13), .B1(N159), .B2(n17), .C1(N283), .C2(n20), .ZN(n103) );
  AOI22_X1 U126 ( .A1(NPC_in[18]), .A2(n8), .B1(N122), .B2(n12), .ZN(n102) );
  NAND2_X1 U127 ( .A1(n104), .A2(n105), .ZN(NPC_out[17]) );
  AOI222_X1 U128 ( .A1(N51), .A2(n13), .B1(N158), .B2(n17), .C1(N282), .C2(n20), .ZN(n105) );
  AOI22_X1 U129 ( .A1(NPC_in[17]), .A2(n8), .B1(N121), .B2(n12), .ZN(n104) );
  NAND2_X1 U130 ( .A1(n106), .A2(n107), .ZN(NPC_out[16]) );
  AOI222_X1 U131 ( .A1(N50), .A2(n13), .B1(N157), .B2(n17), .C1(N281), .C2(n20), .ZN(n107) );
  AOI22_X1 U132 ( .A1(NPC_in[16]), .A2(n8), .B1(N120), .B2(n12), .ZN(n106) );
  NAND2_X1 U133 ( .A1(n108), .A2(n109), .ZN(NPC_out[15]) );
  AOI222_X1 U134 ( .A1(N49), .A2(n13), .B1(N156), .B2(n17), .C1(N280), .C2(n20), .ZN(n109) );
  AOI22_X1 U135 ( .A1(NPC_in[15]), .A2(n8), .B1(N119), .B2(n12), .ZN(n108) );
  NAND2_X1 U136 ( .A1(n110), .A2(n111), .ZN(NPC_out[14]) );
  AOI222_X1 U137 ( .A1(N48), .A2(n13), .B1(N155), .B2(n17), .C1(N279), .C2(n20), .ZN(n111) );
  AOI22_X1 U138 ( .A1(NPC_in[14]), .A2(n8), .B1(N118), .B2(n12), .ZN(n110) );
  NAND2_X1 U139 ( .A1(n112), .A2(n113), .ZN(NPC_out[13]) );
  AOI222_X1 U140 ( .A1(N47), .A2(n13), .B1(N154), .B2(n17), .C1(N278), .C2(n20), .ZN(n113) );
  AOI22_X1 U141 ( .A1(NPC_in[13]), .A2(n8), .B1(N117), .B2(n12), .ZN(n112) );
  NAND2_X1 U142 ( .A1(n114), .A2(n115), .ZN(NPC_out[12]) );
  AOI222_X1 U143 ( .A1(N46), .A2(n13), .B1(N153), .B2(n17), .C1(N277), .C2(n20), .ZN(n115) );
  AOI22_X1 U144 ( .A1(NPC_in[12]), .A2(n8), .B1(N116), .B2(n12), .ZN(n114) );
  NAND2_X1 U145 ( .A1(n116), .A2(n117), .ZN(NPC_out[11]) );
  AOI222_X1 U146 ( .A1(N45), .A2(n13), .B1(N152), .B2(n17), .C1(N276), .C2(n20), .ZN(n117) );
  AOI22_X1 U147 ( .A1(NPC_in[11]), .A2(n8), .B1(N115), .B2(n12), .ZN(n116) );
  NAND2_X1 U148 ( .A1(n118), .A2(n119), .ZN(NPC_out[10]) );
  AOI222_X1 U149 ( .A1(N44), .A2(n13), .B1(N151), .B2(n17), .C1(N275), .C2(n20), .ZN(n119) );
  AOI22_X1 U150 ( .A1(NPC_in[10]), .A2(n8), .B1(N114), .B2(n12), .ZN(n118) );
  NAND2_X1 U151 ( .A1(n120), .A2(n121), .ZN(NPC_out[0]) );
  AOI222_X1 U152 ( .A1(N34), .A2(n13), .B1(N141), .B2(n17), .C1(N265), .C2(n20), .ZN(n121) );
  NOR3_X1 U153 ( .A1(n48), .A2(n9), .A3(n47), .ZN(n59) );
  NOR3_X1 U154 ( .A1(n122), .A2(n9), .A3(n47), .ZN(n58) );
  NAND2_X1 U155 ( .A1(n123), .A2(n124), .ZN(n47) );
  INV_X1 U156 ( .A(n48), .ZN(n122) );
  NAND2_X1 U157 ( .A1(n125), .A2(n126), .ZN(n48) );
  OAI21_X1 U158 ( .B1(n170), .B2(n2), .A(flag_ismul), .ZN(n126) );
  NAND2_X1 U159 ( .A1(n49), .A2(n127), .ZN(n170) );
  NAND4_X1 U160 ( .A1(n131), .A2(n129), .A3(n130), .A4(n128), .ZN(n49) );
  NOR2_X1 U161 ( .A1(n133), .A2(n132), .ZN(n131) );
  XOR2_X1 U162 ( .A(RSA[4]), .B(EXE_RD[4]), .Z(n133) );
  XOR2_X1 U163 ( .A(RSA[2]), .B(EXE_RD[2]), .Z(n132) );
  XNOR2_X1 U164 ( .A(EXE_RD[0]), .B(RSA[0]), .ZN(n130) );
  XNOR2_X1 U165 ( .A(EXE_RD[1]), .B(RSA[1]), .ZN(n129) );
  XOR2_X1 U166 ( .A(EXE_RD[3]), .B(n51), .Z(n128) );
  NAND4_X1 U167 ( .A1(n134), .A2(n135), .A3(n136), .A4(n137), .ZN(n127) );
  NOR2_X1 U168 ( .A1(n138), .A2(n139), .ZN(n137) );
  XOR2_X1 U169 ( .A(RSB[4]), .B(EXE_RD[4]), .Z(n139) );
  XOR2_X1 U170 ( .A(RSB[3]), .B(EXE_RD[3]), .Z(n138) );
  XNOR2_X1 U171 ( .A(EXE_RD[1]), .B(RSB[1]), .ZN(n136) );
  XNOR2_X1 U172 ( .A(EXE_RD[2]), .B(RSB[2]), .ZN(n135) );
  XNOR2_X1 U173 ( .A(EXE_RD[0]), .B(RSB[0]), .ZN(n134) );
  OAI21_X1 U174 ( .B1(n2), .B2(n140), .A(n141), .ZN(n125) );
  OR4_X1 U175 ( .A1(RD_inmul[3]), .A2(RD_inmul[4]), .A3(RD_inmul[2]), .A4(n142), .ZN(n141) );
  OR2_X1 U176 ( .A1(RD_inmul[1]), .A2(RD_inmul[0]), .ZN(n142) );
  OAI33_X1 U177 ( .A1(n143), .A2(n144), .A3(n145), .B1(n146), .B2(n147), .B3(
        n148), .ZN(n140) );
  XOR2_X1 U178 ( .A(RSA[4]), .B(RD_inmul[4]), .Z(n148) );
  XOR2_X1 U179 ( .A(RSA[2]), .B(RD_inmul[2]), .Z(n147) );
  NAND3_X1 U180 ( .A1(n149), .A2(n150), .A3(n151), .ZN(n146) );
  XNOR2_X1 U181 ( .A(RSA[0]), .B(RD_inmul[0]), .ZN(n151) );
  XNOR2_X1 U182 ( .A(RSA[1]), .B(RD_inmul[1]), .ZN(n150) );
  XOR2_X1 U183 ( .A(n51), .B(RD_inmul[3]), .Z(n149) );
  INV_X1 U184 ( .A(RSA[3]), .ZN(n51) );
  XOR2_X1 U185 ( .A(RSB[4]), .B(RD_inmul[4]), .Z(n145) );
  XOR2_X1 U186 ( .A(RSB[3]), .B(RD_inmul[3]), .Z(n144) );
  NAND3_X1 U187 ( .A1(n152), .A2(n153), .A3(n154), .ZN(n143) );
  XNOR2_X1 U188 ( .A(RSB[1]), .B(RD_inmul[1]), .ZN(n154) );
  XNOR2_X1 U189 ( .A(RSB[2]), .B(RD_inmul[2]), .ZN(n153) );
  XNOR2_X1 U190 ( .A(RSB[0]), .B(RD_inmul[0]), .ZN(n152) );
  XOR2_X1 U191 ( .A(RD_inmul[4]), .B(RD[4]), .Z(n160) );
  XOR2_X1 U192 ( .A(RD_inmul[2]), .B(RD[2]), .Z(n159) );
  NAND3_X1 U193 ( .A1(n161), .A2(n162), .A3(n163), .ZN(n158) );
  XOR2_X1 U194 ( .A(n40), .B(RD_inmul[0]), .Z(n163) );
  XOR2_X1 U195 ( .A(n39), .B(RD_inmul[1]), .Z(n162) );
  XOR2_X1 U196 ( .A(n37), .B(RD_inmul[3]), .Z(n161) );
  XOR2_X1 U197 ( .A(RD[4]), .B(EXE_RD[4]), .Z(n157) );
  XOR2_X1 U198 ( .A(RD[2]), .B(EXE_RD[2]), .Z(n156) );
  NAND3_X1 U199 ( .A1(n164), .A2(n165), .A3(n166), .ZN(n155) );
  XOR2_X1 U200 ( .A(n40), .B(EXE_RD[0]), .Z(n166) );
  INV_X1 U201 ( .A(RD[0]), .ZN(n40) );
  XOR2_X1 U202 ( .A(n39), .B(EXE_RD[1]), .Z(n165) );
  INV_X1 U203 ( .A(RD[1]), .ZN(n39) );
  XOR2_X1 U204 ( .A(EXE_RD[3]), .B(n37), .Z(n164) );
  INV_X1 U205 ( .A(RD[3]), .ZN(n37) );
  NOR2_X1 U206 ( .A1(n124), .A2(n9), .ZN(n57) );
  INV_X1 U207 ( .A(Ld), .ZN(n124) );
  AOI22_X1 U208 ( .A1(NPC_in[0]), .A2(n6), .B1(N104), .B2(n10), .ZN(n120) );
  NOR2_X1 U209 ( .A1(n123), .A2(Ld), .ZN(n42) );
  NAND4_X1 U210 ( .A1(n167), .A2(n168), .A3(n25), .A4(n22), .ZN(n123) );
  INV_X1 U211 ( .A(opcode[5]), .ZN(n22) );
  INV_X1 U212 ( .A(opcode[3]), .ZN(n25) );
  NAND2_X1 U213 ( .A1(opcode[4]), .A2(n33), .ZN(n168) );
  MUX2_X1 U214 ( .A(opcode[4]), .B(n33), .S(opcode[2]), .Z(n167) );
  INV_X1 U215 ( .A(opcode[1]), .ZN(n33) );
  AND4_X1 U216 ( .A1(opcode[2]), .A2(opcode[0]), .A3(opcode[4]), .A4(n169), 
        .ZN(n41) );
  NOR3_X1 U217 ( .A1(opcode[1]), .A2(opcode[5]), .A3(opcode[3]), .ZN(n169) );
endmodule


module register_file_NBIT32_NREG32 ( RESET, ENABLE, RD1, RD2, WR, ADD_WR, 
        ADD_RD1, ADD_RD2, DATAIN, OUT1, OUT2 );
  input [4:0] ADD_WR;
  input [4:0] ADD_RD1;
  input [4:0] ADD_RD2;
  input [31:0] DATAIN;
  output [31:0] OUT1;
  output [31:0] OUT2;
  input RESET, ENABLE, RD1, RD2, WR;
  wire   \REGISTERS[0][31] , \REGISTERS[0][30] , \REGISTERS[0][29] ,
         \REGISTERS[0][28] , \REGISTERS[0][27] , \REGISTERS[0][26] ,
         \REGISTERS[0][25] , \REGISTERS[0][24] , \REGISTERS[0][23] ,
         \REGISTERS[0][22] , \REGISTERS[0][21] , \REGISTERS[0][20] ,
         \REGISTERS[0][19] , \REGISTERS[0][18] , \REGISTERS[0][17] ,
         \REGISTERS[0][16] , \REGISTERS[0][15] , \REGISTERS[0][14] ,
         \REGISTERS[0][13] , \REGISTERS[0][12] , \REGISTERS[0][11] ,
         \REGISTERS[0][10] , \REGISTERS[0][9] , \REGISTERS[0][8] ,
         \REGISTERS[0][7] , \REGISTERS[0][6] , \REGISTERS[0][5] ,
         \REGISTERS[0][4] , \REGISTERS[0][3] , \REGISTERS[0][2] ,
         \REGISTERS[0][1] , \REGISTERS[0][0] , \REGISTERS[1][31] ,
         \REGISTERS[1][30] , \REGISTERS[1][29] , \REGISTERS[1][28] ,
         \REGISTERS[1][27] , \REGISTERS[1][26] , \REGISTERS[1][25] ,
         \REGISTERS[1][24] , \REGISTERS[1][23] , \REGISTERS[1][22] ,
         \REGISTERS[1][21] , \REGISTERS[1][20] , \REGISTERS[1][19] ,
         \REGISTERS[1][18] , \REGISTERS[1][17] , \REGISTERS[1][16] ,
         \REGISTERS[1][15] , \REGISTERS[1][14] , \REGISTERS[1][13] ,
         \REGISTERS[1][12] , \REGISTERS[1][11] , \REGISTERS[1][10] ,
         \REGISTERS[1][9] , \REGISTERS[1][8] , \REGISTERS[1][7] ,
         \REGISTERS[1][6] , \REGISTERS[1][5] , \REGISTERS[1][4] ,
         \REGISTERS[1][3] , \REGISTERS[1][2] , \REGISTERS[1][1] ,
         \REGISTERS[1][0] , \REGISTERS[2][31] , \REGISTERS[2][30] ,
         \REGISTERS[2][29] , \REGISTERS[2][28] , \REGISTERS[2][27] ,
         \REGISTERS[2][26] , \REGISTERS[2][25] , \REGISTERS[2][24] ,
         \REGISTERS[2][23] , \REGISTERS[2][22] , \REGISTERS[2][21] ,
         \REGISTERS[2][20] , \REGISTERS[2][19] , \REGISTERS[2][18] ,
         \REGISTERS[2][17] , \REGISTERS[2][16] , \REGISTERS[2][15] ,
         \REGISTERS[2][14] , \REGISTERS[2][13] , \REGISTERS[2][12] ,
         \REGISTERS[2][11] , \REGISTERS[2][10] , \REGISTERS[2][9] ,
         \REGISTERS[2][8] , \REGISTERS[2][7] , \REGISTERS[2][6] ,
         \REGISTERS[2][5] , \REGISTERS[2][4] , \REGISTERS[2][3] ,
         \REGISTERS[2][2] , \REGISTERS[2][1] , \REGISTERS[2][0] ,
         \REGISTERS[3][31] , \REGISTERS[3][30] , \REGISTERS[3][29] ,
         \REGISTERS[3][28] , \REGISTERS[3][27] , \REGISTERS[3][26] ,
         \REGISTERS[3][25] , \REGISTERS[3][24] , \REGISTERS[3][23] ,
         \REGISTERS[3][22] , \REGISTERS[3][21] , \REGISTERS[3][20] ,
         \REGISTERS[3][19] , \REGISTERS[3][18] , \REGISTERS[3][17] ,
         \REGISTERS[3][16] , \REGISTERS[3][15] , \REGISTERS[3][14] ,
         \REGISTERS[3][13] , \REGISTERS[3][12] , \REGISTERS[3][11] ,
         \REGISTERS[3][10] , \REGISTERS[3][9] , \REGISTERS[3][8] ,
         \REGISTERS[3][7] , \REGISTERS[3][6] , \REGISTERS[3][5] ,
         \REGISTERS[3][4] , \REGISTERS[3][3] , \REGISTERS[3][2] ,
         \REGISTERS[3][1] , \REGISTERS[3][0] , \REGISTERS[4][31] ,
         \REGISTERS[4][30] , \REGISTERS[4][29] , \REGISTERS[4][28] ,
         \REGISTERS[4][27] , \REGISTERS[4][26] , \REGISTERS[4][25] ,
         \REGISTERS[4][24] , \REGISTERS[4][23] , \REGISTERS[4][22] ,
         \REGISTERS[4][21] , \REGISTERS[4][20] , \REGISTERS[4][19] ,
         \REGISTERS[4][18] , \REGISTERS[4][17] , \REGISTERS[4][16] ,
         \REGISTERS[4][15] , \REGISTERS[4][14] , \REGISTERS[4][13] ,
         \REGISTERS[4][12] , \REGISTERS[4][11] , \REGISTERS[4][10] ,
         \REGISTERS[4][9] , \REGISTERS[4][8] , \REGISTERS[4][7] ,
         \REGISTERS[4][6] , \REGISTERS[4][5] , \REGISTERS[4][4] ,
         \REGISTERS[4][3] , \REGISTERS[4][2] , \REGISTERS[4][1] ,
         \REGISTERS[4][0] , \REGISTERS[5][31] , \REGISTERS[5][30] ,
         \REGISTERS[5][29] , \REGISTERS[5][28] , \REGISTERS[5][27] ,
         \REGISTERS[5][26] , \REGISTERS[5][25] , \REGISTERS[5][24] ,
         \REGISTERS[5][23] , \REGISTERS[5][22] , \REGISTERS[5][21] ,
         \REGISTERS[5][20] , \REGISTERS[5][19] , \REGISTERS[5][18] ,
         \REGISTERS[5][17] , \REGISTERS[5][16] , \REGISTERS[5][15] ,
         \REGISTERS[5][14] , \REGISTERS[5][13] , \REGISTERS[5][12] ,
         \REGISTERS[5][11] , \REGISTERS[5][10] , \REGISTERS[5][9] ,
         \REGISTERS[5][8] , \REGISTERS[5][7] , \REGISTERS[5][6] ,
         \REGISTERS[5][5] , \REGISTERS[5][4] , \REGISTERS[5][3] ,
         \REGISTERS[5][2] , \REGISTERS[5][1] , \REGISTERS[5][0] ,
         \REGISTERS[6][31] , \REGISTERS[6][30] , \REGISTERS[6][29] ,
         \REGISTERS[6][28] , \REGISTERS[6][27] , \REGISTERS[6][26] ,
         \REGISTERS[6][25] , \REGISTERS[6][24] , \REGISTERS[6][23] ,
         \REGISTERS[6][22] , \REGISTERS[6][21] , \REGISTERS[6][20] ,
         \REGISTERS[6][19] , \REGISTERS[6][18] , \REGISTERS[6][17] ,
         \REGISTERS[6][16] , \REGISTERS[6][15] , \REGISTERS[6][14] ,
         \REGISTERS[6][13] , \REGISTERS[6][12] , \REGISTERS[6][11] ,
         \REGISTERS[6][10] , \REGISTERS[6][9] , \REGISTERS[6][8] ,
         \REGISTERS[6][7] , \REGISTERS[6][6] , \REGISTERS[6][5] ,
         \REGISTERS[6][4] , \REGISTERS[6][3] , \REGISTERS[6][2] ,
         \REGISTERS[6][1] , \REGISTERS[6][0] , \REGISTERS[7][31] ,
         \REGISTERS[7][30] , \REGISTERS[7][29] , \REGISTERS[7][28] ,
         \REGISTERS[7][27] , \REGISTERS[7][26] , \REGISTERS[7][25] ,
         \REGISTERS[7][24] , \REGISTERS[7][23] , \REGISTERS[7][22] ,
         \REGISTERS[7][21] , \REGISTERS[7][20] , \REGISTERS[7][19] ,
         \REGISTERS[7][18] , \REGISTERS[7][17] , \REGISTERS[7][16] ,
         \REGISTERS[7][15] , \REGISTERS[7][14] , \REGISTERS[7][13] ,
         \REGISTERS[7][12] , \REGISTERS[7][11] , \REGISTERS[7][10] ,
         \REGISTERS[7][9] , \REGISTERS[7][8] , \REGISTERS[7][7] ,
         \REGISTERS[7][6] , \REGISTERS[7][5] , \REGISTERS[7][4] ,
         \REGISTERS[7][3] , \REGISTERS[7][2] , \REGISTERS[7][1] ,
         \REGISTERS[7][0] , \REGISTERS[8][31] , \REGISTERS[8][30] ,
         \REGISTERS[8][29] , \REGISTERS[8][28] , \REGISTERS[8][27] ,
         \REGISTERS[8][26] , \REGISTERS[8][25] , \REGISTERS[8][24] ,
         \REGISTERS[8][23] , \REGISTERS[8][22] , \REGISTERS[8][21] ,
         \REGISTERS[8][20] , \REGISTERS[8][19] , \REGISTERS[8][18] ,
         \REGISTERS[8][17] , \REGISTERS[8][16] , \REGISTERS[8][15] ,
         \REGISTERS[8][14] , \REGISTERS[8][13] , \REGISTERS[8][12] ,
         \REGISTERS[8][11] , \REGISTERS[8][10] , \REGISTERS[8][9] ,
         \REGISTERS[8][8] , \REGISTERS[8][7] , \REGISTERS[8][6] ,
         \REGISTERS[8][5] , \REGISTERS[8][4] , \REGISTERS[8][3] ,
         \REGISTERS[8][2] , \REGISTERS[8][1] , \REGISTERS[8][0] ,
         \REGISTERS[9][31] , \REGISTERS[9][30] , \REGISTERS[9][29] ,
         \REGISTERS[9][28] , \REGISTERS[9][27] , \REGISTERS[9][26] ,
         \REGISTERS[9][25] , \REGISTERS[9][24] , \REGISTERS[9][23] ,
         \REGISTERS[9][22] , \REGISTERS[9][21] , \REGISTERS[9][20] ,
         \REGISTERS[9][19] , \REGISTERS[9][18] , \REGISTERS[9][17] ,
         \REGISTERS[9][16] , \REGISTERS[9][15] , \REGISTERS[9][14] ,
         \REGISTERS[9][13] , \REGISTERS[9][12] , \REGISTERS[9][11] ,
         \REGISTERS[9][10] , \REGISTERS[9][9] , \REGISTERS[9][8] ,
         \REGISTERS[9][7] , \REGISTERS[9][6] , \REGISTERS[9][5] ,
         \REGISTERS[9][4] , \REGISTERS[9][3] , \REGISTERS[9][2] ,
         \REGISTERS[9][1] , \REGISTERS[9][0] , \REGISTERS[10][31] ,
         \REGISTERS[10][30] , \REGISTERS[10][29] , \REGISTERS[10][28] ,
         \REGISTERS[10][27] , \REGISTERS[10][26] , \REGISTERS[10][25] ,
         \REGISTERS[10][24] , \REGISTERS[10][23] , \REGISTERS[10][22] ,
         \REGISTERS[10][21] , \REGISTERS[10][20] , \REGISTERS[10][19] ,
         \REGISTERS[10][18] , \REGISTERS[10][17] , \REGISTERS[10][16] ,
         \REGISTERS[10][15] , \REGISTERS[10][14] , \REGISTERS[10][13] ,
         \REGISTERS[10][12] , \REGISTERS[10][11] , \REGISTERS[10][10] ,
         \REGISTERS[10][9] , \REGISTERS[10][8] , \REGISTERS[10][7] ,
         \REGISTERS[10][6] , \REGISTERS[10][5] , \REGISTERS[10][4] ,
         \REGISTERS[10][3] , \REGISTERS[10][2] , \REGISTERS[10][1] ,
         \REGISTERS[10][0] , \REGISTERS[11][31] , \REGISTERS[11][30] ,
         \REGISTERS[11][29] , \REGISTERS[11][28] , \REGISTERS[11][27] ,
         \REGISTERS[11][26] , \REGISTERS[11][25] , \REGISTERS[11][24] ,
         \REGISTERS[11][23] , \REGISTERS[11][22] , \REGISTERS[11][21] ,
         \REGISTERS[11][20] , \REGISTERS[11][19] , \REGISTERS[11][18] ,
         \REGISTERS[11][17] , \REGISTERS[11][16] , \REGISTERS[11][15] ,
         \REGISTERS[11][14] , \REGISTERS[11][13] , \REGISTERS[11][12] ,
         \REGISTERS[11][11] , \REGISTERS[11][10] , \REGISTERS[11][9] ,
         \REGISTERS[11][8] , \REGISTERS[11][7] , \REGISTERS[11][6] ,
         \REGISTERS[11][5] , \REGISTERS[11][4] , \REGISTERS[11][3] ,
         \REGISTERS[11][2] , \REGISTERS[11][1] , \REGISTERS[11][0] ,
         \REGISTERS[12][31] , \REGISTERS[12][30] , \REGISTERS[12][29] ,
         \REGISTERS[12][28] , \REGISTERS[12][27] , \REGISTERS[12][26] ,
         \REGISTERS[12][25] , \REGISTERS[12][24] , \REGISTERS[12][23] ,
         \REGISTERS[12][22] , \REGISTERS[12][21] , \REGISTERS[12][20] ,
         \REGISTERS[12][19] , \REGISTERS[12][18] , \REGISTERS[12][17] ,
         \REGISTERS[12][16] , \REGISTERS[12][15] , \REGISTERS[12][14] ,
         \REGISTERS[12][13] , \REGISTERS[12][12] , \REGISTERS[12][11] ,
         \REGISTERS[12][10] , \REGISTERS[12][9] , \REGISTERS[12][8] ,
         \REGISTERS[12][7] , \REGISTERS[12][6] , \REGISTERS[12][5] ,
         \REGISTERS[12][4] , \REGISTERS[12][3] , \REGISTERS[12][2] ,
         \REGISTERS[12][1] , \REGISTERS[12][0] , \REGISTERS[13][31] ,
         \REGISTERS[13][30] , \REGISTERS[13][29] , \REGISTERS[13][28] ,
         \REGISTERS[13][27] , \REGISTERS[13][26] , \REGISTERS[13][25] ,
         \REGISTERS[13][24] , \REGISTERS[13][23] , \REGISTERS[13][22] ,
         \REGISTERS[13][21] , \REGISTERS[13][20] , \REGISTERS[13][19] ,
         \REGISTERS[13][18] , \REGISTERS[13][17] , \REGISTERS[13][16] ,
         \REGISTERS[13][15] , \REGISTERS[13][14] , \REGISTERS[13][13] ,
         \REGISTERS[13][12] , \REGISTERS[13][11] , \REGISTERS[13][10] ,
         \REGISTERS[13][9] , \REGISTERS[13][8] , \REGISTERS[13][7] ,
         \REGISTERS[13][6] , \REGISTERS[13][5] , \REGISTERS[13][4] ,
         \REGISTERS[13][3] , \REGISTERS[13][2] , \REGISTERS[13][1] ,
         \REGISTERS[13][0] , \REGISTERS[14][31] , \REGISTERS[14][30] ,
         \REGISTERS[14][29] , \REGISTERS[14][28] , \REGISTERS[14][27] ,
         \REGISTERS[14][26] , \REGISTERS[14][25] , \REGISTERS[14][24] ,
         \REGISTERS[14][23] , \REGISTERS[14][22] , \REGISTERS[14][21] ,
         \REGISTERS[14][20] , \REGISTERS[14][19] , \REGISTERS[14][18] ,
         \REGISTERS[14][17] , \REGISTERS[14][16] , \REGISTERS[14][15] ,
         \REGISTERS[14][14] , \REGISTERS[14][13] , \REGISTERS[14][12] ,
         \REGISTERS[14][11] , \REGISTERS[14][10] , \REGISTERS[14][9] ,
         \REGISTERS[14][8] , \REGISTERS[14][7] , \REGISTERS[14][6] ,
         \REGISTERS[14][5] , \REGISTERS[14][4] , \REGISTERS[14][3] ,
         \REGISTERS[14][2] , \REGISTERS[14][1] , \REGISTERS[14][0] ,
         \REGISTERS[15][31] , \REGISTERS[15][30] , \REGISTERS[15][29] ,
         \REGISTERS[15][28] , \REGISTERS[15][27] , \REGISTERS[15][26] ,
         \REGISTERS[15][25] , \REGISTERS[15][24] , \REGISTERS[15][23] ,
         \REGISTERS[15][22] , \REGISTERS[15][21] , \REGISTERS[15][20] ,
         \REGISTERS[15][19] , \REGISTERS[15][18] , \REGISTERS[15][17] ,
         \REGISTERS[15][16] , \REGISTERS[15][15] , \REGISTERS[15][14] ,
         \REGISTERS[15][13] , \REGISTERS[15][12] , \REGISTERS[15][11] ,
         \REGISTERS[15][10] , \REGISTERS[15][9] , \REGISTERS[15][8] ,
         \REGISTERS[15][7] , \REGISTERS[15][6] , \REGISTERS[15][5] ,
         \REGISTERS[15][4] , \REGISTERS[15][3] , \REGISTERS[15][2] ,
         \REGISTERS[15][1] , \REGISTERS[15][0] , \REGISTERS[16][31] ,
         \REGISTERS[16][30] , \REGISTERS[16][29] , \REGISTERS[16][28] ,
         \REGISTERS[16][27] , \REGISTERS[16][26] , \REGISTERS[16][25] ,
         \REGISTERS[16][24] , \REGISTERS[16][23] , \REGISTERS[16][22] ,
         \REGISTERS[16][21] , \REGISTERS[16][20] , \REGISTERS[16][19] ,
         \REGISTERS[16][18] , \REGISTERS[16][17] , \REGISTERS[16][16] ,
         \REGISTERS[16][15] , \REGISTERS[16][14] , \REGISTERS[16][13] ,
         \REGISTERS[16][12] , \REGISTERS[16][11] , \REGISTERS[16][10] ,
         \REGISTERS[16][9] , \REGISTERS[16][8] , \REGISTERS[16][7] ,
         \REGISTERS[16][6] , \REGISTERS[16][5] , \REGISTERS[16][4] ,
         \REGISTERS[16][3] , \REGISTERS[16][2] , \REGISTERS[16][1] ,
         \REGISTERS[16][0] , \REGISTERS[17][31] , \REGISTERS[17][30] ,
         \REGISTERS[17][29] , \REGISTERS[17][28] , \REGISTERS[17][27] ,
         \REGISTERS[17][26] , \REGISTERS[17][25] , \REGISTERS[17][24] ,
         \REGISTERS[17][23] , \REGISTERS[17][22] , \REGISTERS[17][21] ,
         \REGISTERS[17][20] , \REGISTERS[17][19] , \REGISTERS[17][18] ,
         \REGISTERS[17][17] , \REGISTERS[17][16] , \REGISTERS[17][15] ,
         \REGISTERS[17][14] , \REGISTERS[17][13] , \REGISTERS[17][12] ,
         \REGISTERS[17][11] , \REGISTERS[17][10] , \REGISTERS[17][9] ,
         \REGISTERS[17][8] , \REGISTERS[17][7] , \REGISTERS[17][6] ,
         \REGISTERS[17][5] , \REGISTERS[17][4] , \REGISTERS[17][3] ,
         \REGISTERS[17][2] , \REGISTERS[17][1] , \REGISTERS[17][0] ,
         \REGISTERS[18][31] , \REGISTERS[18][30] , \REGISTERS[18][29] ,
         \REGISTERS[18][28] , \REGISTERS[18][27] , \REGISTERS[18][26] ,
         \REGISTERS[18][25] , \REGISTERS[18][24] , \REGISTERS[18][23] ,
         \REGISTERS[18][22] , \REGISTERS[18][21] , \REGISTERS[18][20] ,
         \REGISTERS[18][19] , \REGISTERS[18][18] , \REGISTERS[18][17] ,
         \REGISTERS[18][16] , \REGISTERS[18][15] , \REGISTERS[18][14] ,
         \REGISTERS[18][13] , \REGISTERS[18][12] , \REGISTERS[18][11] ,
         \REGISTERS[18][10] , \REGISTERS[18][9] , \REGISTERS[18][8] ,
         \REGISTERS[18][7] , \REGISTERS[18][6] , \REGISTERS[18][5] ,
         \REGISTERS[18][4] , \REGISTERS[18][3] , \REGISTERS[18][2] ,
         \REGISTERS[18][1] , \REGISTERS[18][0] , \REGISTERS[19][31] ,
         \REGISTERS[19][30] , \REGISTERS[19][29] , \REGISTERS[19][28] ,
         \REGISTERS[19][27] , \REGISTERS[19][26] , \REGISTERS[19][25] ,
         \REGISTERS[19][24] , \REGISTERS[19][23] , \REGISTERS[19][22] ,
         \REGISTERS[19][21] , \REGISTERS[19][20] , \REGISTERS[19][19] ,
         \REGISTERS[19][18] , \REGISTERS[19][17] , \REGISTERS[19][16] ,
         \REGISTERS[19][15] , \REGISTERS[19][14] , \REGISTERS[19][13] ,
         \REGISTERS[19][12] , \REGISTERS[19][11] , \REGISTERS[19][10] ,
         \REGISTERS[19][9] , \REGISTERS[19][8] , \REGISTERS[19][7] ,
         \REGISTERS[19][6] , \REGISTERS[19][5] , \REGISTERS[19][4] ,
         \REGISTERS[19][3] , \REGISTERS[19][2] , \REGISTERS[19][1] ,
         \REGISTERS[19][0] , \REGISTERS[20][31] , \REGISTERS[20][30] ,
         \REGISTERS[20][29] , \REGISTERS[20][28] , \REGISTERS[20][27] ,
         \REGISTERS[20][26] , \REGISTERS[20][25] , \REGISTERS[20][24] ,
         \REGISTERS[20][23] , \REGISTERS[20][22] , \REGISTERS[20][21] ,
         \REGISTERS[20][20] , \REGISTERS[20][19] , \REGISTERS[20][18] ,
         \REGISTERS[20][17] , \REGISTERS[20][16] , \REGISTERS[20][15] ,
         \REGISTERS[20][14] , \REGISTERS[20][13] , \REGISTERS[20][12] ,
         \REGISTERS[20][11] , \REGISTERS[20][10] , \REGISTERS[20][9] ,
         \REGISTERS[20][8] , \REGISTERS[20][7] , \REGISTERS[20][6] ,
         \REGISTERS[20][5] , \REGISTERS[20][4] , \REGISTERS[20][3] ,
         \REGISTERS[20][2] , \REGISTERS[20][1] , \REGISTERS[20][0] ,
         \REGISTERS[21][31] , \REGISTERS[21][30] , \REGISTERS[21][29] ,
         \REGISTERS[21][28] , \REGISTERS[21][27] , \REGISTERS[21][26] ,
         \REGISTERS[21][25] , \REGISTERS[21][24] , \REGISTERS[21][23] ,
         \REGISTERS[21][22] , \REGISTERS[21][21] , \REGISTERS[21][20] ,
         \REGISTERS[21][19] , \REGISTERS[21][18] , \REGISTERS[21][17] ,
         \REGISTERS[21][16] , \REGISTERS[21][15] , \REGISTERS[21][14] ,
         \REGISTERS[21][13] , \REGISTERS[21][12] , \REGISTERS[21][11] ,
         \REGISTERS[21][10] , \REGISTERS[21][9] , \REGISTERS[21][8] ,
         \REGISTERS[21][7] , \REGISTERS[21][6] , \REGISTERS[21][5] ,
         \REGISTERS[21][4] , \REGISTERS[21][3] , \REGISTERS[21][2] ,
         \REGISTERS[21][1] , \REGISTERS[21][0] , \REGISTERS[22][31] ,
         \REGISTERS[22][30] , \REGISTERS[22][29] , \REGISTERS[22][28] ,
         \REGISTERS[22][27] , \REGISTERS[22][26] , \REGISTERS[22][25] ,
         \REGISTERS[22][24] , \REGISTERS[22][23] , \REGISTERS[22][22] ,
         \REGISTERS[22][21] , \REGISTERS[22][20] , \REGISTERS[22][19] ,
         \REGISTERS[22][18] , \REGISTERS[22][17] , \REGISTERS[22][16] ,
         \REGISTERS[22][15] , \REGISTERS[22][14] , \REGISTERS[22][13] ,
         \REGISTERS[22][12] , \REGISTERS[22][11] , \REGISTERS[22][10] ,
         \REGISTERS[22][9] , \REGISTERS[22][8] , \REGISTERS[22][7] ,
         \REGISTERS[22][6] , \REGISTERS[22][5] , \REGISTERS[22][4] ,
         \REGISTERS[22][3] , \REGISTERS[22][2] , \REGISTERS[22][1] ,
         \REGISTERS[22][0] , \REGISTERS[23][31] , \REGISTERS[23][30] ,
         \REGISTERS[23][29] , \REGISTERS[23][28] , \REGISTERS[23][27] ,
         \REGISTERS[23][26] , \REGISTERS[23][25] , \REGISTERS[23][24] ,
         \REGISTERS[23][23] , \REGISTERS[23][22] , \REGISTERS[23][21] ,
         \REGISTERS[23][20] , \REGISTERS[23][19] , \REGISTERS[23][18] ,
         \REGISTERS[23][17] , \REGISTERS[23][16] , \REGISTERS[23][15] ,
         \REGISTERS[23][14] , \REGISTERS[23][13] , \REGISTERS[23][12] ,
         \REGISTERS[23][11] , \REGISTERS[23][10] , \REGISTERS[23][9] ,
         \REGISTERS[23][8] , \REGISTERS[23][7] , \REGISTERS[23][6] ,
         \REGISTERS[23][5] , \REGISTERS[23][4] , \REGISTERS[23][3] ,
         \REGISTERS[23][2] , \REGISTERS[23][1] , \REGISTERS[23][0] ,
         \REGISTERS[24][31] , \REGISTERS[24][30] , \REGISTERS[24][29] ,
         \REGISTERS[24][28] , \REGISTERS[24][27] , \REGISTERS[24][26] ,
         \REGISTERS[24][25] , \REGISTERS[24][24] , \REGISTERS[24][23] ,
         \REGISTERS[24][22] , \REGISTERS[24][21] , \REGISTERS[24][20] ,
         \REGISTERS[24][19] , \REGISTERS[24][18] , \REGISTERS[24][17] ,
         \REGISTERS[24][16] , \REGISTERS[24][15] , \REGISTERS[24][14] ,
         \REGISTERS[24][13] , \REGISTERS[24][12] , \REGISTERS[24][11] ,
         \REGISTERS[24][10] , \REGISTERS[24][9] , \REGISTERS[24][8] ,
         \REGISTERS[24][7] , \REGISTERS[24][6] , \REGISTERS[24][5] ,
         \REGISTERS[24][4] , \REGISTERS[24][3] , \REGISTERS[24][2] ,
         \REGISTERS[24][1] , \REGISTERS[24][0] , \REGISTERS[25][31] ,
         \REGISTERS[25][30] , \REGISTERS[25][29] , \REGISTERS[25][28] ,
         \REGISTERS[25][27] , \REGISTERS[25][26] , \REGISTERS[25][25] ,
         \REGISTERS[25][24] , \REGISTERS[25][23] , \REGISTERS[25][22] ,
         \REGISTERS[25][21] , \REGISTERS[25][20] , \REGISTERS[25][19] ,
         \REGISTERS[25][18] , \REGISTERS[25][17] , \REGISTERS[25][16] ,
         \REGISTERS[25][15] , \REGISTERS[25][14] , \REGISTERS[25][13] ,
         \REGISTERS[25][12] , \REGISTERS[25][11] , \REGISTERS[25][10] ,
         \REGISTERS[25][9] , \REGISTERS[25][8] , \REGISTERS[25][7] ,
         \REGISTERS[25][6] , \REGISTERS[25][5] , \REGISTERS[25][4] ,
         \REGISTERS[25][3] , \REGISTERS[25][2] , \REGISTERS[25][1] ,
         \REGISTERS[25][0] , \REGISTERS[26][31] , \REGISTERS[26][30] ,
         \REGISTERS[26][29] , \REGISTERS[26][28] , \REGISTERS[26][27] ,
         \REGISTERS[26][26] , \REGISTERS[26][25] , \REGISTERS[26][24] ,
         \REGISTERS[26][23] , \REGISTERS[26][22] , \REGISTERS[26][21] ,
         \REGISTERS[26][20] , \REGISTERS[26][19] , \REGISTERS[26][18] ,
         \REGISTERS[26][17] , \REGISTERS[26][16] , \REGISTERS[26][15] ,
         \REGISTERS[26][14] , \REGISTERS[26][13] , \REGISTERS[26][12] ,
         \REGISTERS[26][11] , \REGISTERS[26][10] , \REGISTERS[26][9] ,
         \REGISTERS[26][8] , \REGISTERS[26][7] , \REGISTERS[26][6] ,
         \REGISTERS[26][5] , \REGISTERS[26][4] , \REGISTERS[26][3] ,
         \REGISTERS[26][2] , \REGISTERS[26][1] , \REGISTERS[26][0] ,
         \REGISTERS[27][31] , \REGISTERS[27][30] , \REGISTERS[27][29] ,
         \REGISTERS[27][28] , \REGISTERS[27][27] , \REGISTERS[27][26] ,
         \REGISTERS[27][25] , \REGISTERS[27][24] , \REGISTERS[27][23] ,
         \REGISTERS[27][22] , \REGISTERS[27][21] , \REGISTERS[27][20] ,
         \REGISTERS[27][19] , \REGISTERS[27][18] , \REGISTERS[27][17] ,
         \REGISTERS[27][16] , \REGISTERS[27][15] , \REGISTERS[27][14] ,
         \REGISTERS[27][13] , \REGISTERS[27][12] , \REGISTERS[27][11] ,
         \REGISTERS[27][10] , \REGISTERS[27][9] , \REGISTERS[27][8] ,
         \REGISTERS[27][7] , \REGISTERS[27][6] , \REGISTERS[27][5] ,
         \REGISTERS[27][4] , \REGISTERS[27][3] , \REGISTERS[27][2] ,
         \REGISTERS[27][1] , \REGISTERS[27][0] , \REGISTERS[28][31] ,
         \REGISTERS[28][30] , \REGISTERS[28][29] , \REGISTERS[28][28] ,
         \REGISTERS[28][27] , \REGISTERS[28][26] , \REGISTERS[28][25] ,
         \REGISTERS[28][24] , \REGISTERS[28][23] , \REGISTERS[28][22] ,
         \REGISTERS[28][21] , \REGISTERS[28][20] , \REGISTERS[28][19] ,
         \REGISTERS[28][18] , \REGISTERS[28][17] , \REGISTERS[28][16] ,
         \REGISTERS[28][15] , \REGISTERS[28][14] , \REGISTERS[28][13] ,
         \REGISTERS[28][12] , \REGISTERS[28][11] , \REGISTERS[28][10] ,
         \REGISTERS[28][9] , \REGISTERS[28][8] , \REGISTERS[28][7] ,
         \REGISTERS[28][6] , \REGISTERS[28][5] , \REGISTERS[28][4] ,
         \REGISTERS[28][3] , \REGISTERS[28][2] , \REGISTERS[28][1] ,
         \REGISTERS[28][0] , \REGISTERS[29][31] , \REGISTERS[29][30] ,
         \REGISTERS[29][29] , \REGISTERS[29][28] , \REGISTERS[29][27] ,
         \REGISTERS[29][26] , \REGISTERS[29][25] , \REGISTERS[29][24] ,
         \REGISTERS[29][23] , \REGISTERS[29][22] , \REGISTERS[29][21] ,
         \REGISTERS[29][20] , \REGISTERS[29][19] , \REGISTERS[29][18] ,
         \REGISTERS[29][17] , \REGISTERS[29][16] , \REGISTERS[29][15] ,
         \REGISTERS[29][14] , \REGISTERS[29][13] , \REGISTERS[29][12] ,
         \REGISTERS[29][11] , \REGISTERS[29][10] , \REGISTERS[29][9] ,
         \REGISTERS[29][8] , \REGISTERS[29][7] , \REGISTERS[29][6] ,
         \REGISTERS[29][5] , \REGISTERS[29][4] , \REGISTERS[29][3] ,
         \REGISTERS[29][2] , \REGISTERS[29][1] , \REGISTERS[29][0] ,
         \REGISTERS[30][31] , \REGISTERS[30][30] , \REGISTERS[30][29] ,
         \REGISTERS[30][28] , \REGISTERS[30][27] , \REGISTERS[30][26] ,
         \REGISTERS[30][25] , \REGISTERS[30][24] , \REGISTERS[30][23] ,
         \REGISTERS[30][22] , \REGISTERS[30][21] , \REGISTERS[30][20] ,
         \REGISTERS[30][19] , \REGISTERS[30][18] , \REGISTERS[30][17] ,
         \REGISTERS[30][16] , \REGISTERS[30][15] , \REGISTERS[30][14] ,
         \REGISTERS[30][13] , \REGISTERS[30][12] , \REGISTERS[30][11] ,
         \REGISTERS[30][10] , \REGISTERS[30][9] , \REGISTERS[30][8] ,
         \REGISTERS[30][7] , \REGISTERS[30][6] , \REGISTERS[30][5] ,
         \REGISTERS[30][4] , \REGISTERS[30][3] , \REGISTERS[30][2] ,
         \REGISTERS[30][1] , \REGISTERS[30][0] , \REGISTERS[31][31] ,
         \REGISTERS[31][30] , \REGISTERS[31][29] , \REGISTERS[31][28] ,
         \REGISTERS[31][27] , \REGISTERS[31][26] , \REGISTERS[31][25] ,
         \REGISTERS[31][24] , \REGISTERS[31][23] , \REGISTERS[31][22] ,
         \REGISTERS[31][21] , \REGISTERS[31][20] , \REGISTERS[31][19] ,
         \REGISTERS[31][18] , \REGISTERS[31][17] , \REGISTERS[31][16] ,
         \REGISTERS[31][15] , \REGISTERS[31][14] , \REGISTERS[31][13] ,
         \REGISTERS[31][12] , \REGISTERS[31][11] , \REGISTERS[31][10] ,
         \REGISTERS[31][9] , \REGISTERS[31][8] , \REGISTERS[31][7] ,
         \REGISTERS[31][6] , \REGISTERS[31][5] , \REGISTERS[31][4] ,
         \REGISTERS[31][3] , \REGISTERS[31][2] , \REGISTERS[31][1] ,
         \REGISTERS[31][0] , N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352,
         N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363,
         N364, N365, N366, N367, N368, N369, N370, N371, N372, N373, N374,
         N375, N376, N377, N378, N379, N380, N381, N382, N383, N384, N385,
         N386, N387, N388, N389, N390, N391, N392, N393, N394, N395, N396,
         N397, N398, N399, N400, N401, N402, N403, N404, N405, N406, N407,
         N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, N418,
         N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429,
         N430, N431, N432, N433, N434, N435, N436, N437, N438, N439, N440,
         N441, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
         n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
         n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
         n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
         n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
         n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
         n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
         n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
         n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
         n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
         n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
         n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
         n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
         n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
         n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
         n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
         n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
         n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
         n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
         n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
         n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
         n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
         n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
         n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
         n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
         n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
         n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
         n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
         n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
         n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
         n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
         n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
         n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
         n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
         n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
         n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
         n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
         n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
         n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
         n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718,
         n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
         n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
         n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748,
         n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758,
         n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768,
         n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
         n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788,
         n1789, n1790, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n1791,
         n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801,
         n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811,
         n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821,
         n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831,
         n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841,
         n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851,
         n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861,
         n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
         n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881,
         n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
         n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901,
         n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911,
         n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921,
         n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931,
         n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941,
         n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951,
         n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961,
         n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971,
         n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981,
         n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991,
         n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001,
         n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011,
         n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021,
         n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031,
         n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041,
         n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
         n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061,
         n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071,
         n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081,
         n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091,
         n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101,
         n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
         n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
         n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
         n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
         n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
         n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
         n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
         n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
         n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191,
         n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
         n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
         n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
         n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
         n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
         n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
         n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
         n2262, n2263;

  DLH_X1 \REGISTERS_reg[0][31]  ( .G(n204), .D(n328), .Q(\REGISTERS[0][31] )
         );
  DLH_X1 \REGISTERS_reg[0][30]  ( .G(n204), .D(n332), .Q(\REGISTERS[0][30] )
         );
  DLH_X1 \REGISTERS_reg[0][29]  ( .G(n204), .D(n336), .Q(\REGISTERS[0][29] )
         );
  DLH_X1 \REGISTERS_reg[0][28]  ( .G(n204), .D(n340), .Q(\REGISTERS[0][28] )
         );
  DLH_X1 \REGISTERS_reg[0][27]  ( .G(n204), .D(n344), .Q(\REGISTERS[0][27] )
         );
  DLH_X1 \REGISTERS_reg[0][26]  ( .G(n204), .D(n348), .Q(\REGISTERS[0][26] )
         );
  DLH_X1 \REGISTERS_reg[0][25]  ( .G(n204), .D(n352), .Q(\REGISTERS[0][25] )
         );
  DLH_X1 \REGISTERS_reg[0][24]  ( .G(n204), .D(n356), .Q(\REGISTERS[0][24] )
         );
  DLH_X1 \REGISTERS_reg[0][23]  ( .G(n204), .D(n360), .Q(\REGISTERS[0][23] )
         );
  DLH_X1 \REGISTERS_reg[0][22]  ( .G(n204), .D(n364), .Q(\REGISTERS[0][22] )
         );
  DLH_X1 \REGISTERS_reg[0][21]  ( .G(n205), .D(n368), .Q(\REGISTERS[0][21] )
         );
  DLH_X1 \REGISTERS_reg[0][20]  ( .G(n205), .D(n372), .Q(\REGISTERS[0][20] )
         );
  DLH_X1 \REGISTERS_reg[0][19]  ( .G(n205), .D(n376), .Q(\REGISTERS[0][19] )
         );
  DLH_X1 \REGISTERS_reg[0][18]  ( .G(n205), .D(n380), .Q(\REGISTERS[0][18] )
         );
  DLH_X1 \REGISTERS_reg[0][17]  ( .G(n205), .D(n384), .Q(\REGISTERS[0][17] )
         );
  DLH_X1 \REGISTERS_reg[0][16]  ( .G(n205), .D(n388), .Q(\REGISTERS[0][16] )
         );
  DLH_X1 \REGISTERS_reg[0][15]  ( .G(n205), .D(n392), .Q(\REGISTERS[0][15] )
         );
  DLH_X1 \REGISTERS_reg[0][14]  ( .G(n205), .D(n396), .Q(\REGISTERS[0][14] )
         );
  DLH_X1 \REGISTERS_reg[0][13]  ( .G(n205), .D(n400), .Q(\REGISTERS[0][13] )
         );
  DLH_X1 \REGISTERS_reg[0][12]  ( .G(n205), .D(n404), .Q(\REGISTERS[0][12] )
         );
  DLH_X1 \REGISTERS_reg[0][11]  ( .G(n206), .D(n408), .Q(\REGISTERS[0][11] )
         );
  DLH_X1 \REGISTERS_reg[0][10]  ( .G(n206), .D(n412), .Q(\REGISTERS[0][10] )
         );
  DLH_X1 \REGISTERS_reg[0][9]  ( .G(n206), .D(n416), .Q(\REGISTERS[0][9] ) );
  DLH_X1 \REGISTERS_reg[0][8]  ( .G(n206), .D(n420), .Q(\REGISTERS[0][8] ) );
  DLH_X1 \REGISTERS_reg[0][7]  ( .G(n206), .D(n424), .Q(\REGISTERS[0][7] ) );
  DLH_X1 \REGISTERS_reg[0][6]  ( .G(n206), .D(n428), .Q(\REGISTERS[0][6] ) );
  DLH_X1 \REGISTERS_reg[0][5]  ( .G(n206), .D(n432), .Q(\REGISTERS[0][5] ) );
  DLH_X1 \REGISTERS_reg[0][4]  ( .G(n206), .D(n436), .Q(\REGISTERS[0][4] ) );
  DLH_X1 \REGISTERS_reg[0][3]  ( .G(n206), .D(n440), .Q(\REGISTERS[0][3] ) );
  DLH_X1 \REGISTERS_reg[0][2]  ( .G(n206), .D(n444), .Q(\REGISTERS[0][2] ) );
  DLH_X1 \REGISTERS_reg[0][1]  ( .G(n207), .D(n448), .Q(\REGISTERS[0][1] ) );
  DLH_X1 \REGISTERS_reg[0][0]  ( .G(n207), .D(n452), .Q(\REGISTERS[0][0] ) );
  DLH_X1 \REGISTERS_reg[1][31]  ( .G(n211), .D(n328), .Q(\REGISTERS[1][31] )
         );
  DLH_X1 \REGISTERS_reg[1][30]  ( .G(n211), .D(n332), .Q(\REGISTERS[1][30] )
         );
  DLH_X1 \REGISTERS_reg[1][29]  ( .G(n210), .D(n336), .Q(\REGISTERS[1][29] )
         );
  DLH_X1 \REGISTERS_reg[1][28]  ( .G(n210), .D(n340), .Q(\REGISTERS[1][28] )
         );
  DLH_X1 \REGISTERS_reg[1][27]  ( .G(n210), .D(n344), .Q(\REGISTERS[1][27] )
         );
  DLH_X1 \REGISTERS_reg[1][26]  ( .G(n210), .D(n348), .Q(\REGISTERS[1][26] )
         );
  DLH_X1 \REGISTERS_reg[1][25]  ( .G(n210), .D(n352), .Q(\REGISTERS[1][25] )
         );
  DLH_X1 \REGISTERS_reg[1][24]  ( .G(n210), .D(n356), .Q(\REGISTERS[1][24] )
         );
  DLH_X1 \REGISTERS_reg[1][23]  ( .G(n210), .D(n360), .Q(\REGISTERS[1][23] )
         );
  DLH_X1 \REGISTERS_reg[1][22]  ( .G(n210), .D(n364), .Q(\REGISTERS[1][22] )
         );
  DLH_X1 \REGISTERS_reg[1][21]  ( .G(n210), .D(n368), .Q(\REGISTERS[1][21] )
         );
  DLH_X1 \REGISTERS_reg[1][20]  ( .G(n210), .D(n372), .Q(\REGISTERS[1][20] )
         );
  DLH_X1 \REGISTERS_reg[1][19]  ( .G(n209), .D(n376), .Q(\REGISTERS[1][19] )
         );
  DLH_X1 \REGISTERS_reg[1][18]  ( .G(n209), .D(n380), .Q(\REGISTERS[1][18] )
         );
  DLH_X1 \REGISTERS_reg[1][17]  ( .G(n209), .D(n384), .Q(\REGISTERS[1][17] )
         );
  DLH_X1 \REGISTERS_reg[1][16]  ( .G(n209), .D(n388), .Q(\REGISTERS[1][16] )
         );
  DLH_X1 \REGISTERS_reg[1][15]  ( .G(n209), .D(n392), .Q(\REGISTERS[1][15] )
         );
  DLH_X1 \REGISTERS_reg[1][14]  ( .G(n209), .D(n396), .Q(\REGISTERS[1][14] )
         );
  DLH_X1 \REGISTERS_reg[1][13]  ( .G(n209), .D(n400), .Q(\REGISTERS[1][13] )
         );
  DLH_X1 \REGISTERS_reg[1][12]  ( .G(n209), .D(n404), .Q(\REGISTERS[1][12] )
         );
  DLH_X1 \REGISTERS_reg[1][11]  ( .G(n209), .D(n408), .Q(\REGISTERS[1][11] )
         );
  DLH_X1 \REGISTERS_reg[1][10]  ( .G(n209), .D(n412), .Q(\REGISTERS[1][10] )
         );
  DLH_X1 \REGISTERS_reg[1][9]  ( .G(n208), .D(n416), .Q(\REGISTERS[1][9] ) );
  DLH_X1 \REGISTERS_reg[1][8]  ( .G(n208), .D(n420), .Q(\REGISTERS[1][8] ) );
  DLH_X1 \REGISTERS_reg[1][7]  ( .G(n208), .D(n424), .Q(\REGISTERS[1][7] ) );
  DLH_X1 \REGISTERS_reg[1][6]  ( .G(n208), .D(n428), .Q(\REGISTERS[1][6] ) );
  DLH_X1 \REGISTERS_reg[1][5]  ( .G(n208), .D(n432), .Q(\REGISTERS[1][5] ) );
  DLH_X1 \REGISTERS_reg[1][4]  ( .G(n208), .D(n436), .Q(\REGISTERS[1][4] ) );
  DLH_X1 \REGISTERS_reg[1][3]  ( .G(n208), .D(n440), .Q(\REGISTERS[1][3] ) );
  DLH_X1 \REGISTERS_reg[1][2]  ( .G(n208), .D(n444), .Q(\REGISTERS[1][2] ) );
  DLH_X1 \REGISTERS_reg[1][1]  ( .G(n208), .D(n448), .Q(\REGISTERS[1][1] ) );
  DLH_X1 \REGISTERS_reg[1][0]  ( .G(n208), .D(n452), .Q(\REGISTERS[1][0] ) );
  DLH_X1 \REGISTERS_reg[2][31]  ( .G(n215), .D(n328), .Q(\REGISTERS[2][31] )
         );
  DLH_X1 \REGISTERS_reg[2][30]  ( .G(n215), .D(n332), .Q(\REGISTERS[2][30] )
         );
  DLH_X1 \REGISTERS_reg[2][29]  ( .G(n214), .D(n336), .Q(\REGISTERS[2][29] )
         );
  DLH_X1 \REGISTERS_reg[2][28]  ( .G(n214), .D(n340), .Q(\REGISTERS[2][28] )
         );
  DLH_X1 \REGISTERS_reg[2][27]  ( .G(n214), .D(n344), .Q(\REGISTERS[2][27] )
         );
  DLH_X1 \REGISTERS_reg[2][26]  ( .G(n214), .D(n348), .Q(\REGISTERS[2][26] )
         );
  DLH_X1 \REGISTERS_reg[2][25]  ( .G(n214), .D(n352), .Q(\REGISTERS[2][25] )
         );
  DLH_X1 \REGISTERS_reg[2][24]  ( .G(n214), .D(n356), .Q(\REGISTERS[2][24] )
         );
  DLH_X1 \REGISTERS_reg[2][23]  ( .G(n214), .D(n360), .Q(\REGISTERS[2][23] )
         );
  DLH_X1 \REGISTERS_reg[2][22]  ( .G(n214), .D(n364), .Q(\REGISTERS[2][22] )
         );
  DLH_X1 \REGISTERS_reg[2][21]  ( .G(n214), .D(n368), .Q(\REGISTERS[2][21] )
         );
  DLH_X1 \REGISTERS_reg[2][20]  ( .G(n214), .D(n372), .Q(\REGISTERS[2][20] )
         );
  DLH_X1 \REGISTERS_reg[2][19]  ( .G(n213), .D(n376), .Q(\REGISTERS[2][19] )
         );
  DLH_X1 \REGISTERS_reg[2][18]  ( .G(n213), .D(n380), .Q(\REGISTERS[2][18] )
         );
  DLH_X1 \REGISTERS_reg[2][17]  ( .G(n213), .D(n384), .Q(\REGISTERS[2][17] )
         );
  DLH_X1 \REGISTERS_reg[2][16]  ( .G(n213), .D(n388), .Q(\REGISTERS[2][16] )
         );
  DLH_X1 \REGISTERS_reg[2][15]  ( .G(n213), .D(n392), .Q(\REGISTERS[2][15] )
         );
  DLH_X1 \REGISTERS_reg[2][14]  ( .G(n213), .D(n396), .Q(\REGISTERS[2][14] )
         );
  DLH_X1 \REGISTERS_reg[2][13]  ( .G(n213), .D(n400), .Q(\REGISTERS[2][13] )
         );
  DLH_X1 \REGISTERS_reg[2][12]  ( .G(n213), .D(n404), .Q(\REGISTERS[2][12] )
         );
  DLH_X1 \REGISTERS_reg[2][11]  ( .G(n213), .D(n408), .Q(\REGISTERS[2][11] )
         );
  DLH_X1 \REGISTERS_reg[2][10]  ( .G(n213), .D(n412), .Q(\REGISTERS[2][10] )
         );
  DLH_X1 \REGISTERS_reg[2][9]  ( .G(n212), .D(n416), .Q(\REGISTERS[2][9] ) );
  DLH_X1 \REGISTERS_reg[2][8]  ( .G(n212), .D(n420), .Q(\REGISTERS[2][8] ) );
  DLH_X1 \REGISTERS_reg[2][7]  ( .G(n212), .D(n424), .Q(\REGISTERS[2][7] ) );
  DLH_X1 \REGISTERS_reg[2][6]  ( .G(n212), .D(n428), .Q(\REGISTERS[2][6] ) );
  DLH_X1 \REGISTERS_reg[2][5]  ( .G(n212), .D(n432), .Q(\REGISTERS[2][5] ) );
  DLH_X1 \REGISTERS_reg[2][4]  ( .G(n212), .D(n436), .Q(\REGISTERS[2][4] ) );
  DLH_X1 \REGISTERS_reg[2][3]  ( .G(n212), .D(n440), .Q(\REGISTERS[2][3] ) );
  DLH_X1 \REGISTERS_reg[2][2]  ( .G(n212), .D(n444), .Q(\REGISTERS[2][2] ) );
  DLH_X1 \REGISTERS_reg[2][1]  ( .G(n212), .D(n448), .Q(\REGISTERS[2][1] ) );
  DLH_X1 \REGISTERS_reg[2][0]  ( .G(n212), .D(n452), .Q(\REGISTERS[2][0] ) );
  DLH_X1 \REGISTERS_reg[3][31]  ( .G(n219), .D(n328), .Q(\REGISTERS[3][31] )
         );
  DLH_X1 \REGISTERS_reg[3][30]  ( .G(n219), .D(n332), .Q(\REGISTERS[3][30] )
         );
  DLH_X1 \REGISTERS_reg[3][29]  ( .G(n218), .D(n336), .Q(\REGISTERS[3][29] )
         );
  DLH_X1 \REGISTERS_reg[3][28]  ( .G(n218), .D(n340), .Q(\REGISTERS[3][28] )
         );
  DLH_X1 \REGISTERS_reg[3][27]  ( .G(n218), .D(n344), .Q(\REGISTERS[3][27] )
         );
  DLH_X1 \REGISTERS_reg[3][26]  ( .G(n218), .D(n348), .Q(\REGISTERS[3][26] )
         );
  DLH_X1 \REGISTERS_reg[3][25]  ( .G(n218), .D(n352), .Q(\REGISTERS[3][25] )
         );
  DLH_X1 \REGISTERS_reg[3][24]  ( .G(n218), .D(n356), .Q(\REGISTERS[3][24] )
         );
  DLH_X1 \REGISTERS_reg[3][23]  ( .G(n218), .D(n360), .Q(\REGISTERS[3][23] )
         );
  DLH_X1 \REGISTERS_reg[3][22]  ( .G(n218), .D(n364), .Q(\REGISTERS[3][22] )
         );
  DLH_X1 \REGISTERS_reg[3][21]  ( .G(n218), .D(n368), .Q(\REGISTERS[3][21] )
         );
  DLH_X1 \REGISTERS_reg[3][20]  ( .G(n218), .D(n372), .Q(\REGISTERS[3][20] )
         );
  DLH_X1 \REGISTERS_reg[3][19]  ( .G(n217), .D(n376), .Q(\REGISTERS[3][19] )
         );
  DLH_X1 \REGISTERS_reg[3][18]  ( .G(n217), .D(n380), .Q(\REGISTERS[3][18] )
         );
  DLH_X1 \REGISTERS_reg[3][17]  ( .G(n217), .D(n384), .Q(\REGISTERS[3][17] )
         );
  DLH_X1 \REGISTERS_reg[3][16]  ( .G(n217), .D(n388), .Q(\REGISTERS[3][16] )
         );
  DLH_X1 \REGISTERS_reg[3][15]  ( .G(n217), .D(n392), .Q(\REGISTERS[3][15] )
         );
  DLH_X1 \REGISTERS_reg[3][14]  ( .G(n217), .D(n396), .Q(\REGISTERS[3][14] )
         );
  DLH_X1 \REGISTERS_reg[3][13]  ( .G(n217), .D(n400), .Q(\REGISTERS[3][13] )
         );
  DLH_X1 \REGISTERS_reg[3][12]  ( .G(n217), .D(n404), .Q(\REGISTERS[3][12] )
         );
  DLH_X1 \REGISTERS_reg[3][11]  ( .G(n217), .D(n408), .Q(\REGISTERS[3][11] )
         );
  DLH_X1 \REGISTERS_reg[3][10]  ( .G(n217), .D(n412), .Q(\REGISTERS[3][10] )
         );
  DLH_X1 \REGISTERS_reg[3][9]  ( .G(n216), .D(n416), .Q(\REGISTERS[3][9] ) );
  DLH_X1 \REGISTERS_reg[3][8]  ( .G(n216), .D(n420), .Q(\REGISTERS[3][8] ) );
  DLH_X1 \REGISTERS_reg[3][7]  ( .G(n216), .D(n424), .Q(\REGISTERS[3][7] ) );
  DLH_X1 \REGISTERS_reg[3][6]  ( .G(n216), .D(n428), .Q(\REGISTERS[3][6] ) );
  DLH_X1 \REGISTERS_reg[3][5]  ( .G(n216), .D(n432), .Q(\REGISTERS[3][5] ) );
  DLH_X1 \REGISTERS_reg[3][4]  ( .G(n216), .D(n436), .Q(\REGISTERS[3][4] ) );
  DLH_X1 \REGISTERS_reg[3][3]  ( .G(n216), .D(n440), .Q(\REGISTERS[3][3] ) );
  DLH_X1 \REGISTERS_reg[3][2]  ( .G(n216), .D(n444), .Q(\REGISTERS[3][2] ) );
  DLH_X1 \REGISTERS_reg[3][1]  ( .G(n216), .D(n448), .Q(\REGISTERS[3][1] ) );
  DLH_X1 \REGISTERS_reg[3][0]  ( .G(n216), .D(n452), .Q(\REGISTERS[3][0] ) );
  DLH_X1 \REGISTERS_reg[4][31]  ( .G(n223), .D(n328), .Q(\REGISTERS[4][31] )
         );
  DLH_X1 \REGISTERS_reg[4][30]  ( .G(n223), .D(n332), .Q(\REGISTERS[4][30] )
         );
  DLH_X1 \REGISTERS_reg[4][29]  ( .G(n222), .D(n336), .Q(\REGISTERS[4][29] )
         );
  DLH_X1 \REGISTERS_reg[4][28]  ( .G(n222), .D(n340), .Q(\REGISTERS[4][28] )
         );
  DLH_X1 \REGISTERS_reg[4][27]  ( .G(n222), .D(n344), .Q(\REGISTERS[4][27] )
         );
  DLH_X1 \REGISTERS_reg[4][26]  ( .G(n222), .D(n348), .Q(\REGISTERS[4][26] )
         );
  DLH_X1 \REGISTERS_reg[4][25]  ( .G(n222), .D(n352), .Q(\REGISTERS[4][25] )
         );
  DLH_X1 \REGISTERS_reg[4][24]  ( .G(n222), .D(n356), .Q(\REGISTERS[4][24] )
         );
  DLH_X1 \REGISTERS_reg[4][23]  ( .G(n222), .D(n360), .Q(\REGISTERS[4][23] )
         );
  DLH_X1 \REGISTERS_reg[4][22]  ( .G(n222), .D(n364), .Q(\REGISTERS[4][22] )
         );
  DLH_X1 \REGISTERS_reg[4][21]  ( .G(n222), .D(n368), .Q(\REGISTERS[4][21] )
         );
  DLH_X1 \REGISTERS_reg[4][20]  ( .G(n222), .D(n372), .Q(\REGISTERS[4][20] )
         );
  DLH_X1 \REGISTERS_reg[4][19]  ( .G(n221), .D(n376), .Q(\REGISTERS[4][19] )
         );
  DLH_X1 \REGISTERS_reg[4][18]  ( .G(n221), .D(n380), .Q(\REGISTERS[4][18] )
         );
  DLH_X1 \REGISTERS_reg[4][17]  ( .G(n221), .D(n384), .Q(\REGISTERS[4][17] )
         );
  DLH_X1 \REGISTERS_reg[4][16]  ( .G(n221), .D(n388), .Q(\REGISTERS[4][16] )
         );
  DLH_X1 \REGISTERS_reg[4][15]  ( .G(n221), .D(n392), .Q(\REGISTERS[4][15] )
         );
  DLH_X1 \REGISTERS_reg[4][14]  ( .G(n221), .D(n396), .Q(\REGISTERS[4][14] )
         );
  DLH_X1 \REGISTERS_reg[4][13]  ( .G(n221), .D(n400), .Q(\REGISTERS[4][13] )
         );
  DLH_X1 \REGISTERS_reg[4][12]  ( .G(n221), .D(n404), .Q(\REGISTERS[4][12] )
         );
  DLH_X1 \REGISTERS_reg[4][11]  ( .G(n221), .D(n408), .Q(\REGISTERS[4][11] )
         );
  DLH_X1 \REGISTERS_reg[4][10]  ( .G(n221), .D(n412), .Q(\REGISTERS[4][10] )
         );
  DLH_X1 \REGISTERS_reg[4][9]  ( .G(n220), .D(n416), .Q(\REGISTERS[4][9] ) );
  DLH_X1 \REGISTERS_reg[4][8]  ( .G(n220), .D(n420), .Q(\REGISTERS[4][8] ) );
  DLH_X1 \REGISTERS_reg[4][7]  ( .G(n220), .D(n424), .Q(\REGISTERS[4][7] ) );
  DLH_X1 \REGISTERS_reg[4][6]  ( .G(n220), .D(n428), .Q(\REGISTERS[4][6] ) );
  DLH_X1 \REGISTERS_reg[4][5]  ( .G(n220), .D(n432), .Q(\REGISTERS[4][5] ) );
  DLH_X1 \REGISTERS_reg[4][4]  ( .G(n220), .D(n436), .Q(\REGISTERS[4][4] ) );
  DLH_X1 \REGISTERS_reg[4][3]  ( .G(n220), .D(n440), .Q(\REGISTERS[4][3] ) );
  DLH_X1 \REGISTERS_reg[4][2]  ( .G(n220), .D(n444), .Q(\REGISTERS[4][2] ) );
  DLH_X1 \REGISTERS_reg[4][1]  ( .G(n220), .D(n448), .Q(\REGISTERS[4][1] ) );
  DLH_X1 \REGISTERS_reg[4][0]  ( .G(n220), .D(n452), .Q(\REGISTERS[4][0] ) );
  DLH_X1 \REGISTERS_reg[5][31]  ( .G(n227), .D(n328), .Q(\REGISTERS[5][31] )
         );
  DLH_X1 \REGISTERS_reg[5][30]  ( .G(n227), .D(n332), .Q(\REGISTERS[5][30] )
         );
  DLH_X1 \REGISTERS_reg[5][29]  ( .G(n226), .D(n336), .Q(\REGISTERS[5][29] )
         );
  DLH_X1 \REGISTERS_reg[5][28]  ( .G(n226), .D(n340), .Q(\REGISTERS[5][28] )
         );
  DLH_X1 \REGISTERS_reg[5][27]  ( .G(n226), .D(n344), .Q(\REGISTERS[5][27] )
         );
  DLH_X1 \REGISTERS_reg[5][26]  ( .G(n226), .D(n348), .Q(\REGISTERS[5][26] )
         );
  DLH_X1 \REGISTERS_reg[5][25]  ( .G(n226), .D(n352), .Q(\REGISTERS[5][25] )
         );
  DLH_X1 \REGISTERS_reg[5][24]  ( .G(n226), .D(n356), .Q(\REGISTERS[5][24] )
         );
  DLH_X1 \REGISTERS_reg[5][23]  ( .G(n226), .D(n360), .Q(\REGISTERS[5][23] )
         );
  DLH_X1 \REGISTERS_reg[5][22]  ( .G(n226), .D(n364), .Q(\REGISTERS[5][22] )
         );
  DLH_X1 \REGISTERS_reg[5][21]  ( .G(n226), .D(n368), .Q(\REGISTERS[5][21] )
         );
  DLH_X1 \REGISTERS_reg[5][20]  ( .G(n226), .D(n372), .Q(\REGISTERS[5][20] )
         );
  DLH_X1 \REGISTERS_reg[5][19]  ( .G(n225), .D(n376), .Q(\REGISTERS[5][19] )
         );
  DLH_X1 \REGISTERS_reg[5][18]  ( .G(n225), .D(n380), .Q(\REGISTERS[5][18] )
         );
  DLH_X1 \REGISTERS_reg[5][17]  ( .G(n225), .D(n384), .Q(\REGISTERS[5][17] )
         );
  DLH_X1 \REGISTERS_reg[5][16]  ( .G(n225), .D(n388), .Q(\REGISTERS[5][16] )
         );
  DLH_X1 \REGISTERS_reg[5][15]  ( .G(n225), .D(n392), .Q(\REGISTERS[5][15] )
         );
  DLH_X1 \REGISTERS_reg[5][14]  ( .G(n225), .D(n396), .Q(\REGISTERS[5][14] )
         );
  DLH_X1 \REGISTERS_reg[5][13]  ( .G(n225), .D(n400), .Q(\REGISTERS[5][13] )
         );
  DLH_X1 \REGISTERS_reg[5][12]  ( .G(n225), .D(n404), .Q(\REGISTERS[5][12] )
         );
  DLH_X1 \REGISTERS_reg[5][11]  ( .G(n225), .D(n408), .Q(\REGISTERS[5][11] )
         );
  DLH_X1 \REGISTERS_reg[5][10]  ( .G(n225), .D(n412), .Q(\REGISTERS[5][10] )
         );
  DLH_X1 \REGISTERS_reg[5][9]  ( .G(n224), .D(n416), .Q(\REGISTERS[5][9] ) );
  DLH_X1 \REGISTERS_reg[5][8]  ( .G(n224), .D(n420), .Q(\REGISTERS[5][8] ) );
  DLH_X1 \REGISTERS_reg[5][7]  ( .G(n224), .D(n424), .Q(\REGISTERS[5][7] ) );
  DLH_X1 \REGISTERS_reg[5][6]  ( .G(n224), .D(n428), .Q(\REGISTERS[5][6] ) );
  DLH_X1 \REGISTERS_reg[5][5]  ( .G(n224), .D(n432), .Q(\REGISTERS[5][5] ) );
  DLH_X1 \REGISTERS_reg[5][4]  ( .G(n224), .D(n436), .Q(\REGISTERS[5][4] ) );
  DLH_X1 \REGISTERS_reg[5][3]  ( .G(n224), .D(n440), .Q(\REGISTERS[5][3] ) );
  DLH_X1 \REGISTERS_reg[5][2]  ( .G(n224), .D(n444), .Q(\REGISTERS[5][2] ) );
  DLH_X1 \REGISTERS_reg[5][1]  ( .G(n224), .D(n448), .Q(\REGISTERS[5][1] ) );
  DLH_X1 \REGISTERS_reg[5][0]  ( .G(n224), .D(n452), .Q(\REGISTERS[5][0] ) );
  DLH_X1 \REGISTERS_reg[6][31]  ( .G(n231), .D(n328), .Q(\REGISTERS[6][31] )
         );
  DLH_X1 \REGISTERS_reg[6][30]  ( .G(n231), .D(n332), .Q(\REGISTERS[6][30] )
         );
  DLH_X1 \REGISTERS_reg[6][29]  ( .G(n230), .D(n336), .Q(\REGISTERS[6][29] )
         );
  DLH_X1 \REGISTERS_reg[6][28]  ( .G(n230), .D(n340), .Q(\REGISTERS[6][28] )
         );
  DLH_X1 \REGISTERS_reg[6][27]  ( .G(n230), .D(n344), .Q(\REGISTERS[6][27] )
         );
  DLH_X1 \REGISTERS_reg[6][26]  ( .G(n230), .D(n348), .Q(\REGISTERS[6][26] )
         );
  DLH_X1 \REGISTERS_reg[6][25]  ( .G(n230), .D(n352), .Q(\REGISTERS[6][25] )
         );
  DLH_X1 \REGISTERS_reg[6][24]  ( .G(n230), .D(n356), .Q(\REGISTERS[6][24] )
         );
  DLH_X1 \REGISTERS_reg[6][23]  ( .G(n230), .D(n360), .Q(\REGISTERS[6][23] )
         );
  DLH_X1 \REGISTERS_reg[6][22]  ( .G(n230), .D(n364), .Q(\REGISTERS[6][22] )
         );
  DLH_X1 \REGISTERS_reg[6][21]  ( .G(n230), .D(n368), .Q(\REGISTERS[6][21] )
         );
  DLH_X1 \REGISTERS_reg[6][20]  ( .G(n230), .D(n372), .Q(\REGISTERS[6][20] )
         );
  DLH_X1 \REGISTERS_reg[6][19]  ( .G(n229), .D(n376), .Q(\REGISTERS[6][19] )
         );
  DLH_X1 \REGISTERS_reg[6][18]  ( .G(n229), .D(n380), .Q(\REGISTERS[6][18] )
         );
  DLH_X1 \REGISTERS_reg[6][17]  ( .G(n229), .D(n384), .Q(\REGISTERS[6][17] )
         );
  DLH_X1 \REGISTERS_reg[6][16]  ( .G(n229), .D(n388), .Q(\REGISTERS[6][16] )
         );
  DLH_X1 \REGISTERS_reg[6][15]  ( .G(n229), .D(n392), .Q(\REGISTERS[6][15] )
         );
  DLH_X1 \REGISTERS_reg[6][14]  ( .G(n229), .D(n396), .Q(\REGISTERS[6][14] )
         );
  DLH_X1 \REGISTERS_reg[6][13]  ( .G(n229), .D(n400), .Q(\REGISTERS[6][13] )
         );
  DLH_X1 \REGISTERS_reg[6][12]  ( .G(n229), .D(n404), .Q(\REGISTERS[6][12] )
         );
  DLH_X1 \REGISTERS_reg[6][11]  ( .G(n229), .D(n408), .Q(\REGISTERS[6][11] )
         );
  DLH_X1 \REGISTERS_reg[6][10]  ( .G(n229), .D(n412), .Q(\REGISTERS[6][10] )
         );
  DLH_X1 \REGISTERS_reg[6][9]  ( .G(n228), .D(n416), .Q(\REGISTERS[6][9] ) );
  DLH_X1 \REGISTERS_reg[6][8]  ( .G(n228), .D(n420), .Q(\REGISTERS[6][8] ) );
  DLH_X1 \REGISTERS_reg[6][7]  ( .G(n228), .D(n424), .Q(\REGISTERS[6][7] ) );
  DLH_X1 \REGISTERS_reg[6][6]  ( .G(n228), .D(n428), .Q(\REGISTERS[6][6] ) );
  DLH_X1 \REGISTERS_reg[6][5]  ( .G(n228), .D(n432), .Q(\REGISTERS[6][5] ) );
  DLH_X1 \REGISTERS_reg[6][4]  ( .G(n228), .D(n436), .Q(\REGISTERS[6][4] ) );
  DLH_X1 \REGISTERS_reg[6][3]  ( .G(n228), .D(n440), .Q(\REGISTERS[6][3] ) );
  DLH_X1 \REGISTERS_reg[6][2]  ( .G(n228), .D(n444), .Q(\REGISTERS[6][2] ) );
  DLH_X1 \REGISTERS_reg[6][1]  ( .G(n228), .D(n448), .Q(\REGISTERS[6][1] ) );
  DLH_X1 \REGISTERS_reg[6][0]  ( .G(n228), .D(n452), .Q(\REGISTERS[6][0] ) );
  DLH_X1 \REGISTERS_reg[7][31]  ( .G(n235), .D(n328), .Q(\REGISTERS[7][31] )
         );
  DLH_X1 \REGISTERS_reg[7][30]  ( .G(n235), .D(n332), .Q(\REGISTERS[7][30] )
         );
  DLH_X1 \REGISTERS_reg[7][29]  ( .G(n234), .D(n336), .Q(\REGISTERS[7][29] )
         );
  DLH_X1 \REGISTERS_reg[7][28]  ( .G(n234), .D(n340), .Q(\REGISTERS[7][28] )
         );
  DLH_X1 \REGISTERS_reg[7][27]  ( .G(n234), .D(n344), .Q(\REGISTERS[7][27] )
         );
  DLH_X1 \REGISTERS_reg[7][26]  ( .G(n234), .D(n348), .Q(\REGISTERS[7][26] )
         );
  DLH_X1 \REGISTERS_reg[7][25]  ( .G(n234), .D(n352), .Q(\REGISTERS[7][25] )
         );
  DLH_X1 \REGISTERS_reg[7][24]  ( .G(n234), .D(n356), .Q(\REGISTERS[7][24] )
         );
  DLH_X1 \REGISTERS_reg[7][23]  ( .G(n234), .D(n360), .Q(\REGISTERS[7][23] )
         );
  DLH_X1 \REGISTERS_reg[7][22]  ( .G(n234), .D(n364), .Q(\REGISTERS[7][22] )
         );
  DLH_X1 \REGISTERS_reg[7][21]  ( .G(n234), .D(n368), .Q(\REGISTERS[7][21] )
         );
  DLH_X1 \REGISTERS_reg[7][20]  ( .G(n234), .D(n372), .Q(\REGISTERS[7][20] )
         );
  DLH_X1 \REGISTERS_reg[7][19]  ( .G(n233), .D(n376), .Q(\REGISTERS[7][19] )
         );
  DLH_X1 \REGISTERS_reg[7][18]  ( .G(n233), .D(n380), .Q(\REGISTERS[7][18] )
         );
  DLH_X1 \REGISTERS_reg[7][17]  ( .G(n233), .D(n384), .Q(\REGISTERS[7][17] )
         );
  DLH_X1 \REGISTERS_reg[7][16]  ( .G(n233), .D(n388), .Q(\REGISTERS[7][16] )
         );
  DLH_X1 \REGISTERS_reg[7][15]  ( .G(n233), .D(n392), .Q(\REGISTERS[7][15] )
         );
  DLH_X1 \REGISTERS_reg[7][14]  ( .G(n233), .D(n396), .Q(\REGISTERS[7][14] )
         );
  DLH_X1 \REGISTERS_reg[7][13]  ( .G(n233), .D(n400), .Q(\REGISTERS[7][13] )
         );
  DLH_X1 \REGISTERS_reg[7][12]  ( .G(n233), .D(n404), .Q(\REGISTERS[7][12] )
         );
  DLH_X1 \REGISTERS_reg[7][11]  ( .G(n233), .D(n408), .Q(\REGISTERS[7][11] )
         );
  DLH_X1 \REGISTERS_reg[7][10]  ( .G(n233), .D(n412), .Q(\REGISTERS[7][10] )
         );
  DLH_X1 \REGISTERS_reg[7][9]  ( .G(n232), .D(n416), .Q(\REGISTERS[7][9] ) );
  DLH_X1 \REGISTERS_reg[7][8]  ( .G(n232), .D(n420), .Q(\REGISTERS[7][8] ) );
  DLH_X1 \REGISTERS_reg[7][7]  ( .G(n232), .D(n424), .Q(\REGISTERS[7][7] ) );
  DLH_X1 \REGISTERS_reg[7][6]  ( .G(n232), .D(n428), .Q(\REGISTERS[7][6] ) );
  DLH_X1 \REGISTERS_reg[7][5]  ( .G(n232), .D(n432), .Q(\REGISTERS[7][5] ) );
  DLH_X1 \REGISTERS_reg[7][4]  ( .G(n232), .D(n436), .Q(\REGISTERS[7][4] ) );
  DLH_X1 \REGISTERS_reg[7][3]  ( .G(n232), .D(n440), .Q(\REGISTERS[7][3] ) );
  DLH_X1 \REGISTERS_reg[7][2]  ( .G(n232), .D(n444), .Q(\REGISTERS[7][2] ) );
  DLH_X1 \REGISTERS_reg[7][1]  ( .G(n232), .D(n448), .Q(\REGISTERS[7][1] ) );
  DLH_X1 \REGISTERS_reg[7][0]  ( .G(n232), .D(n452), .Q(\REGISTERS[7][0] ) );
  DLH_X1 \REGISTERS_reg[8][31]  ( .G(n239), .D(n328), .Q(\REGISTERS[8][31] )
         );
  DLH_X1 \REGISTERS_reg[8][30]  ( .G(n239), .D(n332), .Q(\REGISTERS[8][30] )
         );
  DLH_X1 \REGISTERS_reg[8][29]  ( .G(n238), .D(n336), .Q(\REGISTERS[8][29] )
         );
  DLH_X1 \REGISTERS_reg[8][28]  ( .G(n238), .D(n340), .Q(\REGISTERS[8][28] )
         );
  DLH_X1 \REGISTERS_reg[8][27]  ( .G(n238), .D(n344), .Q(\REGISTERS[8][27] )
         );
  DLH_X1 \REGISTERS_reg[8][26]  ( .G(n238), .D(n348), .Q(\REGISTERS[8][26] )
         );
  DLH_X1 \REGISTERS_reg[8][25]  ( .G(n238), .D(n352), .Q(\REGISTERS[8][25] )
         );
  DLH_X1 \REGISTERS_reg[8][24]  ( .G(n238), .D(n356), .Q(\REGISTERS[8][24] )
         );
  DLH_X1 \REGISTERS_reg[8][23]  ( .G(n238), .D(n360), .Q(\REGISTERS[8][23] )
         );
  DLH_X1 \REGISTERS_reg[8][22]  ( .G(n238), .D(n364), .Q(\REGISTERS[8][22] )
         );
  DLH_X1 \REGISTERS_reg[8][21]  ( .G(n238), .D(n368), .Q(\REGISTERS[8][21] )
         );
  DLH_X1 \REGISTERS_reg[8][20]  ( .G(n238), .D(n372), .Q(\REGISTERS[8][20] )
         );
  DLH_X1 \REGISTERS_reg[8][19]  ( .G(n237), .D(n376), .Q(\REGISTERS[8][19] )
         );
  DLH_X1 \REGISTERS_reg[8][18]  ( .G(n237), .D(n380), .Q(\REGISTERS[8][18] )
         );
  DLH_X1 \REGISTERS_reg[8][17]  ( .G(n237), .D(n384), .Q(\REGISTERS[8][17] )
         );
  DLH_X1 \REGISTERS_reg[8][16]  ( .G(n237), .D(n388), .Q(\REGISTERS[8][16] )
         );
  DLH_X1 \REGISTERS_reg[8][15]  ( .G(n237), .D(n392), .Q(\REGISTERS[8][15] )
         );
  DLH_X1 \REGISTERS_reg[8][14]  ( .G(n237), .D(n396), .Q(\REGISTERS[8][14] )
         );
  DLH_X1 \REGISTERS_reg[8][13]  ( .G(n237), .D(n400), .Q(\REGISTERS[8][13] )
         );
  DLH_X1 \REGISTERS_reg[8][12]  ( .G(n237), .D(n404), .Q(\REGISTERS[8][12] )
         );
  DLH_X1 \REGISTERS_reg[8][11]  ( .G(n237), .D(n408), .Q(\REGISTERS[8][11] )
         );
  DLH_X1 \REGISTERS_reg[8][10]  ( .G(n237), .D(n412), .Q(\REGISTERS[8][10] )
         );
  DLH_X1 \REGISTERS_reg[8][9]  ( .G(n236), .D(n416), .Q(\REGISTERS[8][9] ) );
  DLH_X1 \REGISTERS_reg[8][8]  ( .G(n236), .D(n420), .Q(\REGISTERS[8][8] ) );
  DLH_X1 \REGISTERS_reg[8][7]  ( .G(n236), .D(n424), .Q(\REGISTERS[8][7] ) );
  DLH_X1 \REGISTERS_reg[8][6]  ( .G(n236), .D(n428), .Q(\REGISTERS[8][6] ) );
  DLH_X1 \REGISTERS_reg[8][5]  ( .G(n236), .D(n432), .Q(\REGISTERS[8][5] ) );
  DLH_X1 \REGISTERS_reg[8][4]  ( .G(n236), .D(n436), .Q(\REGISTERS[8][4] ) );
  DLH_X1 \REGISTERS_reg[8][3]  ( .G(n236), .D(n440), .Q(\REGISTERS[8][3] ) );
  DLH_X1 \REGISTERS_reg[8][2]  ( .G(n236), .D(n444), .Q(\REGISTERS[8][2] ) );
  DLH_X1 \REGISTERS_reg[8][1]  ( .G(n236), .D(n448), .Q(\REGISTERS[8][1] ) );
  DLH_X1 \REGISTERS_reg[8][0]  ( .G(n236), .D(n452), .Q(\REGISTERS[8][0] ) );
  DLH_X1 \REGISTERS_reg[9][31]  ( .G(n243), .D(n328), .Q(\REGISTERS[9][31] )
         );
  DLH_X1 \REGISTERS_reg[9][30]  ( .G(n243), .D(n332), .Q(\REGISTERS[9][30] )
         );
  DLH_X1 \REGISTERS_reg[9][29]  ( .G(n242), .D(n336), .Q(\REGISTERS[9][29] )
         );
  DLH_X1 \REGISTERS_reg[9][28]  ( .G(n242), .D(n340), .Q(\REGISTERS[9][28] )
         );
  DLH_X1 \REGISTERS_reg[9][27]  ( .G(n242), .D(n344), .Q(\REGISTERS[9][27] )
         );
  DLH_X1 \REGISTERS_reg[9][26]  ( .G(n242), .D(n348), .Q(\REGISTERS[9][26] )
         );
  DLH_X1 \REGISTERS_reg[9][25]  ( .G(n242), .D(n352), .Q(\REGISTERS[9][25] )
         );
  DLH_X1 \REGISTERS_reg[9][24]  ( .G(n242), .D(n356), .Q(\REGISTERS[9][24] )
         );
  DLH_X1 \REGISTERS_reg[9][23]  ( .G(n242), .D(n360), .Q(\REGISTERS[9][23] )
         );
  DLH_X1 \REGISTERS_reg[9][22]  ( .G(n242), .D(n364), .Q(\REGISTERS[9][22] )
         );
  DLH_X1 \REGISTERS_reg[9][21]  ( .G(n242), .D(n368), .Q(\REGISTERS[9][21] )
         );
  DLH_X1 \REGISTERS_reg[9][20]  ( .G(n242), .D(n372), .Q(\REGISTERS[9][20] )
         );
  DLH_X1 \REGISTERS_reg[9][19]  ( .G(n241), .D(n376), .Q(\REGISTERS[9][19] )
         );
  DLH_X1 \REGISTERS_reg[9][18]  ( .G(n241), .D(n380), .Q(\REGISTERS[9][18] )
         );
  DLH_X1 \REGISTERS_reg[9][17]  ( .G(n241), .D(n384), .Q(\REGISTERS[9][17] )
         );
  DLH_X1 \REGISTERS_reg[9][16]  ( .G(n241), .D(n388), .Q(\REGISTERS[9][16] )
         );
  DLH_X1 \REGISTERS_reg[9][15]  ( .G(n241), .D(n392), .Q(\REGISTERS[9][15] )
         );
  DLH_X1 \REGISTERS_reg[9][14]  ( .G(n241), .D(n396), .Q(\REGISTERS[9][14] )
         );
  DLH_X1 \REGISTERS_reg[9][13]  ( .G(n241), .D(n400), .Q(\REGISTERS[9][13] )
         );
  DLH_X1 \REGISTERS_reg[9][12]  ( .G(n241), .D(n404), .Q(\REGISTERS[9][12] )
         );
  DLH_X1 \REGISTERS_reg[9][11]  ( .G(n241), .D(n408), .Q(\REGISTERS[9][11] )
         );
  DLH_X1 \REGISTERS_reg[9][10]  ( .G(n241), .D(n412), .Q(\REGISTERS[9][10] )
         );
  DLH_X1 \REGISTERS_reg[9][9]  ( .G(n240), .D(n416), .Q(\REGISTERS[9][9] ) );
  DLH_X1 \REGISTERS_reg[9][8]  ( .G(n240), .D(n420), .Q(\REGISTERS[9][8] ) );
  DLH_X1 \REGISTERS_reg[9][7]  ( .G(n240), .D(n424), .Q(\REGISTERS[9][7] ) );
  DLH_X1 \REGISTERS_reg[9][6]  ( .G(n240), .D(n428), .Q(\REGISTERS[9][6] ) );
  DLH_X1 \REGISTERS_reg[9][5]  ( .G(n240), .D(n432), .Q(\REGISTERS[9][5] ) );
  DLH_X1 \REGISTERS_reg[9][4]  ( .G(n240), .D(n436), .Q(\REGISTERS[9][4] ) );
  DLH_X1 \REGISTERS_reg[9][3]  ( .G(n240), .D(n440), .Q(\REGISTERS[9][3] ) );
  DLH_X1 \REGISTERS_reg[9][2]  ( .G(n240), .D(n444), .Q(\REGISTERS[9][2] ) );
  DLH_X1 \REGISTERS_reg[9][1]  ( .G(n240), .D(n448), .Q(\REGISTERS[9][1] ) );
  DLH_X1 \REGISTERS_reg[9][0]  ( .G(n240), .D(n452), .Q(\REGISTERS[9][0] ) );
  DLH_X1 \REGISTERS_reg[10][31]  ( .G(n247), .D(n329), .Q(\REGISTERS[10][31] )
         );
  DLH_X1 \REGISTERS_reg[10][30]  ( .G(n247), .D(n333), .Q(\REGISTERS[10][30] )
         );
  DLH_X1 \REGISTERS_reg[10][29]  ( .G(n246), .D(n337), .Q(\REGISTERS[10][29] )
         );
  DLH_X1 \REGISTERS_reg[10][28]  ( .G(n246), .D(n341), .Q(\REGISTERS[10][28] )
         );
  DLH_X1 \REGISTERS_reg[10][27]  ( .G(n246), .D(n345), .Q(\REGISTERS[10][27] )
         );
  DLH_X1 \REGISTERS_reg[10][26]  ( .G(n246), .D(n349), .Q(\REGISTERS[10][26] )
         );
  DLH_X1 \REGISTERS_reg[10][25]  ( .G(n246), .D(n353), .Q(\REGISTERS[10][25] )
         );
  DLH_X1 \REGISTERS_reg[10][24]  ( .G(n246), .D(n357), .Q(\REGISTERS[10][24] )
         );
  DLH_X1 \REGISTERS_reg[10][23]  ( .G(n246), .D(n361), .Q(\REGISTERS[10][23] )
         );
  DLH_X1 \REGISTERS_reg[10][22]  ( .G(n246), .D(n365), .Q(\REGISTERS[10][22] )
         );
  DLH_X1 \REGISTERS_reg[10][21]  ( .G(n246), .D(n369), .Q(\REGISTERS[10][21] )
         );
  DLH_X1 \REGISTERS_reg[10][20]  ( .G(n246), .D(n373), .Q(\REGISTERS[10][20] )
         );
  DLH_X1 \REGISTERS_reg[10][19]  ( .G(n245), .D(n377), .Q(\REGISTERS[10][19] )
         );
  DLH_X1 \REGISTERS_reg[10][18]  ( .G(n245), .D(n381), .Q(\REGISTERS[10][18] )
         );
  DLH_X1 \REGISTERS_reg[10][17]  ( .G(n245), .D(n385), .Q(\REGISTERS[10][17] )
         );
  DLH_X1 \REGISTERS_reg[10][16]  ( .G(n245), .D(n389), .Q(\REGISTERS[10][16] )
         );
  DLH_X1 \REGISTERS_reg[10][15]  ( .G(n245), .D(n393), .Q(\REGISTERS[10][15] )
         );
  DLH_X1 \REGISTERS_reg[10][14]  ( .G(n245), .D(n397), .Q(\REGISTERS[10][14] )
         );
  DLH_X1 \REGISTERS_reg[10][13]  ( .G(n245), .D(n401), .Q(\REGISTERS[10][13] )
         );
  DLH_X1 \REGISTERS_reg[10][12]  ( .G(n245), .D(n405), .Q(\REGISTERS[10][12] )
         );
  DLH_X1 \REGISTERS_reg[10][11]  ( .G(n245), .D(n409), .Q(\REGISTERS[10][11] )
         );
  DLH_X1 \REGISTERS_reg[10][10]  ( .G(n245), .D(n413), .Q(\REGISTERS[10][10] )
         );
  DLH_X1 \REGISTERS_reg[10][9]  ( .G(n244), .D(n417), .Q(\REGISTERS[10][9] )
         );
  DLH_X1 \REGISTERS_reg[10][8]  ( .G(n244), .D(n421), .Q(\REGISTERS[10][8] )
         );
  DLH_X1 \REGISTERS_reg[10][7]  ( .G(n244), .D(n425), .Q(\REGISTERS[10][7] )
         );
  DLH_X1 \REGISTERS_reg[10][6]  ( .G(n244), .D(n429), .Q(\REGISTERS[10][6] )
         );
  DLH_X1 \REGISTERS_reg[10][5]  ( .G(n244), .D(n433), .Q(\REGISTERS[10][5] )
         );
  DLH_X1 \REGISTERS_reg[10][4]  ( .G(n244), .D(n437), .Q(\REGISTERS[10][4] )
         );
  DLH_X1 \REGISTERS_reg[10][3]  ( .G(n244), .D(n441), .Q(\REGISTERS[10][3] )
         );
  DLH_X1 \REGISTERS_reg[10][2]  ( .G(n244), .D(n445), .Q(\REGISTERS[10][2] )
         );
  DLH_X1 \REGISTERS_reg[10][1]  ( .G(n244), .D(n449), .Q(\REGISTERS[10][1] )
         );
  DLH_X1 \REGISTERS_reg[10][0]  ( .G(n244), .D(n453), .Q(\REGISTERS[10][0] )
         );
  DLH_X1 \REGISTERS_reg[11][31]  ( .G(n251), .D(n329), .Q(\REGISTERS[11][31] )
         );
  DLH_X1 \REGISTERS_reg[11][30]  ( .G(n251), .D(n333), .Q(\REGISTERS[11][30] )
         );
  DLH_X1 \REGISTERS_reg[11][29]  ( .G(n250), .D(n337), .Q(\REGISTERS[11][29] )
         );
  DLH_X1 \REGISTERS_reg[11][28]  ( .G(n250), .D(n341), .Q(\REGISTERS[11][28] )
         );
  DLH_X1 \REGISTERS_reg[11][27]  ( .G(n250), .D(n345), .Q(\REGISTERS[11][27] )
         );
  DLH_X1 \REGISTERS_reg[11][26]  ( .G(n250), .D(n349), .Q(\REGISTERS[11][26] )
         );
  DLH_X1 \REGISTERS_reg[11][25]  ( .G(n250), .D(n353), .Q(\REGISTERS[11][25] )
         );
  DLH_X1 \REGISTERS_reg[11][24]  ( .G(n250), .D(n357), .Q(\REGISTERS[11][24] )
         );
  DLH_X1 \REGISTERS_reg[11][23]  ( .G(n250), .D(n361), .Q(\REGISTERS[11][23] )
         );
  DLH_X1 \REGISTERS_reg[11][22]  ( .G(n250), .D(n365), .Q(\REGISTERS[11][22] )
         );
  DLH_X1 \REGISTERS_reg[11][21]  ( .G(n250), .D(n369), .Q(\REGISTERS[11][21] )
         );
  DLH_X1 \REGISTERS_reg[11][20]  ( .G(n250), .D(n373), .Q(\REGISTERS[11][20] )
         );
  DLH_X1 \REGISTERS_reg[11][19]  ( .G(n249), .D(n377), .Q(\REGISTERS[11][19] )
         );
  DLH_X1 \REGISTERS_reg[11][18]  ( .G(n249), .D(n381), .Q(\REGISTERS[11][18] )
         );
  DLH_X1 \REGISTERS_reg[11][17]  ( .G(n249), .D(n385), .Q(\REGISTERS[11][17] )
         );
  DLH_X1 \REGISTERS_reg[11][16]  ( .G(n249), .D(n389), .Q(\REGISTERS[11][16] )
         );
  DLH_X1 \REGISTERS_reg[11][15]  ( .G(n249), .D(n393), .Q(\REGISTERS[11][15] )
         );
  DLH_X1 \REGISTERS_reg[11][14]  ( .G(n249), .D(n397), .Q(\REGISTERS[11][14] )
         );
  DLH_X1 \REGISTERS_reg[11][13]  ( .G(n249), .D(n401), .Q(\REGISTERS[11][13] )
         );
  DLH_X1 \REGISTERS_reg[11][12]  ( .G(n249), .D(n405), .Q(\REGISTERS[11][12] )
         );
  DLH_X1 \REGISTERS_reg[11][11]  ( .G(n249), .D(n409), .Q(\REGISTERS[11][11] )
         );
  DLH_X1 \REGISTERS_reg[11][10]  ( .G(n249), .D(n413), .Q(\REGISTERS[11][10] )
         );
  DLH_X1 \REGISTERS_reg[11][9]  ( .G(n248), .D(n417), .Q(\REGISTERS[11][9] )
         );
  DLH_X1 \REGISTERS_reg[11][8]  ( .G(n248), .D(n421), .Q(\REGISTERS[11][8] )
         );
  DLH_X1 \REGISTERS_reg[11][7]  ( .G(n248), .D(n425), .Q(\REGISTERS[11][7] )
         );
  DLH_X1 \REGISTERS_reg[11][6]  ( .G(n248), .D(n429), .Q(\REGISTERS[11][6] )
         );
  DLH_X1 \REGISTERS_reg[11][5]  ( .G(n248), .D(n433), .Q(\REGISTERS[11][5] )
         );
  DLH_X1 \REGISTERS_reg[11][4]  ( .G(n248), .D(n437), .Q(\REGISTERS[11][4] )
         );
  DLH_X1 \REGISTERS_reg[11][3]  ( .G(n248), .D(n441), .Q(\REGISTERS[11][3] )
         );
  DLH_X1 \REGISTERS_reg[11][2]  ( .G(n248), .D(n445), .Q(\REGISTERS[11][2] )
         );
  DLH_X1 \REGISTERS_reg[11][1]  ( .G(n248), .D(n449), .Q(\REGISTERS[11][1] )
         );
  DLH_X1 \REGISTERS_reg[11][0]  ( .G(n248), .D(n453), .Q(\REGISTERS[11][0] )
         );
  DLH_X1 \REGISTERS_reg[12][31]  ( .G(n255), .D(n329), .Q(\REGISTERS[12][31] )
         );
  DLH_X1 \REGISTERS_reg[12][30]  ( .G(n255), .D(n333), .Q(\REGISTERS[12][30] )
         );
  DLH_X1 \REGISTERS_reg[12][29]  ( .G(n254), .D(n337), .Q(\REGISTERS[12][29] )
         );
  DLH_X1 \REGISTERS_reg[12][28]  ( .G(n254), .D(n341), .Q(\REGISTERS[12][28] )
         );
  DLH_X1 \REGISTERS_reg[12][27]  ( .G(n254), .D(n345), .Q(\REGISTERS[12][27] )
         );
  DLH_X1 \REGISTERS_reg[12][26]  ( .G(n254), .D(n349), .Q(\REGISTERS[12][26] )
         );
  DLH_X1 \REGISTERS_reg[12][25]  ( .G(n254), .D(n353), .Q(\REGISTERS[12][25] )
         );
  DLH_X1 \REGISTERS_reg[12][24]  ( .G(n254), .D(n357), .Q(\REGISTERS[12][24] )
         );
  DLH_X1 \REGISTERS_reg[12][23]  ( .G(n254), .D(n361), .Q(\REGISTERS[12][23] )
         );
  DLH_X1 \REGISTERS_reg[12][22]  ( .G(n254), .D(n365), .Q(\REGISTERS[12][22] )
         );
  DLH_X1 \REGISTERS_reg[12][21]  ( .G(n254), .D(n369), .Q(\REGISTERS[12][21] )
         );
  DLH_X1 \REGISTERS_reg[12][20]  ( .G(n254), .D(n373), .Q(\REGISTERS[12][20] )
         );
  DLH_X1 \REGISTERS_reg[12][19]  ( .G(n253), .D(n377), .Q(\REGISTERS[12][19] )
         );
  DLH_X1 \REGISTERS_reg[12][18]  ( .G(n253), .D(n381), .Q(\REGISTERS[12][18] )
         );
  DLH_X1 \REGISTERS_reg[12][17]  ( .G(n253), .D(n385), .Q(\REGISTERS[12][17] )
         );
  DLH_X1 \REGISTERS_reg[12][16]  ( .G(n253), .D(n389), .Q(\REGISTERS[12][16] )
         );
  DLH_X1 \REGISTERS_reg[12][15]  ( .G(n253), .D(n393), .Q(\REGISTERS[12][15] )
         );
  DLH_X1 \REGISTERS_reg[12][14]  ( .G(n253), .D(n397), .Q(\REGISTERS[12][14] )
         );
  DLH_X1 \REGISTERS_reg[12][13]  ( .G(n253), .D(n401), .Q(\REGISTERS[12][13] )
         );
  DLH_X1 \REGISTERS_reg[12][12]  ( .G(n253), .D(n405), .Q(\REGISTERS[12][12] )
         );
  DLH_X1 \REGISTERS_reg[12][11]  ( .G(n253), .D(n409), .Q(\REGISTERS[12][11] )
         );
  DLH_X1 \REGISTERS_reg[12][10]  ( .G(n253), .D(n413), .Q(\REGISTERS[12][10] )
         );
  DLH_X1 \REGISTERS_reg[12][9]  ( .G(n252), .D(n417), .Q(\REGISTERS[12][9] )
         );
  DLH_X1 \REGISTERS_reg[12][8]  ( .G(n252), .D(n421), .Q(\REGISTERS[12][8] )
         );
  DLH_X1 \REGISTERS_reg[12][7]  ( .G(n252), .D(n425), .Q(\REGISTERS[12][7] )
         );
  DLH_X1 \REGISTERS_reg[12][6]  ( .G(n252), .D(n429), .Q(\REGISTERS[12][6] )
         );
  DLH_X1 \REGISTERS_reg[12][5]  ( .G(n252), .D(n433), .Q(\REGISTERS[12][5] )
         );
  DLH_X1 \REGISTERS_reg[12][4]  ( .G(n252), .D(n437), .Q(\REGISTERS[12][4] )
         );
  DLH_X1 \REGISTERS_reg[12][3]  ( .G(n252), .D(n441), .Q(\REGISTERS[12][3] )
         );
  DLH_X1 \REGISTERS_reg[12][2]  ( .G(n252), .D(n445), .Q(\REGISTERS[12][2] )
         );
  DLH_X1 \REGISTERS_reg[12][1]  ( .G(n252), .D(n449), .Q(\REGISTERS[12][1] )
         );
  DLH_X1 \REGISTERS_reg[12][0]  ( .G(n252), .D(n453), .Q(\REGISTERS[12][0] )
         );
  DLH_X1 \REGISTERS_reg[13][31]  ( .G(n259), .D(n329), .Q(\REGISTERS[13][31] )
         );
  DLH_X1 \REGISTERS_reg[13][30]  ( .G(n259), .D(n333), .Q(\REGISTERS[13][30] )
         );
  DLH_X1 \REGISTERS_reg[13][29]  ( .G(n258), .D(n337), .Q(\REGISTERS[13][29] )
         );
  DLH_X1 \REGISTERS_reg[13][28]  ( .G(n258), .D(n341), .Q(\REGISTERS[13][28] )
         );
  DLH_X1 \REGISTERS_reg[13][27]  ( .G(n258), .D(n345), .Q(\REGISTERS[13][27] )
         );
  DLH_X1 \REGISTERS_reg[13][26]  ( .G(n258), .D(n349), .Q(\REGISTERS[13][26] )
         );
  DLH_X1 \REGISTERS_reg[13][25]  ( .G(n258), .D(n353), .Q(\REGISTERS[13][25] )
         );
  DLH_X1 \REGISTERS_reg[13][24]  ( .G(n258), .D(n357), .Q(\REGISTERS[13][24] )
         );
  DLH_X1 \REGISTERS_reg[13][23]  ( .G(n258), .D(n361), .Q(\REGISTERS[13][23] )
         );
  DLH_X1 \REGISTERS_reg[13][22]  ( .G(n258), .D(n365), .Q(\REGISTERS[13][22] )
         );
  DLH_X1 \REGISTERS_reg[13][21]  ( .G(n258), .D(n369), .Q(\REGISTERS[13][21] )
         );
  DLH_X1 \REGISTERS_reg[13][20]  ( .G(n258), .D(n373), .Q(\REGISTERS[13][20] )
         );
  DLH_X1 \REGISTERS_reg[13][19]  ( .G(n257), .D(n377), .Q(\REGISTERS[13][19] )
         );
  DLH_X1 \REGISTERS_reg[13][18]  ( .G(n257), .D(n381), .Q(\REGISTERS[13][18] )
         );
  DLH_X1 \REGISTERS_reg[13][17]  ( .G(n257), .D(n385), .Q(\REGISTERS[13][17] )
         );
  DLH_X1 \REGISTERS_reg[13][16]  ( .G(n257), .D(n389), .Q(\REGISTERS[13][16] )
         );
  DLH_X1 \REGISTERS_reg[13][15]  ( .G(n257), .D(n393), .Q(\REGISTERS[13][15] )
         );
  DLH_X1 \REGISTERS_reg[13][14]  ( .G(n257), .D(n397), .Q(\REGISTERS[13][14] )
         );
  DLH_X1 \REGISTERS_reg[13][13]  ( .G(n257), .D(n401), .Q(\REGISTERS[13][13] )
         );
  DLH_X1 \REGISTERS_reg[13][12]  ( .G(n257), .D(n405), .Q(\REGISTERS[13][12] )
         );
  DLH_X1 \REGISTERS_reg[13][11]  ( .G(n257), .D(n409), .Q(\REGISTERS[13][11] )
         );
  DLH_X1 \REGISTERS_reg[13][10]  ( .G(n257), .D(n413), .Q(\REGISTERS[13][10] )
         );
  DLH_X1 \REGISTERS_reg[13][9]  ( .G(n256), .D(n417), .Q(\REGISTERS[13][9] )
         );
  DLH_X1 \REGISTERS_reg[13][8]  ( .G(n256), .D(n421), .Q(\REGISTERS[13][8] )
         );
  DLH_X1 \REGISTERS_reg[13][7]  ( .G(n256), .D(n425), .Q(\REGISTERS[13][7] )
         );
  DLH_X1 \REGISTERS_reg[13][6]  ( .G(n256), .D(n429), .Q(\REGISTERS[13][6] )
         );
  DLH_X1 \REGISTERS_reg[13][5]  ( .G(n256), .D(n433), .Q(\REGISTERS[13][5] )
         );
  DLH_X1 \REGISTERS_reg[13][4]  ( .G(n256), .D(n437), .Q(\REGISTERS[13][4] )
         );
  DLH_X1 \REGISTERS_reg[13][3]  ( .G(n256), .D(n441), .Q(\REGISTERS[13][3] )
         );
  DLH_X1 \REGISTERS_reg[13][2]  ( .G(n256), .D(n445), .Q(\REGISTERS[13][2] )
         );
  DLH_X1 \REGISTERS_reg[13][1]  ( .G(n256), .D(n449), .Q(\REGISTERS[13][1] )
         );
  DLH_X1 \REGISTERS_reg[13][0]  ( .G(n256), .D(n453), .Q(\REGISTERS[13][0] )
         );
  DLH_X1 \REGISTERS_reg[14][31]  ( .G(n263), .D(n329), .Q(\REGISTERS[14][31] )
         );
  DLH_X1 \REGISTERS_reg[14][30]  ( .G(n263), .D(n333), .Q(\REGISTERS[14][30] )
         );
  DLH_X1 \REGISTERS_reg[14][29]  ( .G(n262), .D(n337), .Q(\REGISTERS[14][29] )
         );
  DLH_X1 \REGISTERS_reg[14][28]  ( .G(n262), .D(n341), .Q(\REGISTERS[14][28] )
         );
  DLH_X1 \REGISTERS_reg[14][27]  ( .G(n262), .D(n345), .Q(\REGISTERS[14][27] )
         );
  DLH_X1 \REGISTERS_reg[14][26]  ( .G(n262), .D(n349), .Q(\REGISTERS[14][26] )
         );
  DLH_X1 \REGISTERS_reg[14][25]  ( .G(n262), .D(n353), .Q(\REGISTERS[14][25] )
         );
  DLH_X1 \REGISTERS_reg[14][24]  ( .G(n262), .D(n357), .Q(\REGISTERS[14][24] )
         );
  DLH_X1 \REGISTERS_reg[14][23]  ( .G(n262), .D(n361), .Q(\REGISTERS[14][23] )
         );
  DLH_X1 \REGISTERS_reg[14][22]  ( .G(n262), .D(n365), .Q(\REGISTERS[14][22] )
         );
  DLH_X1 \REGISTERS_reg[14][21]  ( .G(n262), .D(n369), .Q(\REGISTERS[14][21] )
         );
  DLH_X1 \REGISTERS_reg[14][20]  ( .G(n262), .D(n373), .Q(\REGISTERS[14][20] )
         );
  DLH_X1 \REGISTERS_reg[14][19]  ( .G(n261), .D(n377), .Q(\REGISTERS[14][19] )
         );
  DLH_X1 \REGISTERS_reg[14][18]  ( .G(n261), .D(n381), .Q(\REGISTERS[14][18] )
         );
  DLH_X1 \REGISTERS_reg[14][17]  ( .G(n261), .D(n385), .Q(\REGISTERS[14][17] )
         );
  DLH_X1 \REGISTERS_reg[14][16]  ( .G(n261), .D(n389), .Q(\REGISTERS[14][16] )
         );
  DLH_X1 \REGISTERS_reg[14][15]  ( .G(n261), .D(n393), .Q(\REGISTERS[14][15] )
         );
  DLH_X1 \REGISTERS_reg[14][14]  ( .G(n261), .D(n397), .Q(\REGISTERS[14][14] )
         );
  DLH_X1 \REGISTERS_reg[14][13]  ( .G(n261), .D(n401), .Q(\REGISTERS[14][13] )
         );
  DLH_X1 \REGISTERS_reg[14][12]  ( .G(n261), .D(n405), .Q(\REGISTERS[14][12] )
         );
  DLH_X1 \REGISTERS_reg[14][11]  ( .G(n261), .D(n409), .Q(\REGISTERS[14][11] )
         );
  DLH_X1 \REGISTERS_reg[14][10]  ( .G(n261), .D(n413), .Q(\REGISTERS[14][10] )
         );
  DLH_X1 \REGISTERS_reg[14][9]  ( .G(n260), .D(n417), .Q(\REGISTERS[14][9] )
         );
  DLH_X1 \REGISTERS_reg[14][8]  ( .G(n260), .D(n421), .Q(\REGISTERS[14][8] )
         );
  DLH_X1 \REGISTERS_reg[14][7]  ( .G(n260), .D(n425), .Q(\REGISTERS[14][7] )
         );
  DLH_X1 \REGISTERS_reg[14][6]  ( .G(n260), .D(n429), .Q(\REGISTERS[14][6] )
         );
  DLH_X1 \REGISTERS_reg[14][5]  ( .G(n260), .D(n433), .Q(\REGISTERS[14][5] )
         );
  DLH_X1 \REGISTERS_reg[14][4]  ( .G(n260), .D(n437), .Q(\REGISTERS[14][4] )
         );
  DLH_X1 \REGISTERS_reg[14][3]  ( .G(n260), .D(n441), .Q(\REGISTERS[14][3] )
         );
  DLH_X1 \REGISTERS_reg[14][2]  ( .G(n260), .D(n445), .Q(\REGISTERS[14][2] )
         );
  DLH_X1 \REGISTERS_reg[14][1]  ( .G(n260), .D(n449), .Q(\REGISTERS[14][1] )
         );
  DLH_X1 \REGISTERS_reg[14][0]  ( .G(n260), .D(n453), .Q(\REGISTERS[14][0] )
         );
  DLH_X1 \REGISTERS_reg[15][31]  ( .G(n267), .D(n329), .Q(\REGISTERS[15][31] )
         );
  DLH_X1 \REGISTERS_reg[15][30]  ( .G(n267), .D(n333), .Q(\REGISTERS[15][30] )
         );
  DLH_X1 \REGISTERS_reg[15][29]  ( .G(n266), .D(n337), .Q(\REGISTERS[15][29] )
         );
  DLH_X1 \REGISTERS_reg[15][28]  ( .G(n266), .D(n341), .Q(\REGISTERS[15][28] )
         );
  DLH_X1 \REGISTERS_reg[15][27]  ( .G(n266), .D(n345), .Q(\REGISTERS[15][27] )
         );
  DLH_X1 \REGISTERS_reg[15][26]  ( .G(n266), .D(n349), .Q(\REGISTERS[15][26] )
         );
  DLH_X1 \REGISTERS_reg[15][25]  ( .G(n266), .D(n353), .Q(\REGISTERS[15][25] )
         );
  DLH_X1 \REGISTERS_reg[15][24]  ( .G(n266), .D(n357), .Q(\REGISTERS[15][24] )
         );
  DLH_X1 \REGISTERS_reg[15][23]  ( .G(n266), .D(n361), .Q(\REGISTERS[15][23] )
         );
  DLH_X1 \REGISTERS_reg[15][22]  ( .G(n266), .D(n365), .Q(\REGISTERS[15][22] )
         );
  DLH_X1 \REGISTERS_reg[15][21]  ( .G(n266), .D(n369), .Q(\REGISTERS[15][21] )
         );
  DLH_X1 \REGISTERS_reg[15][20]  ( .G(n266), .D(n373), .Q(\REGISTERS[15][20] )
         );
  DLH_X1 \REGISTERS_reg[15][19]  ( .G(n265), .D(n377), .Q(\REGISTERS[15][19] )
         );
  DLH_X1 \REGISTERS_reg[15][18]  ( .G(n265), .D(n381), .Q(\REGISTERS[15][18] )
         );
  DLH_X1 \REGISTERS_reg[15][17]  ( .G(n265), .D(n385), .Q(\REGISTERS[15][17] )
         );
  DLH_X1 \REGISTERS_reg[15][16]  ( .G(n265), .D(n389), .Q(\REGISTERS[15][16] )
         );
  DLH_X1 \REGISTERS_reg[15][15]  ( .G(n265), .D(n393), .Q(\REGISTERS[15][15] )
         );
  DLH_X1 \REGISTERS_reg[15][14]  ( .G(n265), .D(n397), .Q(\REGISTERS[15][14] )
         );
  DLH_X1 \REGISTERS_reg[15][13]  ( .G(n265), .D(n401), .Q(\REGISTERS[15][13] )
         );
  DLH_X1 \REGISTERS_reg[15][12]  ( .G(n265), .D(n405), .Q(\REGISTERS[15][12] )
         );
  DLH_X1 \REGISTERS_reg[15][11]  ( .G(n265), .D(n409), .Q(\REGISTERS[15][11] )
         );
  DLH_X1 \REGISTERS_reg[15][10]  ( .G(n265), .D(n413), .Q(\REGISTERS[15][10] )
         );
  DLH_X1 \REGISTERS_reg[15][9]  ( .G(n264), .D(n417), .Q(\REGISTERS[15][9] )
         );
  DLH_X1 \REGISTERS_reg[15][8]  ( .G(n264), .D(n421), .Q(\REGISTERS[15][8] )
         );
  DLH_X1 \REGISTERS_reg[15][7]  ( .G(n264), .D(n425), .Q(\REGISTERS[15][7] )
         );
  DLH_X1 \REGISTERS_reg[15][6]  ( .G(n264), .D(n429), .Q(\REGISTERS[15][6] )
         );
  DLH_X1 \REGISTERS_reg[15][5]  ( .G(n264), .D(n433), .Q(\REGISTERS[15][5] )
         );
  DLH_X1 \REGISTERS_reg[15][4]  ( .G(n264), .D(n437), .Q(\REGISTERS[15][4] )
         );
  DLH_X1 \REGISTERS_reg[15][3]  ( .G(n264), .D(n441), .Q(\REGISTERS[15][3] )
         );
  DLH_X1 \REGISTERS_reg[15][2]  ( .G(n264), .D(n445), .Q(\REGISTERS[15][2] )
         );
  DLH_X1 \REGISTERS_reg[15][1]  ( .G(n264), .D(n449), .Q(\REGISTERS[15][1] )
         );
  DLH_X1 \REGISTERS_reg[15][0]  ( .G(n264), .D(n453), .Q(\REGISTERS[15][0] )
         );
  DLH_X1 \REGISTERS_reg[16][31]  ( .G(n271), .D(n329), .Q(\REGISTERS[16][31] )
         );
  DLH_X1 \REGISTERS_reg[16][30]  ( .G(n271), .D(n333), .Q(\REGISTERS[16][30] )
         );
  DLH_X1 \REGISTERS_reg[16][29]  ( .G(n270), .D(n337), .Q(\REGISTERS[16][29] )
         );
  DLH_X1 \REGISTERS_reg[16][28]  ( .G(n270), .D(n341), .Q(\REGISTERS[16][28] )
         );
  DLH_X1 \REGISTERS_reg[16][27]  ( .G(n270), .D(n345), .Q(\REGISTERS[16][27] )
         );
  DLH_X1 \REGISTERS_reg[16][26]  ( .G(n270), .D(n349), .Q(\REGISTERS[16][26] )
         );
  DLH_X1 \REGISTERS_reg[16][25]  ( .G(n270), .D(n353), .Q(\REGISTERS[16][25] )
         );
  DLH_X1 \REGISTERS_reg[16][24]  ( .G(n270), .D(n357), .Q(\REGISTERS[16][24] )
         );
  DLH_X1 \REGISTERS_reg[16][23]  ( .G(n270), .D(n361), .Q(\REGISTERS[16][23] )
         );
  DLH_X1 \REGISTERS_reg[16][22]  ( .G(n270), .D(n365), .Q(\REGISTERS[16][22] )
         );
  DLH_X1 \REGISTERS_reg[16][21]  ( .G(n270), .D(n369), .Q(\REGISTERS[16][21] )
         );
  DLH_X1 \REGISTERS_reg[16][20]  ( .G(n270), .D(n373), .Q(\REGISTERS[16][20] )
         );
  DLH_X1 \REGISTERS_reg[16][19]  ( .G(n269), .D(n377), .Q(\REGISTERS[16][19] )
         );
  DLH_X1 \REGISTERS_reg[16][18]  ( .G(n269), .D(n381), .Q(\REGISTERS[16][18] )
         );
  DLH_X1 \REGISTERS_reg[16][17]  ( .G(n269), .D(n385), .Q(\REGISTERS[16][17] )
         );
  DLH_X1 \REGISTERS_reg[16][16]  ( .G(n269), .D(n389), .Q(\REGISTERS[16][16] )
         );
  DLH_X1 \REGISTERS_reg[16][15]  ( .G(n269), .D(n393), .Q(\REGISTERS[16][15] )
         );
  DLH_X1 \REGISTERS_reg[16][14]  ( .G(n269), .D(n397), .Q(\REGISTERS[16][14] )
         );
  DLH_X1 \REGISTERS_reg[16][13]  ( .G(n269), .D(n401), .Q(\REGISTERS[16][13] )
         );
  DLH_X1 \REGISTERS_reg[16][12]  ( .G(n269), .D(n405), .Q(\REGISTERS[16][12] )
         );
  DLH_X1 \REGISTERS_reg[16][11]  ( .G(n269), .D(n409), .Q(\REGISTERS[16][11] )
         );
  DLH_X1 \REGISTERS_reg[16][10]  ( .G(n269), .D(n413), .Q(\REGISTERS[16][10] )
         );
  DLH_X1 \REGISTERS_reg[16][9]  ( .G(n268), .D(n417), .Q(\REGISTERS[16][9] )
         );
  DLH_X1 \REGISTERS_reg[16][8]  ( .G(n268), .D(n421), .Q(\REGISTERS[16][8] )
         );
  DLH_X1 \REGISTERS_reg[16][7]  ( .G(n268), .D(n425), .Q(\REGISTERS[16][7] )
         );
  DLH_X1 \REGISTERS_reg[16][6]  ( .G(n268), .D(n429), .Q(\REGISTERS[16][6] )
         );
  DLH_X1 \REGISTERS_reg[16][5]  ( .G(n268), .D(n433), .Q(\REGISTERS[16][5] )
         );
  DLH_X1 \REGISTERS_reg[16][4]  ( .G(n268), .D(n437), .Q(\REGISTERS[16][4] )
         );
  DLH_X1 \REGISTERS_reg[16][3]  ( .G(n268), .D(n441), .Q(\REGISTERS[16][3] )
         );
  DLH_X1 \REGISTERS_reg[16][2]  ( .G(n268), .D(n445), .Q(\REGISTERS[16][2] )
         );
  DLH_X1 \REGISTERS_reg[16][1]  ( .G(n268), .D(n449), .Q(\REGISTERS[16][1] )
         );
  DLH_X1 \REGISTERS_reg[16][0]  ( .G(n268), .D(n453), .Q(\REGISTERS[16][0] )
         );
  DLH_X1 \REGISTERS_reg[17][31]  ( .G(n275), .D(n329), .Q(\REGISTERS[17][31] )
         );
  DLH_X1 \REGISTERS_reg[17][30]  ( .G(n275), .D(n333), .Q(\REGISTERS[17][30] )
         );
  DLH_X1 \REGISTERS_reg[17][29]  ( .G(n274), .D(n337), .Q(\REGISTERS[17][29] )
         );
  DLH_X1 \REGISTERS_reg[17][28]  ( .G(n274), .D(n341), .Q(\REGISTERS[17][28] )
         );
  DLH_X1 \REGISTERS_reg[17][27]  ( .G(n274), .D(n345), .Q(\REGISTERS[17][27] )
         );
  DLH_X1 \REGISTERS_reg[17][26]  ( .G(n274), .D(n349), .Q(\REGISTERS[17][26] )
         );
  DLH_X1 \REGISTERS_reg[17][25]  ( .G(n274), .D(n353), .Q(\REGISTERS[17][25] )
         );
  DLH_X1 \REGISTERS_reg[17][24]  ( .G(n274), .D(n357), .Q(\REGISTERS[17][24] )
         );
  DLH_X1 \REGISTERS_reg[17][23]  ( .G(n274), .D(n361), .Q(\REGISTERS[17][23] )
         );
  DLH_X1 \REGISTERS_reg[17][22]  ( .G(n274), .D(n365), .Q(\REGISTERS[17][22] )
         );
  DLH_X1 \REGISTERS_reg[17][21]  ( .G(n274), .D(n369), .Q(\REGISTERS[17][21] )
         );
  DLH_X1 \REGISTERS_reg[17][20]  ( .G(n274), .D(n373), .Q(\REGISTERS[17][20] )
         );
  DLH_X1 \REGISTERS_reg[17][19]  ( .G(n273), .D(n377), .Q(\REGISTERS[17][19] )
         );
  DLH_X1 \REGISTERS_reg[17][18]  ( .G(n273), .D(n381), .Q(\REGISTERS[17][18] )
         );
  DLH_X1 \REGISTERS_reg[17][17]  ( .G(n273), .D(n385), .Q(\REGISTERS[17][17] )
         );
  DLH_X1 \REGISTERS_reg[17][16]  ( .G(n273), .D(n389), .Q(\REGISTERS[17][16] )
         );
  DLH_X1 \REGISTERS_reg[17][15]  ( .G(n273), .D(n393), .Q(\REGISTERS[17][15] )
         );
  DLH_X1 \REGISTERS_reg[17][14]  ( .G(n273), .D(n397), .Q(\REGISTERS[17][14] )
         );
  DLH_X1 \REGISTERS_reg[17][13]  ( .G(n273), .D(n401), .Q(\REGISTERS[17][13] )
         );
  DLH_X1 \REGISTERS_reg[17][12]  ( .G(n273), .D(n405), .Q(\REGISTERS[17][12] )
         );
  DLH_X1 \REGISTERS_reg[17][11]  ( .G(n273), .D(n409), .Q(\REGISTERS[17][11] )
         );
  DLH_X1 \REGISTERS_reg[17][10]  ( .G(n273), .D(n413), .Q(\REGISTERS[17][10] )
         );
  DLH_X1 \REGISTERS_reg[17][9]  ( .G(n272), .D(n417), .Q(\REGISTERS[17][9] )
         );
  DLH_X1 \REGISTERS_reg[17][8]  ( .G(n272), .D(n421), .Q(\REGISTERS[17][8] )
         );
  DLH_X1 \REGISTERS_reg[17][7]  ( .G(n272), .D(n425), .Q(\REGISTERS[17][7] )
         );
  DLH_X1 \REGISTERS_reg[17][6]  ( .G(n272), .D(n429), .Q(\REGISTERS[17][6] )
         );
  DLH_X1 \REGISTERS_reg[17][5]  ( .G(n272), .D(n433), .Q(\REGISTERS[17][5] )
         );
  DLH_X1 \REGISTERS_reg[17][4]  ( .G(n272), .D(n437), .Q(\REGISTERS[17][4] )
         );
  DLH_X1 \REGISTERS_reg[17][3]  ( .G(n272), .D(n441), .Q(\REGISTERS[17][3] )
         );
  DLH_X1 \REGISTERS_reg[17][2]  ( .G(n272), .D(n445), .Q(\REGISTERS[17][2] )
         );
  DLH_X1 \REGISTERS_reg[17][1]  ( .G(n272), .D(n449), .Q(\REGISTERS[17][1] )
         );
  DLH_X1 \REGISTERS_reg[17][0]  ( .G(n272), .D(n453), .Q(\REGISTERS[17][0] )
         );
  DLH_X1 \REGISTERS_reg[18][31]  ( .G(n279), .D(n329), .Q(\REGISTERS[18][31] )
         );
  DLH_X1 \REGISTERS_reg[18][30]  ( .G(n279), .D(n333), .Q(\REGISTERS[18][30] )
         );
  DLH_X1 \REGISTERS_reg[18][29]  ( .G(n278), .D(n337), .Q(\REGISTERS[18][29] )
         );
  DLH_X1 \REGISTERS_reg[18][28]  ( .G(n278), .D(n341), .Q(\REGISTERS[18][28] )
         );
  DLH_X1 \REGISTERS_reg[18][27]  ( .G(n278), .D(n345), .Q(\REGISTERS[18][27] )
         );
  DLH_X1 \REGISTERS_reg[18][26]  ( .G(n278), .D(n349), .Q(\REGISTERS[18][26] )
         );
  DLH_X1 \REGISTERS_reg[18][25]  ( .G(n278), .D(n353), .Q(\REGISTERS[18][25] )
         );
  DLH_X1 \REGISTERS_reg[18][24]  ( .G(n278), .D(n357), .Q(\REGISTERS[18][24] )
         );
  DLH_X1 \REGISTERS_reg[18][23]  ( .G(n278), .D(n361), .Q(\REGISTERS[18][23] )
         );
  DLH_X1 \REGISTERS_reg[18][22]  ( .G(n278), .D(n365), .Q(\REGISTERS[18][22] )
         );
  DLH_X1 \REGISTERS_reg[18][21]  ( .G(n278), .D(n369), .Q(\REGISTERS[18][21] )
         );
  DLH_X1 \REGISTERS_reg[18][20]  ( .G(n278), .D(n373), .Q(\REGISTERS[18][20] )
         );
  DLH_X1 \REGISTERS_reg[18][19]  ( .G(n277), .D(n377), .Q(\REGISTERS[18][19] )
         );
  DLH_X1 \REGISTERS_reg[18][18]  ( .G(n277), .D(n381), .Q(\REGISTERS[18][18] )
         );
  DLH_X1 \REGISTERS_reg[18][17]  ( .G(n277), .D(n385), .Q(\REGISTERS[18][17] )
         );
  DLH_X1 \REGISTERS_reg[18][16]  ( .G(n277), .D(n389), .Q(\REGISTERS[18][16] )
         );
  DLH_X1 \REGISTERS_reg[18][15]  ( .G(n277), .D(n393), .Q(\REGISTERS[18][15] )
         );
  DLH_X1 \REGISTERS_reg[18][14]  ( .G(n277), .D(n397), .Q(\REGISTERS[18][14] )
         );
  DLH_X1 \REGISTERS_reg[18][13]  ( .G(n277), .D(n401), .Q(\REGISTERS[18][13] )
         );
  DLH_X1 \REGISTERS_reg[18][12]  ( .G(n277), .D(n405), .Q(\REGISTERS[18][12] )
         );
  DLH_X1 \REGISTERS_reg[18][11]  ( .G(n277), .D(n409), .Q(\REGISTERS[18][11] )
         );
  DLH_X1 \REGISTERS_reg[18][10]  ( .G(n277), .D(n413), .Q(\REGISTERS[18][10] )
         );
  DLH_X1 \REGISTERS_reg[18][9]  ( .G(n276), .D(n417), .Q(\REGISTERS[18][9] )
         );
  DLH_X1 \REGISTERS_reg[18][8]  ( .G(n276), .D(n421), .Q(\REGISTERS[18][8] )
         );
  DLH_X1 \REGISTERS_reg[18][7]  ( .G(n276), .D(n425), .Q(\REGISTERS[18][7] )
         );
  DLH_X1 \REGISTERS_reg[18][6]  ( .G(n276), .D(n429), .Q(\REGISTERS[18][6] )
         );
  DLH_X1 \REGISTERS_reg[18][5]  ( .G(n276), .D(n433), .Q(\REGISTERS[18][5] )
         );
  DLH_X1 \REGISTERS_reg[18][4]  ( .G(n276), .D(n437), .Q(\REGISTERS[18][4] )
         );
  DLH_X1 \REGISTERS_reg[18][3]  ( .G(n276), .D(n441), .Q(\REGISTERS[18][3] )
         );
  DLH_X1 \REGISTERS_reg[18][2]  ( .G(n276), .D(n445), .Q(\REGISTERS[18][2] )
         );
  DLH_X1 \REGISTERS_reg[18][1]  ( .G(n276), .D(n449), .Q(\REGISTERS[18][1] )
         );
  DLH_X1 \REGISTERS_reg[18][0]  ( .G(n276), .D(n453), .Q(\REGISTERS[18][0] )
         );
  DLH_X1 \REGISTERS_reg[19][31]  ( .G(n283), .D(n329), .Q(\REGISTERS[19][31] )
         );
  DLH_X1 \REGISTERS_reg[19][30]  ( .G(n283), .D(n333), .Q(\REGISTERS[19][30] )
         );
  DLH_X1 \REGISTERS_reg[19][29]  ( .G(n282), .D(n337), .Q(\REGISTERS[19][29] )
         );
  DLH_X1 \REGISTERS_reg[19][28]  ( .G(n282), .D(n341), .Q(\REGISTERS[19][28] )
         );
  DLH_X1 \REGISTERS_reg[19][27]  ( .G(n282), .D(n345), .Q(\REGISTERS[19][27] )
         );
  DLH_X1 \REGISTERS_reg[19][26]  ( .G(n282), .D(n349), .Q(\REGISTERS[19][26] )
         );
  DLH_X1 \REGISTERS_reg[19][25]  ( .G(n282), .D(n353), .Q(\REGISTERS[19][25] )
         );
  DLH_X1 \REGISTERS_reg[19][24]  ( .G(n282), .D(n357), .Q(\REGISTERS[19][24] )
         );
  DLH_X1 \REGISTERS_reg[19][23]  ( .G(n282), .D(n361), .Q(\REGISTERS[19][23] )
         );
  DLH_X1 \REGISTERS_reg[19][22]  ( .G(n282), .D(n365), .Q(\REGISTERS[19][22] )
         );
  DLH_X1 \REGISTERS_reg[19][21]  ( .G(n282), .D(n369), .Q(\REGISTERS[19][21] )
         );
  DLH_X1 \REGISTERS_reg[19][20]  ( .G(n282), .D(n373), .Q(\REGISTERS[19][20] )
         );
  DLH_X1 \REGISTERS_reg[19][19]  ( .G(n281), .D(n377), .Q(\REGISTERS[19][19] )
         );
  DLH_X1 \REGISTERS_reg[19][18]  ( .G(n281), .D(n381), .Q(\REGISTERS[19][18] )
         );
  DLH_X1 \REGISTERS_reg[19][17]  ( .G(n281), .D(n385), .Q(\REGISTERS[19][17] )
         );
  DLH_X1 \REGISTERS_reg[19][16]  ( .G(n281), .D(n389), .Q(\REGISTERS[19][16] )
         );
  DLH_X1 \REGISTERS_reg[19][15]  ( .G(n281), .D(n393), .Q(\REGISTERS[19][15] )
         );
  DLH_X1 \REGISTERS_reg[19][14]  ( .G(n281), .D(n397), .Q(\REGISTERS[19][14] )
         );
  DLH_X1 \REGISTERS_reg[19][13]  ( .G(n281), .D(n401), .Q(\REGISTERS[19][13] )
         );
  DLH_X1 \REGISTERS_reg[19][12]  ( .G(n281), .D(n405), .Q(\REGISTERS[19][12] )
         );
  DLH_X1 \REGISTERS_reg[19][11]  ( .G(n281), .D(n409), .Q(\REGISTERS[19][11] )
         );
  DLH_X1 \REGISTERS_reg[19][10]  ( .G(n281), .D(n413), .Q(\REGISTERS[19][10] )
         );
  DLH_X1 \REGISTERS_reg[19][9]  ( .G(n280), .D(n417), .Q(\REGISTERS[19][9] )
         );
  DLH_X1 \REGISTERS_reg[19][8]  ( .G(n280), .D(n421), .Q(\REGISTERS[19][8] )
         );
  DLH_X1 \REGISTERS_reg[19][7]  ( .G(n280), .D(n425), .Q(\REGISTERS[19][7] )
         );
  DLH_X1 \REGISTERS_reg[19][6]  ( .G(n280), .D(n429), .Q(\REGISTERS[19][6] )
         );
  DLH_X1 \REGISTERS_reg[19][5]  ( .G(n280), .D(n433), .Q(\REGISTERS[19][5] )
         );
  DLH_X1 \REGISTERS_reg[19][4]  ( .G(n280), .D(n437), .Q(\REGISTERS[19][4] )
         );
  DLH_X1 \REGISTERS_reg[19][3]  ( .G(n280), .D(n441), .Q(\REGISTERS[19][3] )
         );
  DLH_X1 \REGISTERS_reg[19][2]  ( .G(n280), .D(n445), .Q(\REGISTERS[19][2] )
         );
  DLH_X1 \REGISTERS_reg[19][1]  ( .G(n280), .D(n449), .Q(\REGISTERS[19][1] )
         );
  DLH_X1 \REGISTERS_reg[19][0]  ( .G(n280), .D(n453), .Q(\REGISTERS[19][0] )
         );
  DLH_X1 \REGISTERS_reg[20][31]  ( .G(n287), .D(n330), .Q(\REGISTERS[20][31] )
         );
  DLH_X1 \REGISTERS_reg[20][30]  ( .G(n287), .D(n334), .Q(\REGISTERS[20][30] )
         );
  DLH_X1 \REGISTERS_reg[20][29]  ( .G(n286), .D(n338), .Q(\REGISTERS[20][29] )
         );
  DLH_X1 \REGISTERS_reg[20][28]  ( .G(n286), .D(n342), .Q(\REGISTERS[20][28] )
         );
  DLH_X1 \REGISTERS_reg[20][27]  ( .G(n286), .D(n346), .Q(\REGISTERS[20][27] )
         );
  DLH_X1 \REGISTERS_reg[20][26]  ( .G(n286), .D(n350), .Q(\REGISTERS[20][26] )
         );
  DLH_X1 \REGISTERS_reg[20][25]  ( .G(n286), .D(n354), .Q(\REGISTERS[20][25] )
         );
  DLH_X1 \REGISTERS_reg[20][24]  ( .G(n286), .D(n358), .Q(\REGISTERS[20][24] )
         );
  DLH_X1 \REGISTERS_reg[20][23]  ( .G(n286), .D(n362), .Q(\REGISTERS[20][23] )
         );
  DLH_X1 \REGISTERS_reg[20][22]  ( .G(n286), .D(n366), .Q(\REGISTERS[20][22] )
         );
  DLH_X1 \REGISTERS_reg[20][21]  ( .G(n286), .D(n370), .Q(\REGISTERS[20][21] )
         );
  DLH_X1 \REGISTERS_reg[20][20]  ( .G(n286), .D(n374), .Q(\REGISTERS[20][20] )
         );
  DLH_X1 \REGISTERS_reg[20][19]  ( .G(n285), .D(n378), .Q(\REGISTERS[20][19] )
         );
  DLH_X1 \REGISTERS_reg[20][18]  ( .G(n285), .D(n382), .Q(\REGISTERS[20][18] )
         );
  DLH_X1 \REGISTERS_reg[20][17]  ( .G(n285), .D(n386), .Q(\REGISTERS[20][17] )
         );
  DLH_X1 \REGISTERS_reg[20][16]  ( .G(n285), .D(n390), .Q(\REGISTERS[20][16] )
         );
  DLH_X1 \REGISTERS_reg[20][15]  ( .G(n285), .D(n394), .Q(\REGISTERS[20][15] )
         );
  DLH_X1 \REGISTERS_reg[20][14]  ( .G(n285), .D(n398), .Q(\REGISTERS[20][14] )
         );
  DLH_X1 \REGISTERS_reg[20][13]  ( .G(n285), .D(n402), .Q(\REGISTERS[20][13] )
         );
  DLH_X1 \REGISTERS_reg[20][12]  ( .G(n285), .D(n406), .Q(\REGISTERS[20][12] )
         );
  DLH_X1 \REGISTERS_reg[20][11]  ( .G(n285), .D(n410), .Q(\REGISTERS[20][11] )
         );
  DLH_X1 \REGISTERS_reg[20][10]  ( .G(n285), .D(n414), .Q(\REGISTERS[20][10] )
         );
  DLH_X1 \REGISTERS_reg[20][9]  ( .G(n284), .D(n418), .Q(\REGISTERS[20][9] )
         );
  DLH_X1 \REGISTERS_reg[20][8]  ( .G(n284), .D(n422), .Q(\REGISTERS[20][8] )
         );
  DLH_X1 \REGISTERS_reg[20][7]  ( .G(n284), .D(n426), .Q(\REGISTERS[20][7] )
         );
  DLH_X1 \REGISTERS_reg[20][6]  ( .G(n284), .D(n430), .Q(\REGISTERS[20][6] )
         );
  DLH_X1 \REGISTERS_reg[20][5]  ( .G(n284), .D(n434), .Q(\REGISTERS[20][5] )
         );
  DLH_X1 \REGISTERS_reg[20][4]  ( .G(n284), .D(n438), .Q(\REGISTERS[20][4] )
         );
  DLH_X1 \REGISTERS_reg[20][3]  ( .G(n284), .D(n442), .Q(\REGISTERS[20][3] )
         );
  DLH_X1 \REGISTERS_reg[20][2]  ( .G(n284), .D(n446), .Q(\REGISTERS[20][2] )
         );
  DLH_X1 \REGISTERS_reg[20][1]  ( .G(n284), .D(n450), .Q(\REGISTERS[20][1] )
         );
  DLH_X1 \REGISTERS_reg[20][0]  ( .G(n284), .D(n454), .Q(\REGISTERS[20][0] )
         );
  DLH_X1 \REGISTERS_reg[21][31]  ( .G(n291), .D(n330), .Q(\REGISTERS[21][31] )
         );
  DLH_X1 \REGISTERS_reg[21][30]  ( .G(n291), .D(n334), .Q(\REGISTERS[21][30] )
         );
  DLH_X1 \REGISTERS_reg[21][29]  ( .G(n290), .D(n338), .Q(\REGISTERS[21][29] )
         );
  DLH_X1 \REGISTERS_reg[21][28]  ( .G(n290), .D(n342), .Q(\REGISTERS[21][28] )
         );
  DLH_X1 \REGISTERS_reg[21][27]  ( .G(n290), .D(n346), .Q(\REGISTERS[21][27] )
         );
  DLH_X1 \REGISTERS_reg[21][26]  ( .G(n290), .D(n350), .Q(\REGISTERS[21][26] )
         );
  DLH_X1 \REGISTERS_reg[21][25]  ( .G(n290), .D(n354), .Q(\REGISTERS[21][25] )
         );
  DLH_X1 \REGISTERS_reg[21][24]  ( .G(n290), .D(n358), .Q(\REGISTERS[21][24] )
         );
  DLH_X1 \REGISTERS_reg[21][23]  ( .G(n290), .D(n362), .Q(\REGISTERS[21][23] )
         );
  DLH_X1 \REGISTERS_reg[21][22]  ( .G(n290), .D(n366), .Q(\REGISTERS[21][22] )
         );
  DLH_X1 \REGISTERS_reg[21][21]  ( .G(n290), .D(n370), .Q(\REGISTERS[21][21] )
         );
  DLH_X1 \REGISTERS_reg[21][20]  ( .G(n290), .D(n374), .Q(\REGISTERS[21][20] )
         );
  DLH_X1 \REGISTERS_reg[21][19]  ( .G(n289), .D(n378), .Q(\REGISTERS[21][19] )
         );
  DLH_X1 \REGISTERS_reg[21][18]  ( .G(n289), .D(n382), .Q(\REGISTERS[21][18] )
         );
  DLH_X1 \REGISTERS_reg[21][17]  ( .G(n289), .D(n386), .Q(\REGISTERS[21][17] )
         );
  DLH_X1 \REGISTERS_reg[21][16]  ( .G(n289), .D(n390), .Q(\REGISTERS[21][16] )
         );
  DLH_X1 \REGISTERS_reg[21][15]  ( .G(n289), .D(n394), .Q(\REGISTERS[21][15] )
         );
  DLH_X1 \REGISTERS_reg[21][14]  ( .G(n289), .D(n398), .Q(\REGISTERS[21][14] )
         );
  DLH_X1 \REGISTERS_reg[21][13]  ( .G(n289), .D(n402), .Q(\REGISTERS[21][13] )
         );
  DLH_X1 \REGISTERS_reg[21][12]  ( .G(n289), .D(n406), .Q(\REGISTERS[21][12] )
         );
  DLH_X1 \REGISTERS_reg[21][11]  ( .G(n289), .D(n410), .Q(\REGISTERS[21][11] )
         );
  DLH_X1 \REGISTERS_reg[21][10]  ( .G(n289), .D(n414), .Q(\REGISTERS[21][10] )
         );
  DLH_X1 \REGISTERS_reg[21][9]  ( .G(n288), .D(n418), .Q(\REGISTERS[21][9] )
         );
  DLH_X1 \REGISTERS_reg[21][8]  ( .G(n288), .D(n422), .Q(\REGISTERS[21][8] )
         );
  DLH_X1 \REGISTERS_reg[21][7]  ( .G(n288), .D(n426), .Q(\REGISTERS[21][7] )
         );
  DLH_X1 \REGISTERS_reg[21][6]  ( .G(n288), .D(n430), .Q(\REGISTERS[21][6] )
         );
  DLH_X1 \REGISTERS_reg[21][5]  ( .G(n288), .D(n434), .Q(\REGISTERS[21][5] )
         );
  DLH_X1 \REGISTERS_reg[21][4]  ( .G(n288), .D(n438), .Q(\REGISTERS[21][4] )
         );
  DLH_X1 \REGISTERS_reg[21][3]  ( .G(n288), .D(n442), .Q(\REGISTERS[21][3] )
         );
  DLH_X1 \REGISTERS_reg[21][2]  ( .G(n288), .D(n446), .Q(\REGISTERS[21][2] )
         );
  DLH_X1 \REGISTERS_reg[21][1]  ( .G(n288), .D(n450), .Q(\REGISTERS[21][1] )
         );
  DLH_X1 \REGISTERS_reg[21][0]  ( .G(n288), .D(n454), .Q(\REGISTERS[21][0] )
         );
  DLH_X1 \REGISTERS_reg[22][31]  ( .G(n295), .D(n330), .Q(\REGISTERS[22][31] )
         );
  DLH_X1 \REGISTERS_reg[22][30]  ( .G(n295), .D(n334), .Q(\REGISTERS[22][30] )
         );
  DLH_X1 \REGISTERS_reg[22][29]  ( .G(n294), .D(n338), .Q(\REGISTERS[22][29] )
         );
  DLH_X1 \REGISTERS_reg[22][28]  ( .G(n294), .D(n342), .Q(\REGISTERS[22][28] )
         );
  DLH_X1 \REGISTERS_reg[22][27]  ( .G(n294), .D(n346), .Q(\REGISTERS[22][27] )
         );
  DLH_X1 \REGISTERS_reg[22][26]  ( .G(n294), .D(n350), .Q(\REGISTERS[22][26] )
         );
  DLH_X1 \REGISTERS_reg[22][25]  ( .G(n294), .D(n354), .Q(\REGISTERS[22][25] )
         );
  DLH_X1 \REGISTERS_reg[22][24]  ( .G(n294), .D(n358), .Q(\REGISTERS[22][24] )
         );
  DLH_X1 \REGISTERS_reg[22][23]  ( .G(n294), .D(n362), .Q(\REGISTERS[22][23] )
         );
  DLH_X1 \REGISTERS_reg[22][22]  ( .G(n294), .D(n366), .Q(\REGISTERS[22][22] )
         );
  DLH_X1 \REGISTERS_reg[22][21]  ( .G(n294), .D(n370), .Q(\REGISTERS[22][21] )
         );
  DLH_X1 \REGISTERS_reg[22][20]  ( .G(n294), .D(n374), .Q(\REGISTERS[22][20] )
         );
  DLH_X1 \REGISTERS_reg[22][19]  ( .G(n293), .D(n378), .Q(\REGISTERS[22][19] )
         );
  DLH_X1 \REGISTERS_reg[22][18]  ( .G(n293), .D(n382), .Q(\REGISTERS[22][18] )
         );
  DLH_X1 \REGISTERS_reg[22][17]  ( .G(n293), .D(n386), .Q(\REGISTERS[22][17] )
         );
  DLH_X1 \REGISTERS_reg[22][16]  ( .G(n293), .D(n390), .Q(\REGISTERS[22][16] )
         );
  DLH_X1 \REGISTERS_reg[22][15]  ( .G(n293), .D(n394), .Q(\REGISTERS[22][15] )
         );
  DLH_X1 \REGISTERS_reg[22][14]  ( .G(n293), .D(n398), .Q(\REGISTERS[22][14] )
         );
  DLH_X1 \REGISTERS_reg[22][13]  ( .G(n293), .D(n402), .Q(\REGISTERS[22][13] )
         );
  DLH_X1 \REGISTERS_reg[22][12]  ( .G(n293), .D(n406), .Q(\REGISTERS[22][12] )
         );
  DLH_X1 \REGISTERS_reg[22][11]  ( .G(n293), .D(n410), .Q(\REGISTERS[22][11] )
         );
  DLH_X1 \REGISTERS_reg[22][10]  ( .G(n293), .D(n414), .Q(\REGISTERS[22][10] )
         );
  DLH_X1 \REGISTERS_reg[22][9]  ( .G(n292), .D(n418), .Q(\REGISTERS[22][9] )
         );
  DLH_X1 \REGISTERS_reg[22][8]  ( .G(n292), .D(n422), .Q(\REGISTERS[22][8] )
         );
  DLH_X1 \REGISTERS_reg[22][7]  ( .G(n292), .D(n426), .Q(\REGISTERS[22][7] )
         );
  DLH_X1 \REGISTERS_reg[22][6]  ( .G(n292), .D(n430), .Q(\REGISTERS[22][6] )
         );
  DLH_X1 \REGISTERS_reg[22][5]  ( .G(n292), .D(n434), .Q(\REGISTERS[22][5] )
         );
  DLH_X1 \REGISTERS_reg[22][4]  ( .G(n292), .D(n438), .Q(\REGISTERS[22][4] )
         );
  DLH_X1 \REGISTERS_reg[22][3]  ( .G(n292), .D(n442), .Q(\REGISTERS[22][3] )
         );
  DLH_X1 \REGISTERS_reg[22][2]  ( .G(n292), .D(n446), .Q(\REGISTERS[22][2] )
         );
  DLH_X1 \REGISTERS_reg[22][1]  ( .G(n292), .D(n450), .Q(\REGISTERS[22][1] )
         );
  DLH_X1 \REGISTERS_reg[22][0]  ( .G(n292), .D(n454), .Q(\REGISTERS[22][0] )
         );
  DLH_X1 \REGISTERS_reg[23][31]  ( .G(n299), .D(n330), .Q(\REGISTERS[23][31] )
         );
  DLH_X1 \REGISTERS_reg[23][30]  ( .G(n299), .D(n334), .Q(\REGISTERS[23][30] )
         );
  DLH_X1 \REGISTERS_reg[23][29]  ( .G(n298), .D(n338), .Q(\REGISTERS[23][29] )
         );
  DLH_X1 \REGISTERS_reg[23][28]  ( .G(n298), .D(n342), .Q(\REGISTERS[23][28] )
         );
  DLH_X1 \REGISTERS_reg[23][27]  ( .G(n298), .D(n346), .Q(\REGISTERS[23][27] )
         );
  DLH_X1 \REGISTERS_reg[23][26]  ( .G(n298), .D(n350), .Q(\REGISTERS[23][26] )
         );
  DLH_X1 \REGISTERS_reg[23][25]  ( .G(n298), .D(n354), .Q(\REGISTERS[23][25] )
         );
  DLH_X1 \REGISTERS_reg[23][24]  ( .G(n298), .D(n358), .Q(\REGISTERS[23][24] )
         );
  DLH_X1 \REGISTERS_reg[23][23]  ( .G(n298), .D(n362), .Q(\REGISTERS[23][23] )
         );
  DLH_X1 \REGISTERS_reg[23][22]  ( .G(n298), .D(n366), .Q(\REGISTERS[23][22] )
         );
  DLH_X1 \REGISTERS_reg[23][21]  ( .G(n298), .D(n370), .Q(\REGISTERS[23][21] )
         );
  DLH_X1 \REGISTERS_reg[23][20]  ( .G(n298), .D(n374), .Q(\REGISTERS[23][20] )
         );
  DLH_X1 \REGISTERS_reg[23][19]  ( .G(n297), .D(n378), .Q(\REGISTERS[23][19] )
         );
  DLH_X1 \REGISTERS_reg[23][18]  ( .G(n297), .D(n382), .Q(\REGISTERS[23][18] )
         );
  DLH_X1 \REGISTERS_reg[23][17]  ( .G(n297), .D(n386), .Q(\REGISTERS[23][17] )
         );
  DLH_X1 \REGISTERS_reg[23][16]  ( .G(n297), .D(n390), .Q(\REGISTERS[23][16] )
         );
  DLH_X1 \REGISTERS_reg[23][15]  ( .G(n297), .D(n394), .Q(\REGISTERS[23][15] )
         );
  DLH_X1 \REGISTERS_reg[23][14]  ( .G(n297), .D(n398), .Q(\REGISTERS[23][14] )
         );
  DLH_X1 \REGISTERS_reg[23][13]  ( .G(n297), .D(n402), .Q(\REGISTERS[23][13] )
         );
  DLH_X1 \REGISTERS_reg[23][12]  ( .G(n297), .D(n406), .Q(\REGISTERS[23][12] )
         );
  DLH_X1 \REGISTERS_reg[23][11]  ( .G(n297), .D(n410), .Q(\REGISTERS[23][11] )
         );
  DLH_X1 \REGISTERS_reg[23][10]  ( .G(n297), .D(n414), .Q(\REGISTERS[23][10] )
         );
  DLH_X1 \REGISTERS_reg[23][9]  ( .G(n296), .D(n418), .Q(\REGISTERS[23][9] )
         );
  DLH_X1 \REGISTERS_reg[23][8]  ( .G(n296), .D(n422), .Q(\REGISTERS[23][8] )
         );
  DLH_X1 \REGISTERS_reg[23][7]  ( .G(n296), .D(n426), .Q(\REGISTERS[23][7] )
         );
  DLH_X1 \REGISTERS_reg[23][6]  ( .G(n296), .D(n430), .Q(\REGISTERS[23][6] )
         );
  DLH_X1 \REGISTERS_reg[23][5]  ( .G(n296), .D(n434), .Q(\REGISTERS[23][5] )
         );
  DLH_X1 \REGISTERS_reg[23][4]  ( .G(n296), .D(n438), .Q(\REGISTERS[23][4] )
         );
  DLH_X1 \REGISTERS_reg[23][3]  ( .G(n296), .D(n442), .Q(\REGISTERS[23][3] )
         );
  DLH_X1 \REGISTERS_reg[23][2]  ( .G(n296), .D(n446), .Q(\REGISTERS[23][2] )
         );
  DLH_X1 \REGISTERS_reg[23][1]  ( .G(n296), .D(n450), .Q(\REGISTERS[23][1] )
         );
  DLH_X1 \REGISTERS_reg[23][0]  ( .G(n296), .D(n454), .Q(\REGISTERS[23][0] )
         );
  DLH_X1 \REGISTERS_reg[24][31]  ( .G(n303), .D(n330), .Q(\REGISTERS[24][31] )
         );
  DLH_X1 \REGISTERS_reg[24][30]  ( .G(n303), .D(n334), .Q(\REGISTERS[24][30] )
         );
  DLH_X1 \REGISTERS_reg[24][29]  ( .G(n302), .D(n338), .Q(\REGISTERS[24][29] )
         );
  DLH_X1 \REGISTERS_reg[24][28]  ( .G(n302), .D(n342), .Q(\REGISTERS[24][28] )
         );
  DLH_X1 \REGISTERS_reg[24][27]  ( .G(n302), .D(n346), .Q(\REGISTERS[24][27] )
         );
  DLH_X1 \REGISTERS_reg[24][26]  ( .G(n302), .D(n350), .Q(\REGISTERS[24][26] )
         );
  DLH_X1 \REGISTERS_reg[24][25]  ( .G(n302), .D(n354), .Q(\REGISTERS[24][25] )
         );
  DLH_X1 \REGISTERS_reg[24][24]  ( .G(n302), .D(n358), .Q(\REGISTERS[24][24] )
         );
  DLH_X1 \REGISTERS_reg[24][23]  ( .G(n302), .D(n362), .Q(\REGISTERS[24][23] )
         );
  DLH_X1 \REGISTERS_reg[24][22]  ( .G(n302), .D(n366), .Q(\REGISTERS[24][22] )
         );
  DLH_X1 \REGISTERS_reg[24][21]  ( .G(n302), .D(n370), .Q(\REGISTERS[24][21] )
         );
  DLH_X1 \REGISTERS_reg[24][20]  ( .G(n302), .D(n374), .Q(\REGISTERS[24][20] )
         );
  DLH_X1 \REGISTERS_reg[24][19]  ( .G(n301), .D(n378), .Q(\REGISTERS[24][19] )
         );
  DLH_X1 \REGISTERS_reg[24][18]  ( .G(n301), .D(n382), .Q(\REGISTERS[24][18] )
         );
  DLH_X1 \REGISTERS_reg[24][17]  ( .G(n301), .D(n386), .Q(\REGISTERS[24][17] )
         );
  DLH_X1 \REGISTERS_reg[24][16]  ( .G(n301), .D(n390), .Q(\REGISTERS[24][16] )
         );
  DLH_X1 \REGISTERS_reg[24][15]  ( .G(n301), .D(n394), .Q(\REGISTERS[24][15] )
         );
  DLH_X1 \REGISTERS_reg[24][14]  ( .G(n301), .D(n398), .Q(\REGISTERS[24][14] )
         );
  DLH_X1 \REGISTERS_reg[24][13]  ( .G(n301), .D(n402), .Q(\REGISTERS[24][13] )
         );
  DLH_X1 \REGISTERS_reg[24][12]  ( .G(n301), .D(n406), .Q(\REGISTERS[24][12] )
         );
  DLH_X1 \REGISTERS_reg[24][11]  ( .G(n301), .D(n410), .Q(\REGISTERS[24][11] )
         );
  DLH_X1 \REGISTERS_reg[24][10]  ( .G(n301), .D(n414), .Q(\REGISTERS[24][10] )
         );
  DLH_X1 \REGISTERS_reg[24][9]  ( .G(n300), .D(n418), .Q(\REGISTERS[24][9] )
         );
  DLH_X1 \REGISTERS_reg[24][8]  ( .G(n300), .D(n422), .Q(\REGISTERS[24][8] )
         );
  DLH_X1 \REGISTERS_reg[24][7]  ( .G(n300), .D(n426), .Q(\REGISTERS[24][7] )
         );
  DLH_X1 \REGISTERS_reg[24][6]  ( .G(n300), .D(n430), .Q(\REGISTERS[24][6] )
         );
  DLH_X1 \REGISTERS_reg[24][5]  ( .G(n300), .D(n434), .Q(\REGISTERS[24][5] )
         );
  DLH_X1 \REGISTERS_reg[24][4]  ( .G(n300), .D(n438), .Q(\REGISTERS[24][4] )
         );
  DLH_X1 \REGISTERS_reg[24][3]  ( .G(n300), .D(n442), .Q(\REGISTERS[24][3] )
         );
  DLH_X1 \REGISTERS_reg[24][2]  ( .G(n300), .D(n446), .Q(\REGISTERS[24][2] )
         );
  DLH_X1 \REGISTERS_reg[24][1]  ( .G(n300), .D(n450), .Q(\REGISTERS[24][1] )
         );
  DLH_X1 \REGISTERS_reg[24][0]  ( .G(n300), .D(n454), .Q(\REGISTERS[24][0] )
         );
  DLH_X1 \REGISTERS_reg[25][31]  ( .G(n307), .D(n330), .Q(\REGISTERS[25][31] )
         );
  DLH_X1 \REGISTERS_reg[25][30]  ( .G(n307), .D(n334), .Q(\REGISTERS[25][30] )
         );
  DLH_X1 \REGISTERS_reg[25][29]  ( .G(n306), .D(n338), .Q(\REGISTERS[25][29] )
         );
  DLH_X1 \REGISTERS_reg[25][28]  ( .G(n306), .D(n342), .Q(\REGISTERS[25][28] )
         );
  DLH_X1 \REGISTERS_reg[25][27]  ( .G(n306), .D(n346), .Q(\REGISTERS[25][27] )
         );
  DLH_X1 \REGISTERS_reg[25][26]  ( .G(n306), .D(n350), .Q(\REGISTERS[25][26] )
         );
  DLH_X1 \REGISTERS_reg[25][25]  ( .G(n306), .D(n354), .Q(\REGISTERS[25][25] )
         );
  DLH_X1 \REGISTERS_reg[25][24]  ( .G(n306), .D(n358), .Q(\REGISTERS[25][24] )
         );
  DLH_X1 \REGISTERS_reg[25][23]  ( .G(n306), .D(n362), .Q(\REGISTERS[25][23] )
         );
  DLH_X1 \REGISTERS_reg[25][22]  ( .G(n306), .D(n366), .Q(\REGISTERS[25][22] )
         );
  DLH_X1 \REGISTERS_reg[25][21]  ( .G(n306), .D(n370), .Q(\REGISTERS[25][21] )
         );
  DLH_X1 \REGISTERS_reg[25][20]  ( .G(n306), .D(n374), .Q(\REGISTERS[25][20] )
         );
  DLH_X1 \REGISTERS_reg[25][19]  ( .G(n305), .D(n378), .Q(\REGISTERS[25][19] )
         );
  DLH_X1 \REGISTERS_reg[25][18]  ( .G(n305), .D(n382), .Q(\REGISTERS[25][18] )
         );
  DLH_X1 \REGISTERS_reg[25][17]  ( .G(n305), .D(n386), .Q(\REGISTERS[25][17] )
         );
  DLH_X1 \REGISTERS_reg[25][16]  ( .G(n305), .D(n390), .Q(\REGISTERS[25][16] )
         );
  DLH_X1 \REGISTERS_reg[25][15]  ( .G(n305), .D(n394), .Q(\REGISTERS[25][15] )
         );
  DLH_X1 \REGISTERS_reg[25][14]  ( .G(n305), .D(n398), .Q(\REGISTERS[25][14] )
         );
  DLH_X1 \REGISTERS_reg[25][13]  ( .G(n305), .D(n402), .Q(\REGISTERS[25][13] )
         );
  DLH_X1 \REGISTERS_reg[25][12]  ( .G(n305), .D(n406), .Q(\REGISTERS[25][12] )
         );
  DLH_X1 \REGISTERS_reg[25][11]  ( .G(n305), .D(n410), .Q(\REGISTERS[25][11] )
         );
  DLH_X1 \REGISTERS_reg[25][10]  ( .G(n305), .D(n414), .Q(\REGISTERS[25][10] )
         );
  DLH_X1 \REGISTERS_reg[25][9]  ( .G(n304), .D(n418), .Q(\REGISTERS[25][9] )
         );
  DLH_X1 \REGISTERS_reg[25][8]  ( .G(n304), .D(n422), .Q(\REGISTERS[25][8] )
         );
  DLH_X1 \REGISTERS_reg[25][7]  ( .G(n304), .D(n426), .Q(\REGISTERS[25][7] )
         );
  DLH_X1 \REGISTERS_reg[25][6]  ( .G(n304), .D(n430), .Q(\REGISTERS[25][6] )
         );
  DLH_X1 \REGISTERS_reg[25][5]  ( .G(n304), .D(n434), .Q(\REGISTERS[25][5] )
         );
  DLH_X1 \REGISTERS_reg[25][4]  ( .G(n304), .D(n438), .Q(\REGISTERS[25][4] )
         );
  DLH_X1 \REGISTERS_reg[25][3]  ( .G(n304), .D(n442), .Q(\REGISTERS[25][3] )
         );
  DLH_X1 \REGISTERS_reg[25][2]  ( .G(n304), .D(n446), .Q(\REGISTERS[25][2] )
         );
  DLH_X1 \REGISTERS_reg[25][1]  ( .G(n304), .D(n450), .Q(\REGISTERS[25][1] )
         );
  DLH_X1 \REGISTERS_reg[25][0]  ( .G(n304), .D(n454), .Q(\REGISTERS[25][0] )
         );
  DLH_X1 \REGISTERS_reg[26][31]  ( .G(n311), .D(n330), .Q(\REGISTERS[26][31] )
         );
  DLH_X1 \REGISTERS_reg[26][30]  ( .G(n311), .D(n334), .Q(\REGISTERS[26][30] )
         );
  DLH_X1 \REGISTERS_reg[26][29]  ( .G(n310), .D(n338), .Q(\REGISTERS[26][29] )
         );
  DLH_X1 \REGISTERS_reg[26][28]  ( .G(n310), .D(n342), .Q(\REGISTERS[26][28] )
         );
  DLH_X1 \REGISTERS_reg[26][27]  ( .G(n310), .D(n346), .Q(\REGISTERS[26][27] )
         );
  DLH_X1 \REGISTERS_reg[26][26]  ( .G(n310), .D(n350), .Q(\REGISTERS[26][26] )
         );
  DLH_X1 \REGISTERS_reg[26][25]  ( .G(n310), .D(n354), .Q(\REGISTERS[26][25] )
         );
  DLH_X1 \REGISTERS_reg[26][24]  ( .G(n310), .D(n358), .Q(\REGISTERS[26][24] )
         );
  DLH_X1 \REGISTERS_reg[26][23]  ( .G(n310), .D(n362), .Q(\REGISTERS[26][23] )
         );
  DLH_X1 \REGISTERS_reg[26][22]  ( .G(n310), .D(n366), .Q(\REGISTERS[26][22] )
         );
  DLH_X1 \REGISTERS_reg[26][21]  ( .G(n310), .D(n370), .Q(\REGISTERS[26][21] )
         );
  DLH_X1 \REGISTERS_reg[26][20]  ( .G(n310), .D(n374), .Q(\REGISTERS[26][20] )
         );
  DLH_X1 \REGISTERS_reg[26][19]  ( .G(n309), .D(n378), .Q(\REGISTERS[26][19] )
         );
  DLH_X1 \REGISTERS_reg[26][18]  ( .G(n309), .D(n382), .Q(\REGISTERS[26][18] )
         );
  DLH_X1 \REGISTERS_reg[26][17]  ( .G(n309), .D(n386), .Q(\REGISTERS[26][17] )
         );
  DLH_X1 \REGISTERS_reg[26][16]  ( .G(n309), .D(n390), .Q(\REGISTERS[26][16] )
         );
  DLH_X1 \REGISTERS_reg[26][15]  ( .G(n309), .D(n394), .Q(\REGISTERS[26][15] )
         );
  DLH_X1 \REGISTERS_reg[26][14]  ( .G(n309), .D(n398), .Q(\REGISTERS[26][14] )
         );
  DLH_X1 \REGISTERS_reg[26][13]  ( .G(n309), .D(n402), .Q(\REGISTERS[26][13] )
         );
  DLH_X1 \REGISTERS_reg[26][12]  ( .G(n309), .D(n406), .Q(\REGISTERS[26][12] )
         );
  DLH_X1 \REGISTERS_reg[26][11]  ( .G(n309), .D(n410), .Q(\REGISTERS[26][11] )
         );
  DLH_X1 \REGISTERS_reg[26][10]  ( .G(n309), .D(n414), .Q(\REGISTERS[26][10] )
         );
  DLH_X1 \REGISTERS_reg[26][9]  ( .G(n308), .D(n418), .Q(\REGISTERS[26][9] )
         );
  DLH_X1 \REGISTERS_reg[26][8]  ( .G(n308), .D(n422), .Q(\REGISTERS[26][8] )
         );
  DLH_X1 \REGISTERS_reg[26][7]  ( .G(n308), .D(n426), .Q(\REGISTERS[26][7] )
         );
  DLH_X1 \REGISTERS_reg[26][6]  ( .G(n308), .D(n430), .Q(\REGISTERS[26][6] )
         );
  DLH_X1 \REGISTERS_reg[26][5]  ( .G(n308), .D(n434), .Q(\REGISTERS[26][5] )
         );
  DLH_X1 \REGISTERS_reg[26][4]  ( .G(n308), .D(n438), .Q(\REGISTERS[26][4] )
         );
  DLH_X1 \REGISTERS_reg[26][3]  ( .G(n308), .D(n442), .Q(\REGISTERS[26][3] )
         );
  DLH_X1 \REGISTERS_reg[26][2]  ( .G(n308), .D(n446), .Q(\REGISTERS[26][2] )
         );
  DLH_X1 \REGISTERS_reg[26][1]  ( .G(n308), .D(n450), .Q(\REGISTERS[26][1] )
         );
  DLH_X1 \REGISTERS_reg[26][0]  ( .G(n308), .D(n454), .Q(\REGISTERS[26][0] )
         );
  DLH_X1 \REGISTERS_reg[27][31]  ( .G(n315), .D(n330), .Q(\REGISTERS[27][31] )
         );
  DLH_X1 \REGISTERS_reg[27][30]  ( .G(n315), .D(n334), .Q(\REGISTERS[27][30] )
         );
  DLH_X1 \REGISTERS_reg[27][29]  ( .G(n314), .D(n338), .Q(\REGISTERS[27][29] )
         );
  DLH_X1 \REGISTERS_reg[27][28]  ( .G(n314), .D(n342), .Q(\REGISTERS[27][28] )
         );
  DLH_X1 \REGISTERS_reg[27][27]  ( .G(n314), .D(n346), .Q(\REGISTERS[27][27] )
         );
  DLH_X1 \REGISTERS_reg[27][26]  ( .G(n314), .D(n350), .Q(\REGISTERS[27][26] )
         );
  DLH_X1 \REGISTERS_reg[27][25]  ( .G(n314), .D(n354), .Q(\REGISTERS[27][25] )
         );
  DLH_X1 \REGISTERS_reg[27][24]  ( .G(n314), .D(n358), .Q(\REGISTERS[27][24] )
         );
  DLH_X1 \REGISTERS_reg[27][23]  ( .G(n314), .D(n362), .Q(\REGISTERS[27][23] )
         );
  DLH_X1 \REGISTERS_reg[27][22]  ( .G(n314), .D(n366), .Q(\REGISTERS[27][22] )
         );
  DLH_X1 \REGISTERS_reg[27][21]  ( .G(n314), .D(n370), .Q(\REGISTERS[27][21] )
         );
  DLH_X1 \REGISTERS_reg[27][20]  ( .G(n314), .D(n374), .Q(\REGISTERS[27][20] )
         );
  DLH_X1 \REGISTERS_reg[27][19]  ( .G(n313), .D(n378), .Q(\REGISTERS[27][19] )
         );
  DLH_X1 \REGISTERS_reg[27][18]  ( .G(n313), .D(n382), .Q(\REGISTERS[27][18] )
         );
  DLH_X1 \REGISTERS_reg[27][17]  ( .G(n313), .D(n386), .Q(\REGISTERS[27][17] )
         );
  DLH_X1 \REGISTERS_reg[27][16]  ( .G(n313), .D(n390), .Q(\REGISTERS[27][16] )
         );
  DLH_X1 \REGISTERS_reg[27][15]  ( .G(n313), .D(n394), .Q(\REGISTERS[27][15] )
         );
  DLH_X1 \REGISTERS_reg[27][14]  ( .G(n313), .D(n398), .Q(\REGISTERS[27][14] )
         );
  DLH_X1 \REGISTERS_reg[27][13]  ( .G(n313), .D(n402), .Q(\REGISTERS[27][13] )
         );
  DLH_X1 \REGISTERS_reg[27][12]  ( .G(n313), .D(n406), .Q(\REGISTERS[27][12] )
         );
  DLH_X1 \REGISTERS_reg[27][11]  ( .G(n313), .D(n410), .Q(\REGISTERS[27][11] )
         );
  DLH_X1 \REGISTERS_reg[27][10]  ( .G(n313), .D(n414), .Q(\REGISTERS[27][10] )
         );
  DLH_X1 \REGISTERS_reg[27][9]  ( .G(n312), .D(n418), .Q(\REGISTERS[27][9] )
         );
  DLH_X1 \REGISTERS_reg[27][8]  ( .G(n312), .D(n422), .Q(\REGISTERS[27][8] )
         );
  DLH_X1 \REGISTERS_reg[27][7]  ( .G(n312), .D(n426), .Q(\REGISTERS[27][7] )
         );
  DLH_X1 \REGISTERS_reg[27][6]  ( .G(n312), .D(n430), .Q(\REGISTERS[27][6] )
         );
  DLH_X1 \REGISTERS_reg[27][5]  ( .G(n312), .D(n434), .Q(\REGISTERS[27][5] )
         );
  DLH_X1 \REGISTERS_reg[27][4]  ( .G(n312), .D(n438), .Q(\REGISTERS[27][4] )
         );
  DLH_X1 \REGISTERS_reg[27][3]  ( .G(n312), .D(n442), .Q(\REGISTERS[27][3] )
         );
  DLH_X1 \REGISTERS_reg[27][2]  ( .G(n312), .D(n446), .Q(\REGISTERS[27][2] )
         );
  DLH_X1 \REGISTERS_reg[27][1]  ( .G(n312), .D(n450), .Q(\REGISTERS[27][1] )
         );
  DLH_X1 \REGISTERS_reg[27][0]  ( .G(n312), .D(n454), .Q(\REGISTERS[27][0] )
         );
  DLH_X1 \REGISTERS_reg[28][31]  ( .G(n319), .D(n330), .Q(\REGISTERS[28][31] )
         );
  DLH_X1 \REGISTERS_reg[28][30]  ( .G(n319), .D(n334), .Q(\REGISTERS[28][30] )
         );
  DLH_X1 \REGISTERS_reg[28][29]  ( .G(n318), .D(n338), .Q(\REGISTERS[28][29] )
         );
  DLH_X1 \REGISTERS_reg[28][28]  ( .G(n318), .D(n342), .Q(\REGISTERS[28][28] )
         );
  DLH_X1 \REGISTERS_reg[28][27]  ( .G(n318), .D(n346), .Q(\REGISTERS[28][27] )
         );
  DLH_X1 \REGISTERS_reg[28][26]  ( .G(n318), .D(n350), .Q(\REGISTERS[28][26] )
         );
  DLH_X1 \REGISTERS_reg[28][25]  ( .G(n318), .D(n354), .Q(\REGISTERS[28][25] )
         );
  DLH_X1 \REGISTERS_reg[28][24]  ( .G(n318), .D(n358), .Q(\REGISTERS[28][24] )
         );
  DLH_X1 \REGISTERS_reg[28][23]  ( .G(n318), .D(n362), .Q(\REGISTERS[28][23] )
         );
  DLH_X1 \REGISTERS_reg[28][22]  ( .G(n318), .D(n366), .Q(\REGISTERS[28][22] )
         );
  DLH_X1 \REGISTERS_reg[28][21]  ( .G(n318), .D(n370), .Q(\REGISTERS[28][21] )
         );
  DLH_X1 \REGISTERS_reg[28][20]  ( .G(n318), .D(n374), .Q(\REGISTERS[28][20] )
         );
  DLH_X1 \REGISTERS_reg[28][19]  ( .G(n317), .D(n378), .Q(\REGISTERS[28][19] )
         );
  DLH_X1 \REGISTERS_reg[28][18]  ( .G(n317), .D(n382), .Q(\REGISTERS[28][18] )
         );
  DLH_X1 \REGISTERS_reg[28][17]  ( .G(n317), .D(n386), .Q(\REGISTERS[28][17] )
         );
  DLH_X1 \REGISTERS_reg[28][16]  ( .G(n317), .D(n390), .Q(\REGISTERS[28][16] )
         );
  DLH_X1 \REGISTERS_reg[28][15]  ( .G(n317), .D(n394), .Q(\REGISTERS[28][15] )
         );
  DLH_X1 \REGISTERS_reg[28][14]  ( .G(n317), .D(n398), .Q(\REGISTERS[28][14] )
         );
  DLH_X1 \REGISTERS_reg[28][13]  ( .G(n317), .D(n402), .Q(\REGISTERS[28][13] )
         );
  DLH_X1 \REGISTERS_reg[28][12]  ( .G(n317), .D(n406), .Q(\REGISTERS[28][12] )
         );
  DLH_X1 \REGISTERS_reg[28][11]  ( .G(n317), .D(n410), .Q(\REGISTERS[28][11] )
         );
  DLH_X1 \REGISTERS_reg[28][10]  ( .G(n317), .D(n414), .Q(\REGISTERS[28][10] )
         );
  DLH_X1 \REGISTERS_reg[28][9]  ( .G(n316), .D(n418), .Q(\REGISTERS[28][9] )
         );
  DLH_X1 \REGISTERS_reg[28][8]  ( .G(n316), .D(n422), .Q(\REGISTERS[28][8] )
         );
  DLH_X1 \REGISTERS_reg[28][7]  ( .G(n316), .D(n426), .Q(\REGISTERS[28][7] )
         );
  DLH_X1 \REGISTERS_reg[28][6]  ( .G(n316), .D(n430), .Q(\REGISTERS[28][6] )
         );
  DLH_X1 \REGISTERS_reg[28][5]  ( .G(n316), .D(n434), .Q(\REGISTERS[28][5] )
         );
  DLH_X1 \REGISTERS_reg[28][4]  ( .G(n316), .D(n438), .Q(\REGISTERS[28][4] )
         );
  DLH_X1 \REGISTERS_reg[28][3]  ( .G(n316), .D(n442), .Q(\REGISTERS[28][3] )
         );
  DLH_X1 \REGISTERS_reg[28][2]  ( .G(n316), .D(n446), .Q(\REGISTERS[28][2] )
         );
  DLH_X1 \REGISTERS_reg[28][1]  ( .G(n316), .D(n450), .Q(\REGISTERS[28][1] )
         );
  DLH_X1 \REGISTERS_reg[28][0]  ( .G(n316), .D(n454), .Q(\REGISTERS[28][0] )
         );
  DLH_X1 \REGISTERS_reg[29][31]  ( .G(n323), .D(n330), .Q(\REGISTERS[29][31] )
         );
  DLH_X1 \REGISTERS_reg[29][30]  ( .G(n323), .D(n334), .Q(\REGISTERS[29][30] )
         );
  DLH_X1 \REGISTERS_reg[29][29]  ( .G(n322), .D(n338), .Q(\REGISTERS[29][29] )
         );
  DLH_X1 \REGISTERS_reg[29][28]  ( .G(n322), .D(n342), .Q(\REGISTERS[29][28] )
         );
  DLH_X1 \REGISTERS_reg[29][27]  ( .G(n322), .D(n346), .Q(\REGISTERS[29][27] )
         );
  DLH_X1 \REGISTERS_reg[29][26]  ( .G(n322), .D(n350), .Q(\REGISTERS[29][26] )
         );
  DLH_X1 \REGISTERS_reg[29][25]  ( .G(n322), .D(n354), .Q(\REGISTERS[29][25] )
         );
  DLH_X1 \REGISTERS_reg[29][24]  ( .G(n322), .D(n358), .Q(\REGISTERS[29][24] )
         );
  DLH_X1 \REGISTERS_reg[29][23]  ( .G(n322), .D(n362), .Q(\REGISTERS[29][23] )
         );
  DLH_X1 \REGISTERS_reg[29][22]  ( .G(n322), .D(n366), .Q(\REGISTERS[29][22] )
         );
  DLH_X1 \REGISTERS_reg[29][21]  ( .G(n322), .D(n370), .Q(\REGISTERS[29][21] )
         );
  DLH_X1 \REGISTERS_reg[29][20]  ( .G(n322), .D(n374), .Q(\REGISTERS[29][20] )
         );
  DLH_X1 \REGISTERS_reg[29][19]  ( .G(n321), .D(n378), .Q(\REGISTERS[29][19] )
         );
  DLH_X1 \REGISTERS_reg[29][18]  ( .G(n321), .D(n382), .Q(\REGISTERS[29][18] )
         );
  DLH_X1 \REGISTERS_reg[29][17]  ( .G(n321), .D(n386), .Q(\REGISTERS[29][17] )
         );
  DLH_X1 \REGISTERS_reg[29][16]  ( .G(n321), .D(n390), .Q(\REGISTERS[29][16] )
         );
  DLH_X1 \REGISTERS_reg[29][15]  ( .G(n321), .D(n394), .Q(\REGISTERS[29][15] )
         );
  DLH_X1 \REGISTERS_reg[29][14]  ( .G(n321), .D(n398), .Q(\REGISTERS[29][14] )
         );
  DLH_X1 \REGISTERS_reg[29][13]  ( .G(n321), .D(n402), .Q(\REGISTERS[29][13] )
         );
  DLH_X1 \REGISTERS_reg[29][12]  ( .G(n321), .D(n406), .Q(\REGISTERS[29][12] )
         );
  DLH_X1 \REGISTERS_reg[29][11]  ( .G(n321), .D(n410), .Q(\REGISTERS[29][11] )
         );
  DLH_X1 \REGISTERS_reg[29][10]  ( .G(n321), .D(n414), .Q(\REGISTERS[29][10] )
         );
  DLH_X1 \REGISTERS_reg[29][9]  ( .G(n320), .D(n418), .Q(\REGISTERS[29][9] )
         );
  DLH_X1 \REGISTERS_reg[29][8]  ( .G(n320), .D(n422), .Q(\REGISTERS[29][8] )
         );
  DLH_X1 \REGISTERS_reg[29][7]  ( .G(n320), .D(n426), .Q(\REGISTERS[29][7] )
         );
  DLH_X1 \REGISTERS_reg[29][6]  ( .G(n320), .D(n430), .Q(\REGISTERS[29][6] )
         );
  DLH_X1 \REGISTERS_reg[29][5]  ( .G(n320), .D(n434), .Q(\REGISTERS[29][5] )
         );
  DLH_X1 \REGISTERS_reg[29][4]  ( .G(n320), .D(n438), .Q(\REGISTERS[29][4] )
         );
  DLH_X1 \REGISTERS_reg[29][3]  ( .G(n320), .D(n442), .Q(\REGISTERS[29][3] )
         );
  DLH_X1 \REGISTERS_reg[29][2]  ( .G(n320), .D(n446), .Q(\REGISTERS[29][2] )
         );
  DLH_X1 \REGISTERS_reg[29][1]  ( .G(n320), .D(n450), .Q(\REGISTERS[29][1] )
         );
  DLH_X1 \REGISTERS_reg[29][0]  ( .G(n320), .D(n454), .Q(\REGISTERS[29][0] )
         );
  DLH_X1 \REGISTERS_reg[30][31]  ( .G(n327), .D(n331), .Q(\REGISTERS[30][31] )
         );
  DLH_X1 \REGISTERS_reg[30][30]  ( .G(n327), .D(n335), .Q(\REGISTERS[30][30] )
         );
  DLH_X1 \REGISTERS_reg[30][29]  ( .G(n326), .D(n339), .Q(\REGISTERS[30][29] )
         );
  DLH_X1 \REGISTERS_reg[30][28]  ( .G(n326), .D(n343), .Q(\REGISTERS[30][28] )
         );
  DLH_X1 \REGISTERS_reg[30][27]  ( .G(n326), .D(n347), .Q(\REGISTERS[30][27] )
         );
  DLH_X1 \REGISTERS_reg[30][26]  ( .G(n326), .D(n351), .Q(\REGISTERS[30][26] )
         );
  DLH_X1 \REGISTERS_reg[30][25]  ( .G(n326), .D(n355), .Q(\REGISTERS[30][25] )
         );
  DLH_X1 \REGISTERS_reg[30][24]  ( .G(n326), .D(n359), .Q(\REGISTERS[30][24] )
         );
  DLH_X1 \REGISTERS_reg[30][23]  ( .G(n326), .D(n363), .Q(\REGISTERS[30][23] )
         );
  DLH_X1 \REGISTERS_reg[30][22]  ( .G(n326), .D(n367), .Q(\REGISTERS[30][22] )
         );
  DLH_X1 \REGISTERS_reg[30][21]  ( .G(n326), .D(n371), .Q(\REGISTERS[30][21] )
         );
  DLH_X1 \REGISTERS_reg[30][20]  ( .G(n326), .D(n375), .Q(\REGISTERS[30][20] )
         );
  DLH_X1 \REGISTERS_reg[30][19]  ( .G(n325), .D(n379), .Q(\REGISTERS[30][19] )
         );
  DLH_X1 \REGISTERS_reg[30][18]  ( .G(n325), .D(n383), .Q(\REGISTERS[30][18] )
         );
  DLH_X1 \REGISTERS_reg[30][17]  ( .G(n325), .D(n387), .Q(\REGISTERS[30][17] )
         );
  DLH_X1 \REGISTERS_reg[30][16]  ( .G(n325), .D(n391), .Q(\REGISTERS[30][16] )
         );
  DLH_X1 \REGISTERS_reg[30][15]  ( .G(n325), .D(n395), .Q(\REGISTERS[30][15] )
         );
  DLH_X1 \REGISTERS_reg[30][14]  ( .G(n325), .D(n399), .Q(\REGISTERS[30][14] )
         );
  DLH_X1 \REGISTERS_reg[30][13]  ( .G(n325), .D(n403), .Q(\REGISTERS[30][13] )
         );
  DLH_X1 \REGISTERS_reg[30][12]  ( .G(n325), .D(n407), .Q(\REGISTERS[30][12] )
         );
  DLH_X1 \REGISTERS_reg[30][11]  ( .G(n325), .D(n411), .Q(\REGISTERS[30][11] )
         );
  DLH_X1 \REGISTERS_reg[30][10]  ( .G(n325), .D(n415), .Q(\REGISTERS[30][10] )
         );
  DLH_X1 \REGISTERS_reg[30][9]  ( .G(n324), .D(n419), .Q(\REGISTERS[30][9] )
         );
  DLH_X1 \REGISTERS_reg[30][8]  ( .G(n324), .D(n423), .Q(\REGISTERS[30][8] )
         );
  DLH_X1 \REGISTERS_reg[30][7]  ( .G(n324), .D(n427), .Q(\REGISTERS[30][7] )
         );
  DLH_X1 \REGISTERS_reg[30][6]  ( .G(n324), .D(n431), .Q(\REGISTERS[30][6] )
         );
  DLH_X1 \REGISTERS_reg[30][5]  ( .G(n324), .D(n435), .Q(\REGISTERS[30][5] )
         );
  DLH_X1 \REGISTERS_reg[30][4]  ( .G(n324), .D(n439), .Q(\REGISTERS[30][4] )
         );
  DLH_X1 \REGISTERS_reg[30][3]  ( .G(n324), .D(n443), .Q(\REGISTERS[30][3] )
         );
  DLH_X1 \REGISTERS_reg[30][2]  ( .G(n324), .D(n447), .Q(\REGISTERS[30][2] )
         );
  DLH_X1 \REGISTERS_reg[30][1]  ( .G(n324), .D(n451), .Q(\REGISTERS[30][1] )
         );
  DLH_X1 \REGISTERS_reg[30][0]  ( .G(n324), .D(n455), .Q(\REGISTERS[30][0] )
         );
  DLH_X1 \REGISTERS_reg[31][31]  ( .G(n459), .D(n331), .Q(\REGISTERS[31][31] )
         );
  DLH_X1 \REGISTERS_reg[31][30]  ( .G(n459), .D(n335), .Q(\REGISTERS[31][30] )
         );
  DLH_X1 \REGISTERS_reg[31][29]  ( .G(n458), .D(n339), .Q(\REGISTERS[31][29] )
         );
  DLH_X1 \REGISTERS_reg[31][28]  ( .G(n458), .D(n343), .Q(\REGISTERS[31][28] )
         );
  DLH_X1 \REGISTERS_reg[31][27]  ( .G(n458), .D(n347), .Q(\REGISTERS[31][27] )
         );
  DLH_X1 \REGISTERS_reg[31][26]  ( .G(n458), .D(n351), .Q(\REGISTERS[31][26] )
         );
  DLH_X1 \REGISTERS_reg[31][25]  ( .G(n458), .D(n355), .Q(\REGISTERS[31][25] )
         );
  DLH_X1 \REGISTERS_reg[31][24]  ( .G(n458), .D(n359), .Q(\REGISTERS[31][24] )
         );
  DLH_X1 \REGISTERS_reg[31][23]  ( .G(n458), .D(n363), .Q(\REGISTERS[31][23] )
         );
  DLH_X1 \REGISTERS_reg[31][22]  ( .G(n458), .D(n367), .Q(\REGISTERS[31][22] )
         );
  DLH_X1 \REGISTERS_reg[31][21]  ( .G(n458), .D(n371), .Q(\REGISTERS[31][21] )
         );
  DLH_X1 \REGISTERS_reg[31][20]  ( .G(n458), .D(n375), .Q(\REGISTERS[31][20] )
         );
  DLH_X1 \REGISTERS_reg[31][19]  ( .G(n457), .D(n379), .Q(\REGISTERS[31][19] )
         );
  DLH_X1 \REGISTERS_reg[31][18]  ( .G(n457), .D(n383), .Q(\REGISTERS[31][18] )
         );
  DLH_X1 \REGISTERS_reg[31][17]  ( .G(n457), .D(n387), .Q(\REGISTERS[31][17] )
         );
  DLH_X1 \REGISTERS_reg[31][16]  ( .G(n457), .D(n391), .Q(\REGISTERS[31][16] )
         );
  DLH_X1 \REGISTERS_reg[31][15]  ( .G(n457), .D(n395), .Q(\REGISTERS[31][15] )
         );
  DLH_X1 \REGISTERS_reg[31][14]  ( .G(n457), .D(n399), .Q(\REGISTERS[31][14] )
         );
  DLH_X1 \REGISTERS_reg[31][13]  ( .G(n457), .D(n403), .Q(\REGISTERS[31][13] )
         );
  DLH_X1 \REGISTERS_reg[31][12]  ( .G(n457), .D(n407), .Q(\REGISTERS[31][12] )
         );
  DLH_X1 \REGISTERS_reg[31][11]  ( .G(n457), .D(n411), .Q(\REGISTERS[31][11] )
         );
  DLH_X1 \REGISTERS_reg[31][10]  ( .G(n457), .D(n415), .Q(\REGISTERS[31][10] )
         );
  DLH_X1 \REGISTERS_reg[31][9]  ( .G(n456), .D(n419), .Q(\REGISTERS[31][9] )
         );
  DLH_X1 \REGISTERS_reg[31][8]  ( .G(n456), .D(n423), .Q(\REGISTERS[31][8] )
         );
  DLH_X1 \REGISTERS_reg[31][7]  ( .G(n456), .D(n427), .Q(\REGISTERS[31][7] )
         );
  DLH_X1 \REGISTERS_reg[31][6]  ( .G(n456), .D(n431), .Q(\REGISTERS[31][6] )
         );
  DLH_X1 \REGISTERS_reg[31][5]  ( .G(n456), .D(n435), .Q(\REGISTERS[31][5] )
         );
  DLH_X1 \REGISTERS_reg[31][4]  ( .G(n456), .D(n439), .Q(\REGISTERS[31][4] )
         );
  DLH_X1 \REGISTERS_reg[31][3]  ( .G(n456), .D(n443), .Q(\REGISTERS[31][3] )
         );
  DLH_X1 \REGISTERS_reg[31][2]  ( .G(n456), .D(n447), .Q(\REGISTERS[31][2] )
         );
  DLH_X1 \REGISTERS_reg[31][1]  ( .G(n456), .D(n451), .Q(\REGISTERS[31][1] )
         );
  DLH_X1 \REGISTERS_reg[31][0]  ( .G(n456), .D(n455), .Q(\REGISTERS[31][0] )
         );
  DLH_X1 \OUT1_reg[31]  ( .G(n200), .D(N408), .Q(OUT1[31]) );
  DLH_X1 \OUT1_reg[30]  ( .G(n200), .D(N407), .Q(OUT1[30]) );
  DLH_X1 \OUT1_reg[29]  ( .G(n200), .D(N406), .Q(OUT1[29]) );
  DLH_X1 \OUT1_reg[28]  ( .G(n200), .D(N405), .Q(OUT1[28]) );
  DLH_X1 \OUT1_reg[27]  ( .G(n200), .D(N404), .Q(OUT1[27]) );
  DLH_X1 \OUT1_reg[26]  ( .G(n200), .D(N403), .Q(OUT1[26]) );
  DLH_X1 \OUT1_reg[25]  ( .G(n200), .D(N402), .Q(OUT1[25]) );
  DLH_X1 \OUT1_reg[24]  ( .G(n200), .D(N401), .Q(OUT1[24]) );
  DLH_X1 \OUT1_reg[23]  ( .G(n200), .D(N400), .Q(OUT1[23]) );
  DLH_X1 \OUT1_reg[22]  ( .G(n200), .D(N399), .Q(OUT1[22]) );
  DLH_X1 \OUT1_reg[21]  ( .G(n201), .D(N398), .Q(OUT1[21]) );
  DLH_X1 \OUT1_reg[20]  ( .G(n201), .D(N397), .Q(OUT1[20]) );
  DLH_X1 \OUT1_reg[19]  ( .G(n201), .D(N396), .Q(OUT1[19]) );
  DLH_X1 \OUT1_reg[18]  ( .G(n201), .D(N395), .Q(OUT1[18]) );
  DLH_X1 \OUT1_reg[17]  ( .G(n201), .D(N394), .Q(OUT1[17]) );
  DLH_X1 \OUT1_reg[16]  ( .G(n201), .D(N393), .Q(OUT1[16]) );
  DLH_X1 \OUT1_reg[15]  ( .G(n201), .D(N392), .Q(OUT1[15]) );
  DLH_X1 \OUT1_reg[14]  ( .G(n201), .D(N391), .Q(OUT1[14]) );
  DLH_X1 \OUT1_reg[13]  ( .G(n201), .D(N390), .Q(OUT1[13]) );
  DLH_X1 \OUT1_reg[12]  ( .G(n201), .D(N389), .Q(OUT1[12]) );
  DLH_X1 \OUT1_reg[11]  ( .G(n202), .D(N388), .Q(OUT1[11]) );
  DLH_X1 \OUT1_reg[10]  ( .G(n202), .D(N387), .Q(OUT1[10]) );
  DLH_X1 \OUT1_reg[9]  ( .G(n202), .D(N386), .Q(OUT1[9]) );
  DLH_X1 \OUT1_reg[8]  ( .G(n202), .D(N385), .Q(OUT1[8]) );
  DLH_X1 \OUT1_reg[7]  ( .G(n202), .D(N384), .Q(OUT1[7]) );
  DLH_X1 \OUT1_reg[6]  ( .G(n202), .D(N383), .Q(OUT1[6]) );
  DLH_X1 \OUT1_reg[5]  ( .G(n202), .D(N382), .Q(OUT1[5]) );
  DLH_X1 \OUT1_reg[4]  ( .G(n202), .D(N381), .Q(OUT1[4]) );
  DLH_X1 \OUT1_reg[3]  ( .G(n202), .D(N380), .Q(OUT1[3]) );
  DLH_X1 \OUT1_reg[2]  ( .G(n202), .D(N379), .Q(OUT1[2]) );
  DLH_X1 \OUT1_reg[1]  ( .G(n203), .D(N378), .Q(OUT1[1]) );
  DLH_X1 \OUT1_reg[0]  ( .G(n203), .D(N377), .Q(OUT1[0]) );
  DLH_X1 \OUT2_reg[31]  ( .G(n196), .D(N441), .Q(OUT2[31]) );
  DLH_X1 \OUT2_reg[30]  ( .G(n196), .D(N440), .Q(OUT2[30]) );
  DLH_X1 \OUT2_reg[29]  ( .G(n196), .D(N439), .Q(OUT2[29]) );
  DLH_X1 \OUT2_reg[28]  ( .G(n196), .D(N438), .Q(OUT2[28]) );
  DLH_X1 \OUT2_reg[27]  ( .G(n196), .D(N437), .Q(OUT2[27]) );
  DLH_X1 \OUT2_reg[26]  ( .G(n196), .D(N436), .Q(OUT2[26]) );
  DLH_X1 \OUT2_reg[25]  ( .G(n196), .D(N435), .Q(OUT2[25]) );
  DLH_X1 \OUT2_reg[24]  ( .G(n196), .D(N434), .Q(OUT2[24]) );
  DLH_X1 \OUT2_reg[23]  ( .G(n196), .D(N433), .Q(OUT2[23]) );
  DLH_X1 \OUT2_reg[22]  ( .G(n196), .D(N432), .Q(OUT2[22]) );
  DLH_X1 \OUT2_reg[21]  ( .G(n197), .D(N431), .Q(OUT2[21]) );
  DLH_X1 \OUT2_reg[20]  ( .G(n197), .D(N430), .Q(OUT2[20]) );
  DLH_X1 \OUT2_reg[19]  ( .G(n197), .D(N429), .Q(OUT2[19]) );
  DLH_X1 \OUT2_reg[18]  ( .G(n197), .D(N428), .Q(OUT2[18]) );
  DLH_X1 \OUT2_reg[17]  ( .G(n197), .D(N427), .Q(OUT2[17]) );
  DLH_X1 \OUT2_reg[16]  ( .G(n197), .D(N426), .Q(OUT2[16]) );
  DLH_X1 \OUT2_reg[15]  ( .G(n197), .D(N425), .Q(OUT2[15]) );
  DLH_X1 \OUT2_reg[14]  ( .G(n197), .D(N424), .Q(OUT2[14]) );
  DLH_X1 \OUT2_reg[13]  ( .G(n197), .D(N423), .Q(OUT2[13]) );
  DLH_X1 \OUT2_reg[12]  ( .G(n197), .D(N422), .Q(OUT2[12]) );
  DLH_X1 \OUT2_reg[11]  ( .G(n198), .D(N421), .Q(OUT2[11]) );
  DLH_X1 \OUT2_reg[10]  ( .G(n198), .D(N420), .Q(OUT2[10]) );
  DLH_X1 \OUT2_reg[9]  ( .G(n198), .D(N419), .Q(OUT2[9]) );
  DLH_X1 \OUT2_reg[8]  ( .G(n198), .D(N418), .Q(OUT2[8]) );
  DLH_X1 \OUT2_reg[7]  ( .G(n198), .D(N417), .Q(OUT2[7]) );
  DLH_X1 \OUT2_reg[6]  ( .G(n198), .D(N416), .Q(OUT2[6]) );
  DLH_X1 \OUT2_reg[5]  ( .G(n198), .D(N415), .Q(OUT2[5]) );
  DLH_X1 \OUT2_reg[4]  ( .G(n198), .D(N414), .Q(OUT2[4]) );
  DLH_X1 \OUT2_reg[3]  ( .G(n198), .D(N413), .Q(OUT2[3]) );
  DLH_X1 \OUT2_reg[2]  ( .G(n198), .D(N412), .Q(OUT2[2]) );
  DLH_X1 \OUT2_reg[1]  ( .G(n199), .D(N411), .Q(OUT2[1]) );
  DLH_X1 \OUT2_reg[0]  ( .G(n199), .D(N410), .Q(OUT2[0]) );
  NAND3_X1 U1911 ( .A1(n2262), .A2(n2263), .A3(WR), .ZN(n1778) );
  NAND3_X1 U1912 ( .A1(WR), .A2(n2263), .A3(ADD_WR[3]), .ZN(n1787) );
  NAND3_X1 U1913 ( .A1(WR), .A2(n2262), .A3(ADD_WR[4]), .ZN(n1788) );
  NAND3_X1 U1914 ( .A1(n2260), .A2(n2261), .A3(ADD_WR[0]), .ZN(n1779) );
  NAND3_X1 U1915 ( .A1(n2259), .A2(n2261), .A3(ADD_WR[1]), .ZN(n1780) );
  NAND3_X1 U1916 ( .A1(ADD_WR[0]), .A2(n2261), .A3(ADD_WR[1]), .ZN(n1781) );
  NAND3_X1 U1917 ( .A1(n2259), .A2(n2260), .A3(ADD_WR[2]), .ZN(n1782) );
  NAND3_X1 U1918 ( .A1(ADD_WR[0]), .A2(n2260), .A3(ADD_WR[2]), .ZN(n1783) );
  NAND3_X1 U1919 ( .A1(ADD_WR[1]), .A2(n2259), .A3(ADD_WR[2]), .ZN(n1784) );
  NAND3_X1 U1920 ( .A1(n2260), .A2(n2261), .A3(n2259), .ZN(n1786) );
  NAND3_X1 U1921 ( .A1(ADD_WR[3]), .A2(WR), .A3(ADD_WR[4]), .ZN(n1789) );
  NAND3_X1 U1922 ( .A1(ADD_WR[1]), .A2(ADD_WR[0]), .A3(ADD_WR[2]), .ZN(n1785)
         );
  NOR2_X1 U3 ( .A1(n2253), .A2(ADD_RD2[1]), .ZN(n1130) );
  NOR2_X1 U4 ( .A1(n2257), .A2(ADD_RD1[1]), .ZN(n1755) );
  NOR2_X1 U5 ( .A1(ADD_RD2[1]), .A2(ADD_RD2[2]), .ZN(n1127) );
  BUF_X1 U6 ( .A(n549), .Z(n154) );
  BUF_X1 U7 ( .A(n549), .Z(n155) );
  BUF_X1 U8 ( .A(n1167), .Z(n76) );
  BUF_X1 U9 ( .A(n1191), .Z(n28) );
  BUF_X1 U10 ( .A(n1201), .Z(n4) );
  BUF_X1 U11 ( .A(n1167), .Z(n77) );
  BUF_X1 U12 ( .A(n1191), .Z(n29) );
  BUF_X1 U13 ( .A(n1201), .Z(n5) );
  BUF_X1 U14 ( .A(n1174), .Z(n60) );
  BUF_X1 U15 ( .A(n542), .Z(n172) );
  BUF_X1 U16 ( .A(n566), .Z(n124) );
  BUF_X1 U17 ( .A(n576), .Z(n100) );
  BUF_X1 U18 ( .A(n542), .Z(n173) );
  BUF_X1 U19 ( .A(n566), .Z(n125) );
  BUF_X1 U20 ( .A(n576), .Z(n101) );
  BUF_X1 U21 ( .A(n549), .Z(n156) );
  BUF_X1 U22 ( .A(n1167), .Z(n78) );
  BUF_X1 U23 ( .A(n1191), .Z(n30) );
  BUF_X1 U24 ( .A(n1201), .Z(n6) );
  BUF_X1 U25 ( .A(n542), .Z(n174) );
  BUF_X1 U26 ( .A(n566), .Z(n126) );
  BUF_X1 U27 ( .A(n576), .Z(n102) );
  BUF_X1 U28 ( .A(n1174), .Z(n58) );
  BUF_X1 U29 ( .A(n1174), .Z(n59) );
  INV_X1 U30 ( .A(n473), .ZN(n462) );
  INV_X1 U31 ( .A(n473), .ZN(n463) );
  INV_X1 U32 ( .A(n473), .ZN(n464) );
  BUF_X1 U33 ( .A(n1161), .Z(n91) );
  BUF_X1 U34 ( .A(n1166), .Z(n79) );
  BUF_X1 U35 ( .A(n1171), .Z(n67) );
  BUF_X1 U36 ( .A(n1176), .Z(n55) );
  BUF_X1 U37 ( .A(n1185), .Z(n43) );
  BUF_X1 U38 ( .A(n1190), .Z(n31) );
  BUF_X1 U39 ( .A(n1195), .Z(n19) );
  BUF_X1 U40 ( .A(n1200), .Z(n7) );
  BUF_X1 U41 ( .A(n1161), .Z(n92) );
  BUF_X1 U42 ( .A(n1166), .Z(n80) );
  BUF_X1 U43 ( .A(n1171), .Z(n68) );
  BUF_X1 U44 ( .A(n1176), .Z(n56) );
  BUF_X1 U45 ( .A(n1185), .Z(n44) );
  BUF_X1 U46 ( .A(n1190), .Z(n32) );
  BUF_X1 U47 ( .A(n1195), .Z(n20) );
  BUF_X1 U48 ( .A(n1200), .Z(n8) );
  BUF_X1 U49 ( .A(n1158), .Z(n97) );
  BUF_X1 U50 ( .A(n1182), .Z(n49) );
  BUF_X1 U51 ( .A(n1192), .Z(n25) );
  BUF_X1 U52 ( .A(n1168), .Z(n73) );
  BUF_X1 U53 ( .A(n1163), .Z(n85) );
  BUF_X1 U54 ( .A(n1187), .Z(n37) );
  BUF_X1 U55 ( .A(n1197), .Z(n13) );
  BUF_X1 U56 ( .A(n1173), .Z(n61) );
  BUF_X1 U57 ( .A(n534), .Z(n190) );
  BUF_X1 U58 ( .A(n539), .Z(n178) );
  BUF_X1 U59 ( .A(n544), .Z(n166) );
  BUF_X1 U60 ( .A(n558), .Z(n142) );
  BUF_X1 U61 ( .A(n563), .Z(n130) );
  BUF_X1 U62 ( .A(n568), .Z(n118) );
  BUF_X1 U63 ( .A(n573), .Z(n106) );
  BUF_X1 U64 ( .A(n534), .Z(n191) );
  BUF_X1 U65 ( .A(n539), .Z(n179) );
  BUF_X1 U66 ( .A(n544), .Z(n167) );
  BUF_X1 U67 ( .A(n558), .Z(n143) );
  BUF_X1 U68 ( .A(n563), .Z(n131) );
  BUF_X1 U69 ( .A(n568), .Z(n119) );
  BUF_X1 U70 ( .A(n573), .Z(n107) );
  BUF_X1 U71 ( .A(n1162), .Z(n88) );
  BUF_X1 U72 ( .A(n1172), .Z(n64) );
  BUF_X1 U73 ( .A(n1177), .Z(n52) );
  BUF_X1 U74 ( .A(n1186), .Z(n40) );
  BUF_X1 U75 ( .A(n1196), .Z(n16) );
  BUF_X1 U76 ( .A(n1162), .Z(n89) );
  BUF_X1 U77 ( .A(n1172), .Z(n65) );
  BUF_X1 U78 ( .A(n1177), .Z(n53) );
  BUF_X1 U79 ( .A(n1186), .Z(n41) );
  BUF_X1 U80 ( .A(n1196), .Z(n17) );
  BUF_X1 U81 ( .A(n1159), .Z(n96) );
  BUF_X1 U82 ( .A(n1183), .Z(n48) );
  BUF_X1 U83 ( .A(n1193), .Z(n24) );
  BUF_X1 U84 ( .A(n1169), .Z(n72) );
  BUF_X1 U85 ( .A(n1164), .Z(n84) );
  BUF_X1 U86 ( .A(n1188), .Z(n36) );
  BUF_X1 U87 ( .A(n1198), .Z(n12) );
  BUF_X1 U88 ( .A(n1161), .Z(n93) );
  BUF_X1 U89 ( .A(n1171), .Z(n69) );
  BUF_X1 U90 ( .A(n1166), .Z(n81) );
  BUF_X1 U91 ( .A(n1176), .Z(n57) );
  BUF_X1 U92 ( .A(n1185), .Z(n45) );
  BUF_X1 U93 ( .A(n1190), .Z(n33) );
  BUF_X1 U94 ( .A(n1195), .Z(n21) );
  BUF_X1 U95 ( .A(n1200), .Z(n9) );
  BUF_X1 U96 ( .A(n1158), .Z(n99) );
  BUF_X1 U97 ( .A(n1182), .Z(n51) );
  BUF_X1 U98 ( .A(n1192), .Z(n27) );
  BUF_X1 U99 ( .A(n1168), .Z(n75) );
  BUF_X1 U100 ( .A(n1163), .Z(n87) );
  BUF_X1 U101 ( .A(n1187), .Z(n39) );
  BUF_X1 U102 ( .A(n1197), .Z(n15) );
  BUF_X1 U103 ( .A(n1173), .Z(n63) );
  BUF_X1 U104 ( .A(n533), .Z(n193) );
  BUF_X1 U105 ( .A(n557), .Z(n145) );
  BUF_X1 U106 ( .A(n567), .Z(n121) );
  BUF_X1 U107 ( .A(n533), .Z(n194) );
  BUF_X1 U108 ( .A(n557), .Z(n146) );
  BUF_X1 U109 ( .A(n567), .Z(n122) );
  BUF_X1 U110 ( .A(n538), .Z(n181) );
  BUF_X1 U111 ( .A(n562), .Z(n133) );
  BUF_X1 U112 ( .A(n572), .Z(n109) );
  BUF_X1 U113 ( .A(n538), .Z(n182) );
  BUF_X1 U114 ( .A(n562), .Z(n134) );
  BUF_X1 U115 ( .A(n572), .Z(n110) );
  BUF_X1 U116 ( .A(n543), .Z(n169) );
  BUF_X1 U117 ( .A(n543), .Z(n170) );
  BUF_X1 U118 ( .A(n536), .Z(n187) );
  BUF_X1 U119 ( .A(n541), .Z(n175) );
  BUF_X1 U120 ( .A(n546), .Z(n163) );
  BUF_X1 U121 ( .A(n551), .Z(n151) );
  BUF_X1 U122 ( .A(n560), .Z(n139) );
  BUF_X1 U123 ( .A(n565), .Z(n127) );
  BUF_X1 U124 ( .A(n570), .Z(n115) );
  BUF_X1 U125 ( .A(n575), .Z(n103) );
  BUF_X1 U126 ( .A(n536), .Z(n188) );
  BUF_X1 U127 ( .A(n541), .Z(n176) );
  BUF_X1 U128 ( .A(n546), .Z(n164) );
  BUF_X1 U129 ( .A(n551), .Z(n152) );
  BUF_X1 U130 ( .A(n560), .Z(n140) );
  BUF_X1 U131 ( .A(n565), .Z(n128) );
  BUF_X1 U132 ( .A(n570), .Z(n116) );
  BUF_X1 U133 ( .A(n575), .Z(n104) );
  BUF_X1 U134 ( .A(n548), .Z(n157) );
  BUF_X1 U135 ( .A(n548), .Z(n158) );
  BUF_X1 U136 ( .A(n537), .Z(n184) );
  BUF_X1 U137 ( .A(n547), .Z(n160) );
  BUF_X1 U138 ( .A(n552), .Z(n148) );
  BUF_X1 U139 ( .A(n561), .Z(n136) );
  BUF_X1 U140 ( .A(n571), .Z(n112) );
  BUF_X1 U141 ( .A(n537), .Z(n185) );
  BUF_X1 U142 ( .A(n547), .Z(n161) );
  BUF_X1 U143 ( .A(n552), .Z(n149) );
  BUF_X1 U144 ( .A(n561), .Z(n137) );
  BUF_X1 U145 ( .A(n571), .Z(n113) );
  BUF_X1 U146 ( .A(n534), .Z(n192) );
  BUF_X1 U147 ( .A(n539), .Z(n180) );
  BUF_X1 U148 ( .A(n544), .Z(n168) );
  BUF_X1 U149 ( .A(n558), .Z(n144) );
  BUF_X1 U150 ( .A(n563), .Z(n132) );
  BUF_X1 U151 ( .A(n568), .Z(n120) );
  BUF_X1 U152 ( .A(n573), .Z(n108) );
  BUF_X1 U153 ( .A(n1162), .Z(n90) );
  BUF_X1 U154 ( .A(n1172), .Z(n66) );
  BUF_X1 U155 ( .A(n1177), .Z(n54) );
  BUF_X1 U156 ( .A(n1186), .Z(n42) );
  BUF_X1 U157 ( .A(n1196), .Z(n18) );
  BUF_X1 U158 ( .A(n533), .Z(n195) );
  BUF_X1 U159 ( .A(n557), .Z(n147) );
  BUF_X1 U160 ( .A(n567), .Z(n123) );
  BUF_X1 U161 ( .A(n538), .Z(n183) );
  BUF_X1 U162 ( .A(n562), .Z(n135) );
  BUF_X1 U163 ( .A(n572), .Z(n111) );
  BUF_X1 U164 ( .A(n543), .Z(n171) );
  BUF_X1 U165 ( .A(n536), .Z(n189) );
  BUF_X1 U166 ( .A(n541), .Z(n177) );
  BUF_X1 U167 ( .A(n546), .Z(n165) );
  BUF_X1 U168 ( .A(n551), .Z(n153) );
  BUF_X1 U169 ( .A(n560), .Z(n141) );
  BUF_X1 U170 ( .A(n565), .Z(n129) );
  BUF_X1 U171 ( .A(n570), .Z(n117) );
  BUF_X1 U172 ( .A(n575), .Z(n105) );
  BUF_X1 U173 ( .A(n548), .Z(n159) );
  BUF_X1 U174 ( .A(n537), .Z(n186) );
  BUF_X1 U175 ( .A(n547), .Z(n162) );
  BUF_X1 U176 ( .A(n552), .Z(n150) );
  BUF_X1 U177 ( .A(n561), .Z(n138) );
  BUF_X1 U178 ( .A(n571), .Z(n114) );
  BUF_X1 U179 ( .A(n1159), .Z(n94) );
  BUF_X1 U180 ( .A(n1183), .Z(n46) );
  BUF_X1 U181 ( .A(n1193), .Z(n22) );
  BUF_X1 U182 ( .A(n1159), .Z(n95) );
  BUF_X1 U183 ( .A(n1183), .Z(n47) );
  BUF_X1 U184 ( .A(n1193), .Z(n23) );
  BUF_X1 U185 ( .A(n1169), .Z(n70) );
  BUF_X1 U186 ( .A(n1169), .Z(n71) );
  BUF_X1 U187 ( .A(n1164), .Z(n82) );
  BUF_X1 U188 ( .A(n1188), .Z(n34) );
  BUF_X1 U189 ( .A(n1198), .Z(n10) );
  BUF_X1 U190 ( .A(n1164), .Z(n83) );
  BUF_X1 U191 ( .A(n1188), .Z(n35) );
  BUF_X1 U192 ( .A(n1198), .Z(n11) );
  BUF_X1 U193 ( .A(n1158), .Z(n98) );
  BUF_X1 U194 ( .A(n1182), .Z(n50) );
  BUF_X1 U195 ( .A(n1192), .Z(n26) );
  BUF_X1 U196 ( .A(n1168), .Z(n74) );
  BUF_X1 U197 ( .A(n1163), .Z(n86) );
  BUF_X1 U198 ( .A(n1173), .Z(n62) );
  BUF_X1 U199 ( .A(n1187), .Z(n38) );
  BUF_X1 U200 ( .A(n1197), .Z(n14) );
  NAND2_X1 U201 ( .A1(n1758), .A2(n1754), .ZN(n1174) );
  AND2_X1 U202 ( .A1(n1124), .A2(n1129), .ZN(n542) );
  AND2_X1 U203 ( .A1(n1142), .A2(n1129), .ZN(n566) );
  AND2_X1 U204 ( .A1(n1147), .A2(n1129), .ZN(n576) );
  NAND2_X1 U205 ( .A1(n1133), .A2(n1129), .ZN(n549) );
  AND2_X1 U206 ( .A1(n1749), .A2(n1754), .ZN(n1167) );
  AND2_X1 U207 ( .A1(n1767), .A2(n1754), .ZN(n1191) );
  AND2_X1 U208 ( .A1(n1772), .A2(n1754), .ZN(n1201) );
  NOR2_X1 U209 ( .A1(n2253), .A2(n2252), .ZN(n1129) );
  NOR2_X1 U210 ( .A1(n2257), .A2(n2256), .ZN(n1754) );
  NAND2_X1 U211 ( .A1(n1752), .A2(n1758), .ZN(n1169) );
  NAND2_X1 U212 ( .A1(n1752), .A2(n1759), .ZN(n1168) );
  NAND2_X1 U213 ( .A1(n1749), .A2(n1752), .ZN(n1159) );
  NAND2_X1 U214 ( .A1(n1767), .A2(n1752), .ZN(n1183) );
  NAND2_X1 U215 ( .A1(n1772), .A2(n1752), .ZN(n1193) );
  NAND2_X1 U216 ( .A1(n1751), .A2(n1752), .ZN(n1158) );
  NAND2_X1 U217 ( .A1(n1768), .A2(n1752), .ZN(n1182) );
  NAND2_X1 U218 ( .A1(n1773), .A2(n1752), .ZN(n1192) );
  NAND2_X1 U219 ( .A1(n1127), .A2(n1134), .ZN(n543) );
  NAND2_X1 U220 ( .A1(n1127), .A2(n1133), .ZN(n544) );
  NAND2_X1 U221 ( .A1(n1129), .A2(n1134), .ZN(n548) );
  NAND2_X1 U222 ( .A1(n1126), .A2(n1127), .ZN(n533) );
  NAND2_X1 U223 ( .A1(n1143), .A2(n1127), .ZN(n557) );
  NAND2_X1 U224 ( .A1(n1148), .A2(n1127), .ZN(n567) );
  NAND2_X1 U225 ( .A1(n1754), .A2(n1759), .ZN(n1173) );
  NAND2_X1 U226 ( .A1(n1126), .A2(n1130), .ZN(n538) );
  NAND2_X1 U227 ( .A1(n1143), .A2(n1130), .ZN(n562) );
  NAND2_X1 U228 ( .A1(n1148), .A2(n1130), .ZN(n572) );
  NAND2_X1 U229 ( .A1(n1749), .A2(n1755), .ZN(n1164) );
  NAND2_X1 U230 ( .A1(n1767), .A2(n1755), .ZN(n1188) );
  NAND2_X1 U231 ( .A1(n1772), .A2(n1755), .ZN(n1198) );
  NAND2_X1 U232 ( .A1(n1751), .A2(n1755), .ZN(n1163) );
  NAND2_X1 U233 ( .A1(n1768), .A2(n1755), .ZN(n1187) );
  NAND2_X1 U234 ( .A1(n1773), .A2(n1755), .ZN(n1197) );
  BUF_X1 U235 ( .A(n461), .Z(n473) );
  NAND2_X1 U236 ( .A1(n1124), .A2(n1127), .ZN(n534) );
  NAND2_X1 U237 ( .A1(n1142), .A2(n1127), .ZN(n558) );
  NAND2_X1 U238 ( .A1(n1147), .A2(n1127), .ZN(n568) );
  AND2_X1 U239 ( .A1(n1136), .A2(n2251), .ZN(n1133) );
  AND2_X1 U240 ( .A1(n1761), .A2(n2255), .ZN(n1758) );
  AND2_X1 U241 ( .A1(n1145), .A2(n2251), .ZN(n1142) );
  AND2_X1 U242 ( .A1(n1150), .A2(n2251), .ZN(n1147) );
  AND2_X1 U243 ( .A1(n1770), .A2(n2255), .ZN(n1767) );
  AND2_X1 U244 ( .A1(n1775), .A2(n2255), .ZN(n1772) );
  AND2_X1 U245 ( .A1(n1131), .A2(n2251), .ZN(n1124) );
  AND2_X1 U246 ( .A1(n1756), .A2(n2255), .ZN(n1749) );
  NAND2_X1 U247 ( .A1(n1124), .A2(n1130), .ZN(n539) );
  NAND2_X1 U248 ( .A1(n1142), .A2(n1130), .ZN(n563) );
  NAND2_X1 U249 ( .A1(n1147), .A2(n1130), .ZN(n573) );
  AND2_X1 U250 ( .A1(n1130), .A2(n1134), .ZN(n551) );
  AND2_X1 U251 ( .A1(n1130), .A2(n1133), .ZN(n552) );
  AND2_X1 U252 ( .A1(n1125), .A2(n1134), .ZN(n546) );
  AND2_X1 U253 ( .A1(n1125), .A2(n1133), .ZN(n547) );
  AND2_X1 U254 ( .A1(n1126), .A2(n1129), .ZN(n541) );
  AND2_X1 U255 ( .A1(n1143), .A2(n1129), .ZN(n565) );
  AND2_X1 U256 ( .A1(n1148), .A2(n1129), .ZN(n575) );
  AND2_X1 U257 ( .A1(n1126), .A2(n1125), .ZN(n536) );
  AND2_X1 U258 ( .A1(n1124), .A2(n1125), .ZN(n537) );
  AND2_X1 U259 ( .A1(n1143), .A2(n1125), .ZN(n560) );
  AND2_X1 U260 ( .A1(n1142), .A2(n1125), .ZN(n561) );
  AND2_X1 U261 ( .A1(n1148), .A2(n1125), .ZN(n570) );
  AND2_X1 U262 ( .A1(n1147), .A2(n1125), .ZN(n571) );
  BUF_X1 U263 ( .A(n461), .Z(n471) );
  BUF_X1 U264 ( .A(n461), .Z(n470) );
  BUF_X1 U265 ( .A(n460), .Z(n469) );
  BUF_X1 U266 ( .A(n460), .Z(n468) );
  BUF_X1 U267 ( .A(n460), .Z(n467) );
  BUF_X1 U268 ( .A(n460), .Z(n466) );
  BUF_X1 U269 ( .A(n460), .Z(n465) );
  BUF_X1 U270 ( .A(n461), .Z(n472) );
  BUF_X1 U271 ( .A(n461), .Z(n474) );
  AND2_X1 U272 ( .A1(n1750), .A2(n1759), .ZN(n1171) );
  AND2_X1 U273 ( .A1(n1750), .A2(n1758), .ZN(n1172) );
  AND2_X1 U274 ( .A1(n1755), .A2(n1759), .ZN(n1176) );
  AND2_X1 U275 ( .A1(n1755), .A2(n1758), .ZN(n1177) );
  AND2_X1 U276 ( .A1(n1751), .A2(n1750), .ZN(n1161) );
  AND2_X1 U277 ( .A1(n1749), .A2(n1750), .ZN(n1162) );
  AND2_X1 U278 ( .A1(n1768), .A2(n1750), .ZN(n1185) );
  AND2_X1 U279 ( .A1(n1767), .A2(n1750), .ZN(n1186) );
  AND2_X1 U280 ( .A1(n1773), .A2(n1750), .ZN(n1195) );
  AND2_X1 U281 ( .A1(n1772), .A2(n1750), .ZN(n1196) );
  AND2_X1 U282 ( .A1(n1751), .A2(n1754), .ZN(n1166) );
  AND2_X1 U283 ( .A1(n1768), .A2(n1754), .ZN(n1190) );
  AND2_X1 U284 ( .A1(n1773), .A2(n1754), .ZN(n1200) );
  NAND2_X1 U285 ( .A1(n472), .A2(n1151), .ZN(N409) );
  NAND2_X1 U286 ( .A1(RD2), .A2(ENABLE), .ZN(n1151) );
  NAND2_X1 U287 ( .A1(n473), .A2(n1776), .ZN(N376) );
  NAND2_X1 U288 ( .A1(RD1), .A2(ENABLE), .ZN(n1776) );
  NOR2_X1 U289 ( .A1(n2252), .A2(ADD_RD2[2]), .ZN(n1125) );
  INV_X1 U290 ( .A(ADD_RD2[0]), .ZN(n2251) );
  BUF_X1 U291 ( .A(n1790), .Z(n2) );
  BUF_X1 U292 ( .A(n1790), .Z(n1) );
  INV_X1 U293 ( .A(ADD_RD2[1]), .ZN(n2252) );
  INV_X1 U294 ( .A(ADD_RD2[2]), .ZN(n2253) );
  BUF_X1 U295 ( .A(n1790), .Z(n3) );
  NOR2_X1 U296 ( .A1(ADD_RD2[3]), .A2(ADD_RD2[4]), .ZN(n1145) );
  NOR2_X1 U297 ( .A1(n2254), .A2(ADD_RD2[4]), .ZN(n1150) );
  INV_X1 U298 ( .A(ADD_RD1[0]), .ZN(n2255) );
  AND2_X1 U299 ( .A1(ADD_RD2[0]), .A2(n1136), .ZN(n1134) );
  INV_X1 U300 ( .A(ADD_RD2[3]), .ZN(n2254) );
  AND2_X1 U301 ( .A1(ADD_RD1[0]), .A2(n1761), .ZN(n1759) );
  AND2_X1 U302 ( .A1(n1131), .A2(ADD_RD2[0]), .ZN(n1126) );
  AND2_X1 U303 ( .A1(n1145), .A2(ADD_RD2[0]), .ZN(n1143) );
  AND2_X1 U304 ( .A1(n1150), .A2(ADD_RD2[0]), .ZN(n1148) );
  AND2_X1 U305 ( .A1(n1756), .A2(ADD_RD1[0]), .ZN(n1751) );
  AND2_X1 U306 ( .A1(n1770), .A2(ADD_RD1[0]), .ZN(n1768) );
  AND2_X1 U307 ( .A1(n1775), .A2(ADD_RD1[0]), .ZN(n1773) );
  NOR2_X1 U308 ( .A1(ADD_RD1[3]), .A2(ADD_RD1[4]), .ZN(n1770) );
  NOR2_X1 U309 ( .A1(n2258), .A2(ADD_RD1[4]), .ZN(n1775) );
  INV_X1 U310 ( .A(ADD_RD1[1]), .ZN(n2256) );
  BUF_X1 U311 ( .A(N313), .Z(n454) );
  BUF_X1 U312 ( .A(N314), .Z(n450) );
  BUF_X1 U313 ( .A(N315), .Z(n446) );
  BUF_X1 U314 ( .A(N316), .Z(n442) );
  BUF_X1 U315 ( .A(N317), .Z(n438) );
  BUF_X1 U316 ( .A(N318), .Z(n434) );
  BUF_X1 U317 ( .A(N319), .Z(n430) );
  BUF_X1 U318 ( .A(N320), .Z(n426) );
  BUF_X1 U319 ( .A(N321), .Z(n422) );
  BUF_X1 U320 ( .A(N322), .Z(n418) );
  BUF_X1 U321 ( .A(N323), .Z(n414) );
  BUF_X1 U322 ( .A(N324), .Z(n410) );
  BUF_X1 U323 ( .A(N325), .Z(n406) );
  BUF_X1 U324 ( .A(N326), .Z(n402) );
  BUF_X1 U325 ( .A(N327), .Z(n398) );
  BUF_X1 U326 ( .A(N328), .Z(n394) );
  BUF_X1 U327 ( .A(N329), .Z(n390) );
  BUF_X1 U328 ( .A(N330), .Z(n386) );
  BUF_X1 U329 ( .A(N331), .Z(n382) );
  BUF_X1 U330 ( .A(N332), .Z(n378) );
  BUF_X1 U331 ( .A(N333), .Z(n374) );
  BUF_X1 U332 ( .A(N334), .Z(n370) );
  BUF_X1 U333 ( .A(N335), .Z(n366) );
  BUF_X1 U334 ( .A(N336), .Z(n362) );
  BUF_X1 U335 ( .A(N337), .Z(n358) );
  BUF_X1 U336 ( .A(N338), .Z(n354) );
  BUF_X1 U337 ( .A(N339), .Z(n350) );
  BUF_X1 U338 ( .A(N340), .Z(n346) );
  BUF_X1 U339 ( .A(N341), .Z(n342) );
  BUF_X1 U340 ( .A(N342), .Z(n338) );
  BUF_X1 U341 ( .A(N343), .Z(n334) );
  BUF_X1 U342 ( .A(N344), .Z(n330) );
  BUF_X1 U343 ( .A(N313), .Z(n453) );
  BUF_X1 U344 ( .A(N314), .Z(n449) );
  BUF_X1 U345 ( .A(N315), .Z(n445) );
  BUF_X1 U346 ( .A(N316), .Z(n441) );
  BUF_X1 U347 ( .A(N317), .Z(n437) );
  BUF_X1 U348 ( .A(N318), .Z(n433) );
  BUF_X1 U349 ( .A(N319), .Z(n429) );
  BUF_X1 U350 ( .A(N320), .Z(n425) );
  BUF_X1 U351 ( .A(N321), .Z(n421) );
  BUF_X1 U352 ( .A(N322), .Z(n417) );
  BUF_X1 U353 ( .A(N323), .Z(n413) );
  BUF_X1 U354 ( .A(N324), .Z(n409) );
  BUF_X1 U355 ( .A(N325), .Z(n405) );
  BUF_X1 U356 ( .A(N326), .Z(n401) );
  BUF_X1 U357 ( .A(N327), .Z(n397) );
  BUF_X1 U358 ( .A(N328), .Z(n393) );
  BUF_X1 U359 ( .A(N329), .Z(n389) );
  BUF_X1 U360 ( .A(N330), .Z(n385) );
  BUF_X1 U361 ( .A(N331), .Z(n381) );
  BUF_X1 U362 ( .A(N332), .Z(n377) );
  BUF_X1 U363 ( .A(N333), .Z(n373) );
  BUF_X1 U364 ( .A(N334), .Z(n369) );
  BUF_X1 U365 ( .A(N335), .Z(n365) );
  BUF_X1 U366 ( .A(N336), .Z(n361) );
  BUF_X1 U367 ( .A(N337), .Z(n357) );
  BUF_X1 U368 ( .A(N338), .Z(n353) );
  BUF_X1 U369 ( .A(N339), .Z(n349) );
  BUF_X1 U370 ( .A(N340), .Z(n345) );
  BUF_X1 U371 ( .A(N341), .Z(n341) );
  BUF_X1 U372 ( .A(N342), .Z(n337) );
  BUF_X1 U373 ( .A(N343), .Z(n333) );
  BUF_X1 U374 ( .A(N344), .Z(n329) );
  BUF_X1 U375 ( .A(N313), .Z(n452) );
  BUF_X1 U376 ( .A(N314), .Z(n448) );
  BUF_X1 U377 ( .A(N315), .Z(n444) );
  BUF_X1 U378 ( .A(N316), .Z(n440) );
  BUF_X1 U379 ( .A(N317), .Z(n436) );
  BUF_X1 U380 ( .A(N318), .Z(n432) );
  BUF_X1 U381 ( .A(N319), .Z(n428) );
  BUF_X1 U382 ( .A(N320), .Z(n424) );
  BUF_X1 U383 ( .A(N321), .Z(n420) );
  BUF_X1 U384 ( .A(N322), .Z(n416) );
  BUF_X1 U385 ( .A(N323), .Z(n412) );
  BUF_X1 U386 ( .A(N324), .Z(n408) );
  BUF_X1 U387 ( .A(N325), .Z(n404) );
  BUF_X1 U388 ( .A(N326), .Z(n400) );
  BUF_X1 U389 ( .A(N327), .Z(n396) );
  BUF_X1 U390 ( .A(N328), .Z(n392) );
  BUF_X1 U391 ( .A(N329), .Z(n388) );
  BUF_X1 U392 ( .A(N330), .Z(n384) );
  BUF_X1 U393 ( .A(N331), .Z(n380) );
  BUF_X1 U394 ( .A(N332), .Z(n376) );
  BUF_X1 U395 ( .A(N333), .Z(n372) );
  BUF_X1 U396 ( .A(N334), .Z(n368) );
  BUF_X1 U397 ( .A(N335), .Z(n364) );
  BUF_X1 U398 ( .A(N336), .Z(n360) );
  BUF_X1 U399 ( .A(N337), .Z(n356) );
  BUF_X1 U400 ( .A(N338), .Z(n352) );
  BUF_X1 U401 ( .A(N339), .Z(n348) );
  BUF_X1 U402 ( .A(N340), .Z(n344) );
  BUF_X1 U403 ( .A(N341), .Z(n340) );
  BUF_X1 U404 ( .A(N342), .Z(n336) );
  BUF_X1 U405 ( .A(N343), .Z(n332) );
  BUF_X1 U406 ( .A(N344), .Z(n328) );
  INV_X1 U407 ( .A(ADD_RD1[3]), .ZN(n2258) );
  AND2_X1 U408 ( .A1(ADD_RD2[4]), .A2(ADD_RD2[3]), .ZN(n1136) );
  AND2_X1 U409 ( .A1(ADD_RD2[4]), .A2(n2254), .ZN(n1131) );
  AND2_X1 U410 ( .A1(ADD_RD1[4]), .A2(ADD_RD1[3]), .ZN(n1761) );
  AND2_X1 U411 ( .A1(ADD_RD1[4]), .A2(n2258), .ZN(n1756) );
  BUF_X1 U412 ( .A(RESET), .Z(n460) );
  BUF_X1 U413 ( .A(RESET), .Z(n461) );
  OAI21_X1 U414 ( .B1(n1778), .B2(n1785), .A(n466), .ZN(N368) );
  OAI21_X1 U415 ( .B1(n1778), .B2(n1784), .A(n466), .ZN(N369) );
  OAI21_X1 U416 ( .B1(n1778), .B2(n1783), .A(n466), .ZN(N370) );
  OAI21_X1 U417 ( .B1(n1778), .B2(n1782), .A(n465), .ZN(N371) );
  OAI21_X1 U418 ( .B1(n1778), .B2(n1781), .A(n465), .ZN(N372) );
  OAI21_X1 U419 ( .B1(n1778), .B2(n1780), .A(n465), .ZN(N373) );
  OAI21_X1 U420 ( .B1(n1778), .B2(n1779), .A(n465), .ZN(N374) );
  OAI21_X1 U421 ( .B1(n1785), .B2(n1789), .A(n472), .ZN(N312) );
  OAI21_X1 U422 ( .B1(n1784), .B2(n1789), .A(n470), .ZN(N345) );
  OAI21_X1 U423 ( .B1(n1783), .B2(n1789), .A(n472), .ZN(N346) );
  OAI21_X1 U424 ( .B1(n1782), .B2(n1789), .A(n472), .ZN(N347) );
  OAI21_X1 U425 ( .B1(n1781), .B2(n1789), .A(n471), .ZN(N348) );
  OAI21_X1 U426 ( .B1(n1780), .B2(n1789), .A(n471), .ZN(N349) );
  OAI21_X1 U427 ( .B1(n1779), .B2(n1789), .A(n471), .ZN(N350) );
  OAI21_X1 U428 ( .B1(n1786), .B2(n1789), .A(n471), .ZN(N351) );
  OAI21_X1 U429 ( .B1(n1785), .B2(n1787), .A(n468), .ZN(N360) );
  OAI21_X1 U430 ( .B1(n1784), .B2(n1787), .A(n468), .ZN(N361) );
  OAI21_X1 U431 ( .B1(n1783), .B2(n1787), .A(n468), .ZN(N362) );
  OAI21_X1 U432 ( .B1(n1782), .B2(n1787), .A(n467), .ZN(N363) );
  OAI21_X1 U433 ( .B1(n1781), .B2(n1787), .A(n467), .ZN(N364) );
  OAI21_X1 U434 ( .B1(n1780), .B2(n1787), .A(n467), .ZN(N365) );
  OAI21_X1 U435 ( .B1(n1779), .B2(n1787), .A(n467), .ZN(N366) );
  OAI21_X1 U436 ( .B1(n1786), .B2(n1787), .A(n466), .ZN(N367) );
  OAI21_X1 U437 ( .B1(n1785), .B2(n1788), .A(n470), .ZN(N352) );
  OAI21_X1 U438 ( .B1(n1784), .B2(n1788), .A(n470), .ZN(N353) );
  OAI21_X1 U439 ( .B1(n1783), .B2(n1788), .A(n470), .ZN(N354) );
  OAI21_X1 U440 ( .B1(n1782), .B2(n1788), .A(n469), .ZN(N355) );
  OAI21_X1 U441 ( .B1(n1781), .B2(n1788), .A(n469), .ZN(N356) );
  OAI21_X1 U442 ( .B1(n1780), .B2(n1788), .A(n469), .ZN(N357) );
  OAI21_X1 U443 ( .B1(n1779), .B2(n1788), .A(n469), .ZN(N358) );
  OAI21_X1 U444 ( .B1(n1786), .B2(n1788), .A(n468), .ZN(N359) );
  AOI21_X1 U445 ( .B1(n1117), .B2(n1118), .A(n464), .ZN(N410) );
  NOR4_X1 U446 ( .A1(n1137), .A2(n1138), .A3(n1139), .A4(n1140), .ZN(n1117) );
  NOR4_X1 U447 ( .A1(n1119), .A2(n1120), .A3(n1121), .A4(n1122), .ZN(n1118) );
  OAI221_X1 U448 ( .B1(n109), .B2(n1994), .C1(n106), .C2(n1962), .A(n1149), 
        .ZN(n1137) );
  AOI21_X1 U449 ( .B1(n1742), .B2(n1743), .A(n462), .ZN(N377) );
  NOR4_X1 U450 ( .A1(n1762), .A2(n1763), .A3(n1764), .A4(n1765), .ZN(n1742) );
  NOR4_X1 U451 ( .A1(n1744), .A2(n1745), .A3(n1746), .A4(n1747), .ZN(n1743) );
  OAI221_X1 U452 ( .B1(n1994), .B2(n13), .C1(n1962), .C2(n10), .A(n1774), .ZN(
        n1762) );
  AOI21_X1 U453 ( .B1(n1724), .B2(n1725), .A(n462), .ZN(N378) );
  NOR4_X1 U454 ( .A1(n1734), .A2(n1735), .A3(n1736), .A4(n1737), .ZN(n1724) );
  NOR4_X1 U455 ( .A1(n1726), .A2(n1727), .A3(n1728), .A4(n1729), .ZN(n1725) );
  OAI221_X1 U456 ( .B1(n1993), .B2(n13), .C1(n1961), .C2(n10), .A(n1741), .ZN(
        n1734) );
  AOI21_X1 U457 ( .B1(n1706), .B2(n1707), .A(n462), .ZN(N379) );
  NOR4_X1 U458 ( .A1(n1716), .A2(n1717), .A3(n1718), .A4(n1719), .ZN(n1706) );
  NOR4_X1 U459 ( .A1(n1708), .A2(n1709), .A3(n1710), .A4(n1711), .ZN(n1707) );
  OAI221_X1 U460 ( .B1(n1992), .B2(n13), .C1(n1960), .C2(n10), .A(n1723), .ZN(
        n1716) );
  AOI21_X1 U461 ( .B1(n1688), .B2(n1689), .A(n462), .ZN(N380) );
  NOR4_X1 U462 ( .A1(n1698), .A2(n1699), .A3(n1700), .A4(n1701), .ZN(n1688) );
  NOR4_X1 U463 ( .A1(n1690), .A2(n1691), .A3(n1692), .A4(n1693), .ZN(n1689) );
  OAI221_X1 U464 ( .B1(n1991), .B2(n13), .C1(n1959), .C2(n10), .A(n1705), .ZN(
        n1698) );
  AOI21_X1 U465 ( .B1(n1670), .B2(n1671), .A(n462), .ZN(N381) );
  NOR4_X1 U466 ( .A1(n1680), .A2(n1681), .A3(n1682), .A4(n1683), .ZN(n1670) );
  NOR4_X1 U467 ( .A1(n1672), .A2(n1673), .A3(n1674), .A4(n1675), .ZN(n1671) );
  OAI221_X1 U468 ( .B1(n1990), .B2(n13), .C1(n1958), .C2(n10), .A(n1687), .ZN(
        n1680) );
  AOI21_X1 U469 ( .B1(n1652), .B2(n1653), .A(n462), .ZN(N382) );
  NOR4_X1 U470 ( .A1(n1662), .A2(n1663), .A3(n1664), .A4(n1665), .ZN(n1652) );
  NOR4_X1 U471 ( .A1(n1654), .A2(n1655), .A3(n1656), .A4(n1657), .ZN(n1653) );
  OAI221_X1 U472 ( .B1(n1989), .B2(n13), .C1(n1957), .C2(n10), .A(n1669), .ZN(
        n1662) );
  AOI21_X1 U473 ( .B1(n1634), .B2(n1635), .A(n462), .ZN(N383) );
  NOR4_X1 U474 ( .A1(n1644), .A2(n1645), .A3(n1646), .A4(n1647), .ZN(n1634) );
  NOR4_X1 U475 ( .A1(n1636), .A2(n1637), .A3(n1638), .A4(n1639), .ZN(n1635) );
  OAI221_X1 U476 ( .B1(n1988), .B2(n13), .C1(n1956), .C2(n10), .A(n1651), .ZN(
        n1644) );
  AOI21_X1 U477 ( .B1(n1616), .B2(n1617), .A(n462), .ZN(N384) );
  NOR4_X1 U478 ( .A1(n1626), .A2(n1627), .A3(n1628), .A4(n1629), .ZN(n1616) );
  NOR4_X1 U479 ( .A1(n1618), .A2(n1619), .A3(n1620), .A4(n1621), .ZN(n1617) );
  OAI221_X1 U480 ( .B1(n1987), .B2(n13), .C1(n1955), .C2(n10), .A(n1633), .ZN(
        n1626) );
  AOI21_X1 U481 ( .B1(n1598), .B2(n1599), .A(n462), .ZN(N385) );
  NOR4_X1 U482 ( .A1(n1608), .A2(n1609), .A3(n1610), .A4(n1611), .ZN(n1598) );
  NOR4_X1 U483 ( .A1(n1600), .A2(n1601), .A3(n1602), .A4(n1603), .ZN(n1599) );
  OAI221_X1 U484 ( .B1(n1986), .B2(n13), .C1(n1954), .C2(n10), .A(n1615), .ZN(
        n1608) );
  AOI21_X1 U485 ( .B1(n1580), .B2(n1581), .A(n462), .ZN(N386) );
  NOR4_X1 U486 ( .A1(n1590), .A2(n1591), .A3(n1592), .A4(n1593), .ZN(n1580) );
  NOR4_X1 U487 ( .A1(n1582), .A2(n1583), .A3(n1584), .A4(n1585), .ZN(n1581) );
  OAI221_X1 U488 ( .B1(n1985), .B2(n13), .C1(n1953), .C2(n10), .A(n1597), .ZN(
        n1590) );
  AOI21_X1 U489 ( .B1(n1562), .B2(n1563), .A(n462), .ZN(N387) );
  NOR4_X1 U490 ( .A1(n1572), .A2(n1573), .A3(n1574), .A4(n1575), .ZN(n1562) );
  NOR4_X1 U491 ( .A1(n1564), .A2(n1565), .A3(n1566), .A4(n1567), .ZN(n1563) );
  OAI221_X1 U492 ( .B1(n1984), .B2(n13), .C1(n1952), .C2(n10), .A(n1579), .ZN(
        n1572) );
  AOI21_X1 U493 ( .B1(n1544), .B2(n1545), .A(n463), .ZN(N388) );
  NOR4_X1 U494 ( .A1(n1554), .A2(n1555), .A3(n1556), .A4(n1557), .ZN(n1544) );
  NOR4_X1 U495 ( .A1(n1546), .A2(n1547), .A3(n1548), .A4(n1549), .ZN(n1545) );
  OAI221_X1 U496 ( .B1(n1983), .B2(n14), .C1(n1951), .C2(n11), .A(n1561), .ZN(
        n1554) );
  AOI21_X1 U497 ( .B1(n1526), .B2(n1527), .A(n463), .ZN(N389) );
  NOR4_X1 U498 ( .A1(n1536), .A2(n1537), .A3(n1538), .A4(n1539), .ZN(n1526) );
  NOR4_X1 U499 ( .A1(n1528), .A2(n1529), .A3(n1530), .A4(n1531), .ZN(n1527) );
  OAI221_X1 U500 ( .B1(n1982), .B2(n14), .C1(n1950), .C2(n11), .A(n1543), .ZN(
        n1536) );
  AOI21_X1 U501 ( .B1(n1508), .B2(n1509), .A(n463), .ZN(N390) );
  NOR4_X1 U502 ( .A1(n1518), .A2(n1519), .A3(n1520), .A4(n1521), .ZN(n1508) );
  NOR4_X1 U503 ( .A1(n1510), .A2(n1511), .A3(n1512), .A4(n1513), .ZN(n1509) );
  OAI221_X1 U504 ( .B1(n1981), .B2(n14), .C1(n1949), .C2(n11), .A(n1525), .ZN(
        n1518) );
  AOI21_X1 U505 ( .B1(n1490), .B2(n1491), .A(n463), .ZN(N391) );
  NOR4_X1 U506 ( .A1(n1500), .A2(n1501), .A3(n1502), .A4(n1503), .ZN(n1490) );
  NOR4_X1 U507 ( .A1(n1492), .A2(n1493), .A3(n1494), .A4(n1495), .ZN(n1491) );
  OAI221_X1 U508 ( .B1(n1980), .B2(n14), .C1(n1948), .C2(n11), .A(n1507), .ZN(
        n1500) );
  AOI21_X1 U509 ( .B1(n1472), .B2(n1473), .A(n463), .ZN(N392) );
  NOR4_X1 U510 ( .A1(n1482), .A2(n1483), .A3(n1484), .A4(n1485), .ZN(n1472) );
  NOR4_X1 U511 ( .A1(n1474), .A2(n1475), .A3(n1476), .A4(n1477), .ZN(n1473) );
  OAI221_X1 U512 ( .B1(n1979), .B2(n14), .C1(n1947), .C2(n11), .A(n1489), .ZN(
        n1482) );
  AOI21_X1 U513 ( .B1(n1454), .B2(n1455), .A(n463), .ZN(N393) );
  NOR4_X1 U514 ( .A1(n1464), .A2(n1465), .A3(n1466), .A4(n1467), .ZN(n1454) );
  NOR4_X1 U515 ( .A1(n1456), .A2(n1457), .A3(n1458), .A4(n1459), .ZN(n1455) );
  OAI221_X1 U516 ( .B1(n1978), .B2(n14), .C1(n1946), .C2(n11), .A(n1471), .ZN(
        n1464) );
  AOI21_X1 U517 ( .B1(n1436), .B2(n1437), .A(n463), .ZN(N394) );
  NOR4_X1 U518 ( .A1(n1446), .A2(n1447), .A3(n1448), .A4(n1449), .ZN(n1436) );
  NOR4_X1 U519 ( .A1(n1438), .A2(n1439), .A3(n1440), .A4(n1441), .ZN(n1437) );
  OAI221_X1 U520 ( .B1(n1977), .B2(n14), .C1(n1945), .C2(n11), .A(n1453), .ZN(
        n1446) );
  AOI21_X1 U521 ( .B1(n1418), .B2(n1419), .A(n463), .ZN(N395) );
  NOR4_X1 U522 ( .A1(n1428), .A2(n1429), .A3(n1430), .A4(n1431), .ZN(n1418) );
  NOR4_X1 U523 ( .A1(n1420), .A2(n1421), .A3(n1422), .A4(n1423), .ZN(n1419) );
  OAI221_X1 U524 ( .B1(n1976), .B2(n14), .C1(n1944), .C2(n11), .A(n1435), .ZN(
        n1428) );
  AOI21_X1 U525 ( .B1(n1400), .B2(n1401), .A(n463), .ZN(N396) );
  NOR4_X1 U526 ( .A1(n1410), .A2(n1411), .A3(n1412), .A4(n1413), .ZN(n1400) );
  NOR4_X1 U527 ( .A1(n1402), .A2(n1403), .A3(n1404), .A4(n1405), .ZN(n1401) );
  OAI221_X1 U528 ( .B1(n1975), .B2(n14), .C1(n1943), .C2(n11), .A(n1417), .ZN(
        n1410) );
  AOI21_X1 U529 ( .B1(n1382), .B2(n1383), .A(n463), .ZN(N397) );
  NOR4_X1 U530 ( .A1(n1392), .A2(n1393), .A3(n1394), .A4(n1395), .ZN(n1382) );
  NOR4_X1 U531 ( .A1(n1384), .A2(n1385), .A3(n1386), .A4(n1387), .ZN(n1383) );
  OAI221_X1 U532 ( .B1(n1974), .B2(n14), .C1(n1942), .C2(n11), .A(n1399), .ZN(
        n1392) );
  AOI21_X1 U533 ( .B1(n1364), .B2(n1365), .A(n463), .ZN(N398) );
  NOR4_X1 U534 ( .A1(n1374), .A2(n1375), .A3(n1376), .A4(n1377), .ZN(n1364) );
  NOR4_X1 U535 ( .A1(n1366), .A2(n1367), .A3(n1368), .A4(n1369), .ZN(n1365) );
  OAI221_X1 U536 ( .B1(n1973), .B2(n14), .C1(n1941), .C2(n11), .A(n1381), .ZN(
        n1374) );
  AOI21_X1 U537 ( .B1(n1346), .B2(n1347), .A(n464), .ZN(N399) );
  NOR4_X1 U538 ( .A1(n1356), .A2(n1357), .A3(n1358), .A4(n1359), .ZN(n1346) );
  NOR4_X1 U539 ( .A1(n1348), .A2(n1349), .A3(n1350), .A4(n1351), .ZN(n1347) );
  OAI221_X1 U540 ( .B1(n1972), .B2(n15), .C1(n1940), .C2(n12), .A(n1363), .ZN(
        n1356) );
  AOI21_X1 U541 ( .B1(n1328), .B2(n1329), .A(n464), .ZN(N400) );
  NOR4_X1 U542 ( .A1(n1338), .A2(n1339), .A3(n1340), .A4(n1341), .ZN(n1328) );
  NOR4_X1 U543 ( .A1(n1330), .A2(n1331), .A3(n1332), .A4(n1333), .ZN(n1329) );
  OAI221_X1 U544 ( .B1(n1971), .B2(n15), .C1(n1939), .C2(n12), .A(n1345), .ZN(
        n1338) );
  AOI21_X1 U545 ( .B1(n1310), .B2(n1311), .A(n464), .ZN(N401) );
  NOR4_X1 U546 ( .A1(n1320), .A2(n1321), .A3(n1322), .A4(n1323), .ZN(n1310) );
  NOR4_X1 U547 ( .A1(n1312), .A2(n1313), .A3(n1314), .A4(n1315), .ZN(n1311) );
  OAI221_X1 U548 ( .B1(n1970), .B2(n15), .C1(n1938), .C2(n12), .A(n1327), .ZN(
        n1320) );
  AOI21_X1 U549 ( .B1(n1292), .B2(n1293), .A(n464), .ZN(N402) );
  NOR4_X1 U550 ( .A1(n1302), .A2(n1303), .A3(n1304), .A4(n1305), .ZN(n1292) );
  NOR4_X1 U551 ( .A1(n1294), .A2(n1295), .A3(n1296), .A4(n1297), .ZN(n1293) );
  OAI221_X1 U552 ( .B1(n1969), .B2(n15), .C1(n1937), .C2(n12), .A(n1309), .ZN(
        n1302) );
  AOI21_X1 U553 ( .B1(n1274), .B2(n1275), .A(n464), .ZN(N403) );
  NOR4_X1 U554 ( .A1(n1284), .A2(n1285), .A3(n1286), .A4(n1287), .ZN(n1274) );
  NOR4_X1 U555 ( .A1(n1276), .A2(n1277), .A3(n1278), .A4(n1279), .ZN(n1275) );
  OAI221_X1 U556 ( .B1(n1968), .B2(n15), .C1(n1936), .C2(n12), .A(n1291), .ZN(
        n1284) );
  AOI21_X1 U557 ( .B1(n1256), .B2(n1257), .A(n464), .ZN(N404) );
  NOR4_X1 U558 ( .A1(n1266), .A2(n1267), .A3(n1268), .A4(n1269), .ZN(n1256) );
  NOR4_X1 U559 ( .A1(n1258), .A2(n1259), .A3(n1260), .A4(n1261), .ZN(n1257) );
  OAI221_X1 U560 ( .B1(n1967), .B2(n15), .C1(n1935), .C2(n12), .A(n1273), .ZN(
        n1266) );
  AOI21_X1 U561 ( .B1(n1238), .B2(n1239), .A(n464), .ZN(N405) );
  NOR4_X1 U562 ( .A1(n1248), .A2(n1249), .A3(n1250), .A4(n1251), .ZN(n1238) );
  NOR4_X1 U563 ( .A1(n1240), .A2(n1241), .A3(n1242), .A4(n1243), .ZN(n1239) );
  OAI221_X1 U564 ( .B1(n1966), .B2(n15), .C1(n1934), .C2(n12), .A(n1255), .ZN(
        n1248) );
  AOI21_X1 U565 ( .B1(n1220), .B2(n1221), .A(n464), .ZN(N406) );
  NOR4_X1 U566 ( .A1(n1230), .A2(n1231), .A3(n1232), .A4(n1233), .ZN(n1220) );
  NOR4_X1 U567 ( .A1(n1222), .A2(n1223), .A3(n1224), .A4(n1225), .ZN(n1221) );
  OAI221_X1 U568 ( .B1(n1965), .B2(n15), .C1(n1933), .C2(n12), .A(n1237), .ZN(
        n1230) );
  AOI21_X1 U569 ( .B1(n1202), .B2(n1203), .A(n464), .ZN(N407) );
  NOR4_X1 U570 ( .A1(n1212), .A2(n1213), .A3(n1214), .A4(n1215), .ZN(n1202) );
  NOR4_X1 U571 ( .A1(n1204), .A2(n1205), .A3(n1206), .A4(n1207), .ZN(n1203) );
  OAI221_X1 U572 ( .B1(n1964), .B2(n15), .C1(n1932), .C2(n12), .A(n1219), .ZN(
        n1212) );
  AOI21_X1 U573 ( .B1(n1152), .B2(n1153), .A(n464), .ZN(N408) );
  NOR4_X1 U574 ( .A1(n1178), .A2(n1179), .A3(n1180), .A4(n1181), .ZN(n1152) );
  NOR4_X1 U575 ( .A1(n1154), .A2(n1155), .A3(n1156), .A4(n1157), .ZN(n1153) );
  OAI221_X1 U576 ( .B1(n1963), .B2(n15), .C1(n1931), .C2(n12), .A(n1199), .ZN(
        n1178) );
  AOI21_X1 U577 ( .B1(n1099), .B2(n1100), .A(n464), .ZN(N411) );
  NOR4_X1 U578 ( .A1(n1109), .A2(n1110), .A3(n1111), .A4(n1112), .ZN(n1099) );
  NOR4_X1 U579 ( .A1(n1101), .A2(n1102), .A3(n1103), .A4(n1104), .ZN(n1100) );
  OAI221_X1 U580 ( .B1(n109), .B2(n1993), .C1(n106), .C2(n1961), .A(n1116), 
        .ZN(n1109) );
  AOI21_X1 U581 ( .B1(n1081), .B2(n1082), .A(n462), .ZN(N412) );
  NOR4_X1 U582 ( .A1(n1091), .A2(n1092), .A3(n1093), .A4(n1094), .ZN(n1081) );
  NOR4_X1 U583 ( .A1(n1083), .A2(n1084), .A3(n1085), .A4(n1086), .ZN(n1082) );
  OAI221_X1 U584 ( .B1(n109), .B2(n1992), .C1(n106), .C2(n1960), .A(n1098), 
        .ZN(n1091) );
  AOI21_X1 U585 ( .B1(n1063), .B2(n1064), .A(n463), .ZN(N413) );
  NOR4_X1 U586 ( .A1(n1073), .A2(n1074), .A3(n1075), .A4(n1076), .ZN(n1063) );
  NOR4_X1 U587 ( .A1(n1065), .A2(n1066), .A3(n1067), .A4(n1068), .ZN(n1064) );
  OAI221_X1 U588 ( .B1(n109), .B2(n1991), .C1(n106), .C2(n1959), .A(n1080), 
        .ZN(n1073) );
  AOI21_X1 U589 ( .B1(n1045), .B2(n1046), .A(n464), .ZN(N414) );
  NOR4_X1 U590 ( .A1(n1055), .A2(n1056), .A3(n1057), .A4(n1058), .ZN(n1045) );
  NOR4_X1 U591 ( .A1(n1047), .A2(n1048), .A3(n1049), .A4(n1050), .ZN(n1046) );
  OAI221_X1 U592 ( .B1(n109), .B2(n1990), .C1(n106), .C2(n1958), .A(n1062), 
        .ZN(n1055) );
  AOI21_X1 U593 ( .B1(n1027), .B2(n1028), .A(n462), .ZN(N415) );
  NOR4_X1 U594 ( .A1(n1037), .A2(n1038), .A3(n1039), .A4(n1040), .ZN(n1027) );
  NOR4_X1 U595 ( .A1(n1029), .A2(n1030), .A3(n1031), .A4(n1032), .ZN(n1028) );
  OAI221_X1 U596 ( .B1(n109), .B2(n1989), .C1(n106), .C2(n1957), .A(n1044), 
        .ZN(n1037) );
  AOI21_X1 U597 ( .B1(n1009), .B2(n1010), .A(n463), .ZN(N416) );
  NOR4_X1 U598 ( .A1(n1019), .A2(n1020), .A3(n1021), .A4(n1022), .ZN(n1009) );
  NOR4_X1 U599 ( .A1(n1011), .A2(n1012), .A3(n1013), .A4(n1014), .ZN(n1010) );
  OAI221_X1 U600 ( .B1(n109), .B2(n1988), .C1(n106), .C2(n1956), .A(n1026), 
        .ZN(n1019) );
  AOI21_X1 U601 ( .B1(n991), .B2(n992), .A(n464), .ZN(N417) );
  NOR4_X1 U602 ( .A1(n1001), .A2(n1002), .A3(n1003), .A4(n1004), .ZN(n991) );
  NOR4_X1 U603 ( .A1(n993), .A2(n994), .A3(n995), .A4(n996), .ZN(n992) );
  OAI221_X1 U604 ( .B1(n109), .B2(n1987), .C1(n106), .C2(n1955), .A(n1008), 
        .ZN(n1001) );
  AOI21_X1 U605 ( .B1(n973), .B2(n974), .A(n462), .ZN(N418) );
  NOR4_X1 U606 ( .A1(n983), .A2(n984), .A3(n985), .A4(n986), .ZN(n973) );
  NOR4_X1 U607 ( .A1(n975), .A2(n976), .A3(n977), .A4(n978), .ZN(n974) );
  OAI221_X1 U608 ( .B1(n109), .B2(n1986), .C1(n106), .C2(n1954), .A(n990), 
        .ZN(n983) );
  AOI21_X1 U609 ( .B1(n955), .B2(n956), .A(n463), .ZN(N419) );
  NOR4_X1 U610 ( .A1(n965), .A2(n966), .A3(n967), .A4(n968), .ZN(n955) );
  NOR4_X1 U611 ( .A1(n957), .A2(n958), .A3(n959), .A4(n960), .ZN(n956) );
  OAI221_X1 U612 ( .B1(n109), .B2(n1985), .C1(n106), .C2(n1953), .A(n972), 
        .ZN(n965) );
  AOI21_X1 U613 ( .B1(n937), .B2(n938), .A(n464), .ZN(N420) );
  NOR4_X1 U614 ( .A1(n947), .A2(n948), .A3(n949), .A4(n950), .ZN(n937) );
  NOR4_X1 U615 ( .A1(n939), .A2(n940), .A3(n941), .A4(n942), .ZN(n938) );
  OAI221_X1 U616 ( .B1(n109), .B2(n1984), .C1(n106), .C2(n1952), .A(n954), 
        .ZN(n947) );
  AOI21_X1 U617 ( .B1(n919), .B2(n920), .A(n462), .ZN(N421) );
  NOR4_X1 U618 ( .A1(n929), .A2(n930), .A3(n931), .A4(n932), .ZN(n919) );
  NOR4_X1 U619 ( .A1(n921), .A2(n922), .A3(n923), .A4(n924), .ZN(n920) );
  OAI221_X1 U620 ( .B1(n109), .B2(n1983), .C1(n107), .C2(n1951), .A(n936), 
        .ZN(n929) );
  AOI21_X1 U621 ( .B1(n901), .B2(n902), .A(n463), .ZN(N422) );
  NOR4_X1 U622 ( .A1(n911), .A2(n912), .A3(n913), .A4(n914), .ZN(n901) );
  NOR4_X1 U623 ( .A1(n903), .A2(n904), .A3(n905), .A4(n906), .ZN(n902) );
  OAI221_X1 U624 ( .B1(n110), .B2(n1982), .C1(n107), .C2(n1950), .A(n918), 
        .ZN(n911) );
  AOI21_X1 U625 ( .B1(n883), .B2(n884), .A(n464), .ZN(N423) );
  NOR4_X1 U626 ( .A1(n893), .A2(n894), .A3(n895), .A4(n896), .ZN(n883) );
  NOR4_X1 U627 ( .A1(n885), .A2(n886), .A3(n887), .A4(n888), .ZN(n884) );
  OAI221_X1 U628 ( .B1(n110), .B2(n1981), .C1(n107), .C2(n1949), .A(n900), 
        .ZN(n893) );
  AOI21_X1 U629 ( .B1(n865), .B2(n866), .A(n462), .ZN(N424) );
  NOR4_X1 U630 ( .A1(n875), .A2(n876), .A3(n877), .A4(n878), .ZN(n865) );
  NOR4_X1 U631 ( .A1(n867), .A2(n868), .A3(n869), .A4(n870), .ZN(n866) );
  OAI221_X1 U632 ( .B1(n110), .B2(n1980), .C1(n107), .C2(n1948), .A(n882), 
        .ZN(n875) );
  AOI21_X1 U633 ( .B1(n847), .B2(n848), .A(n462), .ZN(N425) );
  NOR4_X1 U634 ( .A1(n857), .A2(n858), .A3(n859), .A4(n860), .ZN(n847) );
  NOR4_X1 U635 ( .A1(n849), .A2(n850), .A3(n851), .A4(n852), .ZN(n848) );
  OAI221_X1 U636 ( .B1(n110), .B2(n1979), .C1(n107), .C2(n1947), .A(n864), 
        .ZN(n857) );
  AOI21_X1 U637 ( .B1(n829), .B2(n830), .A(n463), .ZN(N426) );
  NOR4_X1 U638 ( .A1(n839), .A2(n840), .A3(n841), .A4(n842), .ZN(n829) );
  NOR4_X1 U639 ( .A1(n831), .A2(n832), .A3(n833), .A4(n834), .ZN(n830) );
  OAI221_X1 U640 ( .B1(n110), .B2(n1978), .C1(n107), .C2(n1946), .A(n846), 
        .ZN(n839) );
  AOI21_X1 U641 ( .B1(n811), .B2(n812), .A(n464), .ZN(N427) );
  NOR4_X1 U642 ( .A1(n821), .A2(n822), .A3(n823), .A4(n824), .ZN(n811) );
  NOR4_X1 U643 ( .A1(n813), .A2(n814), .A3(n815), .A4(n816), .ZN(n812) );
  OAI221_X1 U644 ( .B1(n110), .B2(n1977), .C1(n107), .C2(n1945), .A(n828), 
        .ZN(n821) );
  AOI21_X1 U645 ( .B1(n793), .B2(n794), .A(n463), .ZN(N428) );
  NOR4_X1 U646 ( .A1(n803), .A2(n804), .A3(n805), .A4(n806), .ZN(n793) );
  NOR4_X1 U647 ( .A1(n795), .A2(n796), .A3(n797), .A4(n798), .ZN(n794) );
  OAI221_X1 U648 ( .B1(n110), .B2(n1976), .C1(n107), .C2(n1944), .A(n810), 
        .ZN(n803) );
  AOI21_X1 U649 ( .B1(n775), .B2(n776), .A(n462), .ZN(N429) );
  NOR4_X1 U650 ( .A1(n785), .A2(n786), .A3(n787), .A4(n788), .ZN(n775) );
  NOR4_X1 U651 ( .A1(n777), .A2(n778), .A3(n779), .A4(n780), .ZN(n776) );
  OAI221_X1 U652 ( .B1(n110), .B2(n1975), .C1(n107), .C2(n1943), .A(n792), 
        .ZN(n785) );
  AOI21_X1 U653 ( .B1(n757), .B2(n758), .A(n463), .ZN(N430) );
  NOR4_X1 U654 ( .A1(n767), .A2(n768), .A3(n769), .A4(n770), .ZN(n757) );
  NOR4_X1 U655 ( .A1(n759), .A2(n760), .A3(n761), .A4(n762), .ZN(n758) );
  OAI221_X1 U656 ( .B1(n110), .B2(n1974), .C1(n107), .C2(n1942), .A(n774), 
        .ZN(n767) );
  AOI21_X1 U657 ( .B1(n739), .B2(n740), .A(n464), .ZN(N431) );
  NOR4_X1 U658 ( .A1(n749), .A2(n750), .A3(n751), .A4(n752), .ZN(n739) );
  NOR4_X1 U659 ( .A1(n741), .A2(n742), .A3(n743), .A4(n744), .ZN(n740) );
  OAI221_X1 U660 ( .B1(n110), .B2(n1973), .C1(n107), .C2(n1941), .A(n756), 
        .ZN(n749) );
  AOI21_X1 U661 ( .B1(n721), .B2(n722), .A(n464), .ZN(N432) );
  NOR4_X1 U662 ( .A1(n731), .A2(n732), .A3(n733), .A4(n734), .ZN(n721) );
  NOR4_X1 U663 ( .A1(n723), .A2(n724), .A3(n725), .A4(n726), .ZN(n722) );
  OAI221_X1 U664 ( .B1(n110), .B2(n1972), .C1(n108), .C2(n1940), .A(n738), 
        .ZN(n731) );
  AOI21_X1 U665 ( .B1(n703), .B2(n704), .A(n462), .ZN(N433) );
  NOR4_X1 U666 ( .A1(n713), .A2(n714), .A3(n715), .A4(n716), .ZN(n703) );
  NOR4_X1 U667 ( .A1(n705), .A2(n706), .A3(n707), .A4(n708), .ZN(n704) );
  OAI221_X1 U668 ( .B1(n110), .B2(n1971), .C1(n108), .C2(n1939), .A(n720), 
        .ZN(n713) );
  AOI21_X1 U669 ( .B1(n685), .B2(n686), .A(n463), .ZN(N434) );
  NOR4_X1 U670 ( .A1(n695), .A2(n696), .A3(n697), .A4(n698), .ZN(n685) );
  NOR4_X1 U671 ( .A1(n687), .A2(n688), .A3(n689), .A4(n690), .ZN(n686) );
  OAI221_X1 U672 ( .B1(n111), .B2(n1970), .C1(n108), .C2(n1938), .A(n702), 
        .ZN(n695) );
  AOI21_X1 U673 ( .B1(n667), .B2(n668), .A(n464), .ZN(N435) );
  NOR4_X1 U674 ( .A1(n677), .A2(n678), .A3(n679), .A4(n680), .ZN(n667) );
  NOR4_X1 U675 ( .A1(n669), .A2(n670), .A3(n671), .A4(n672), .ZN(n668) );
  OAI221_X1 U676 ( .B1(n111), .B2(n1969), .C1(n108), .C2(n1937), .A(n684), 
        .ZN(n677) );
  AOI21_X1 U677 ( .B1(n649), .B2(n650), .A(n462), .ZN(N436) );
  NOR4_X1 U678 ( .A1(n659), .A2(n660), .A3(n661), .A4(n662), .ZN(n649) );
  NOR4_X1 U679 ( .A1(n651), .A2(n652), .A3(n653), .A4(n654), .ZN(n650) );
  OAI221_X1 U680 ( .B1(n111), .B2(n1968), .C1(n108), .C2(n1936), .A(n666), 
        .ZN(n659) );
  AOI21_X1 U681 ( .B1(n631), .B2(n632), .A(n462), .ZN(N437) );
  NOR4_X1 U682 ( .A1(n641), .A2(n642), .A3(n643), .A4(n644), .ZN(n631) );
  NOR4_X1 U683 ( .A1(n633), .A2(n634), .A3(n635), .A4(n636), .ZN(n632) );
  OAI221_X1 U684 ( .B1(n111), .B2(n1967), .C1(n108), .C2(n1935), .A(n648), 
        .ZN(n641) );
  AOI21_X1 U685 ( .B1(n613), .B2(n614), .A(n462), .ZN(N438) );
  NOR4_X1 U686 ( .A1(n623), .A2(n624), .A3(n625), .A4(n626), .ZN(n613) );
  NOR4_X1 U687 ( .A1(n615), .A2(n616), .A3(n617), .A4(n618), .ZN(n614) );
  OAI221_X1 U688 ( .B1(n111), .B2(n1966), .C1(n108), .C2(n1934), .A(n630), 
        .ZN(n623) );
  AOI21_X1 U689 ( .B1(n595), .B2(n596), .A(n463), .ZN(N439) );
  NOR4_X1 U690 ( .A1(n605), .A2(n606), .A3(n607), .A4(n608), .ZN(n595) );
  NOR4_X1 U691 ( .A1(n597), .A2(n598), .A3(n599), .A4(n600), .ZN(n596) );
  OAI221_X1 U692 ( .B1(n111), .B2(n1965), .C1(n108), .C2(n1933), .A(n612), 
        .ZN(n605) );
  AOI21_X1 U693 ( .B1(n577), .B2(n578), .A(n464), .ZN(N440) );
  NOR4_X1 U694 ( .A1(n587), .A2(n588), .A3(n589), .A4(n590), .ZN(n577) );
  NOR4_X1 U695 ( .A1(n579), .A2(n580), .A3(n581), .A4(n582), .ZN(n578) );
  OAI221_X1 U696 ( .B1(n111), .B2(n1964), .C1(n108), .C2(n1932), .A(n594), 
        .ZN(n587) );
  AOI21_X1 U697 ( .B1(n527), .B2(n528), .A(n463), .ZN(N441) );
  NOR4_X1 U698 ( .A1(n553), .A2(n554), .A3(n555), .A4(n556), .ZN(n527) );
  NOR4_X1 U699 ( .A1(n529), .A2(n530), .A3(n531), .A4(n532), .ZN(n528) );
  OAI221_X1 U700 ( .B1(n111), .B2(n1963), .C1(n108), .C2(n1931), .A(n574), 
        .ZN(n553) );
  AND2_X1 U701 ( .A1(DATAIN[10]), .A2(n2), .ZN(N323) );
  AND2_X1 U702 ( .A1(DATAIN[11]), .A2(n2), .ZN(N324) );
  AND2_X1 U703 ( .A1(DATAIN[12]), .A2(n2), .ZN(N325) );
  AND2_X1 U704 ( .A1(DATAIN[13]), .A2(n2), .ZN(N326) );
  AND2_X1 U705 ( .A1(DATAIN[14]), .A2(n2), .ZN(N327) );
  AND2_X1 U706 ( .A1(DATAIN[15]), .A2(n2), .ZN(N328) );
  AND2_X1 U707 ( .A1(DATAIN[16]), .A2(n2), .ZN(N329) );
  AND2_X1 U708 ( .A1(DATAIN[17]), .A2(n2), .ZN(N330) );
  AND2_X1 U709 ( .A1(DATAIN[18]), .A2(n2), .ZN(N331) );
  AND2_X1 U710 ( .A1(DATAIN[19]), .A2(n2), .ZN(N332) );
  AND2_X1 U711 ( .A1(DATAIN[20]), .A2(n2), .ZN(N333) );
  AND2_X1 U712 ( .A1(DATAIN[21]), .A2(n1), .ZN(N334) );
  AND2_X1 U713 ( .A1(DATAIN[22]), .A2(n1), .ZN(N335) );
  AND2_X1 U714 ( .A1(DATAIN[23]), .A2(n1), .ZN(N336) );
  AND2_X1 U715 ( .A1(DATAIN[24]), .A2(n1), .ZN(N337) );
  AND2_X1 U716 ( .A1(DATAIN[25]), .A2(n1), .ZN(N338) );
  AND2_X1 U717 ( .A1(DATAIN[26]), .A2(n1), .ZN(N339) );
  AND2_X1 U718 ( .A1(DATAIN[27]), .A2(n1), .ZN(N340) );
  AND2_X1 U719 ( .A1(DATAIN[28]), .A2(n1), .ZN(N341) );
  AND2_X1 U720 ( .A1(DATAIN[29]), .A2(n1), .ZN(N342) );
  AND2_X1 U721 ( .A1(DATAIN[30]), .A2(n1), .ZN(N343) );
  AND2_X1 U722 ( .A1(DATAIN[31]), .A2(n1), .ZN(N344) );
  AND2_X1 U723 ( .A1(DATAIN[0]), .A2(n3), .ZN(N313) );
  AND2_X1 U724 ( .A1(DATAIN[1]), .A2(n3), .ZN(N314) );
  AND2_X1 U725 ( .A1(DATAIN[2]), .A2(n3), .ZN(N315) );
  AND2_X1 U726 ( .A1(DATAIN[3]), .A2(n3), .ZN(N316) );
  AND2_X1 U727 ( .A1(DATAIN[4]), .A2(n3), .ZN(N317) );
  AND2_X1 U728 ( .A1(DATAIN[5]), .A2(n3), .ZN(N318) );
  AND2_X1 U729 ( .A1(DATAIN[6]), .A2(n3), .ZN(N319) );
  AND2_X1 U730 ( .A1(DATAIN[7]), .A2(n3), .ZN(N320) );
  AND2_X1 U731 ( .A1(DATAIN[8]), .A2(n3), .ZN(N321) );
  AND2_X1 U732 ( .A1(DATAIN[9]), .A2(n3), .ZN(N322) );
  NAND2_X1 U733 ( .A1(n473), .A2(n1777), .ZN(N375) );
  AND2_X1 U734 ( .A1(n474), .A2(n1777), .ZN(n1790) );
  OAI221_X1 U735 ( .B1(n195), .B2(n2034), .C1(n192), .C2(n2002), .A(n691), 
        .ZN(n690) );
  AOI22_X1 U736 ( .A1(\REGISTERS[19][24] ), .A2(n189), .B1(\REGISTERS[18][24] ), .B2(n186), .ZN(n691) );
  OAI221_X1 U737 ( .B1(n147), .B2(n514), .C1(n144), .C2(n482), .A(n699), .ZN(
        n698) );
  AOI22_X1 U738 ( .A1(\REGISTERS[3][24] ), .A2(n141), .B1(\REGISTERS[2][24] ), 
        .B2(n138), .ZN(n699) );
  OAI221_X1 U739 ( .B1(n195), .B2(n2033), .C1(n192), .C2(n2001), .A(n673), 
        .ZN(n672) );
  AOI22_X1 U740 ( .A1(\REGISTERS[19][25] ), .A2(n189), .B1(\REGISTERS[18][25] ), .B2(n186), .ZN(n673) );
  OAI221_X1 U741 ( .B1(n147), .B2(n513), .C1(n144), .C2(n481), .A(n681), .ZN(
        n680) );
  AOI22_X1 U742 ( .A1(\REGISTERS[3][25] ), .A2(n141), .B1(\REGISTERS[2][25] ), 
        .B2(n138), .ZN(n681) );
  OAI221_X1 U743 ( .B1(n195), .B2(n2032), .C1(n192), .C2(n2000), .A(n655), 
        .ZN(n654) );
  AOI22_X1 U744 ( .A1(\REGISTERS[19][26] ), .A2(n189), .B1(\REGISTERS[18][26] ), .B2(n186), .ZN(n655) );
  OAI221_X1 U745 ( .B1(n147), .B2(n512), .C1(n144), .C2(n480), .A(n663), .ZN(
        n662) );
  AOI22_X1 U746 ( .A1(\REGISTERS[3][26] ), .A2(n141), .B1(\REGISTERS[2][26] ), 
        .B2(n138), .ZN(n663) );
  OAI221_X1 U747 ( .B1(n195), .B2(n2031), .C1(n192), .C2(n1999), .A(n637), 
        .ZN(n636) );
  AOI22_X1 U748 ( .A1(\REGISTERS[19][27] ), .A2(n189), .B1(\REGISTERS[18][27] ), .B2(n186), .ZN(n637) );
  OAI221_X1 U749 ( .B1(n147), .B2(n511), .C1(n144), .C2(n479), .A(n645), .ZN(
        n644) );
  AOI22_X1 U750 ( .A1(\REGISTERS[3][27] ), .A2(n141), .B1(\REGISTERS[2][27] ), 
        .B2(n138), .ZN(n645) );
  OAI221_X1 U751 ( .B1(n195), .B2(n2030), .C1(n192), .C2(n1998), .A(n619), 
        .ZN(n618) );
  AOI22_X1 U752 ( .A1(\REGISTERS[19][28] ), .A2(n189), .B1(\REGISTERS[18][28] ), .B2(n186), .ZN(n619) );
  OAI221_X1 U753 ( .B1(n147), .B2(n510), .C1(n144), .C2(n478), .A(n627), .ZN(
        n626) );
  AOI22_X1 U754 ( .A1(\REGISTERS[3][28] ), .A2(n141), .B1(\REGISTERS[2][28] ), 
        .B2(n138), .ZN(n627) );
  OAI221_X1 U755 ( .B1(n195), .B2(n2029), .C1(n192), .C2(n1997), .A(n601), 
        .ZN(n600) );
  AOI22_X1 U756 ( .A1(\REGISTERS[19][29] ), .A2(n189), .B1(\REGISTERS[18][29] ), .B2(n186), .ZN(n601) );
  OAI221_X1 U757 ( .B1(n147), .B2(n509), .C1(n144), .C2(n477), .A(n609), .ZN(
        n608) );
  AOI22_X1 U758 ( .A1(\REGISTERS[3][29] ), .A2(n141), .B1(\REGISTERS[2][29] ), 
        .B2(n138), .ZN(n609) );
  OAI221_X1 U759 ( .B1(n195), .B2(n2028), .C1(n192), .C2(n1996), .A(n583), 
        .ZN(n582) );
  AOI22_X1 U760 ( .A1(\REGISTERS[19][30] ), .A2(n189), .B1(\REGISTERS[18][30] ), .B2(n186), .ZN(n583) );
  OAI221_X1 U761 ( .B1(n147), .B2(n508), .C1(n144), .C2(n476), .A(n591), .ZN(
        n590) );
  AOI22_X1 U762 ( .A1(\REGISTERS[3][30] ), .A2(n141), .B1(\REGISTERS[2][30] ), 
        .B2(n138), .ZN(n591) );
  OAI221_X1 U763 ( .B1(n195), .B2(n2027), .C1(n192), .C2(n1995), .A(n535), 
        .ZN(n532) );
  AOI22_X1 U764 ( .A1(\REGISTERS[19][31] ), .A2(n189), .B1(\REGISTERS[18][31] ), .B2(n186), .ZN(n535) );
  OAI221_X1 U765 ( .B1(n147), .B2(n507), .C1(n144), .C2(n475), .A(n559), .ZN(
        n556) );
  AOI22_X1 U766 ( .A1(\REGISTERS[3][31] ), .A2(n141), .B1(\REGISTERS[2][31] ), 
        .B2(n138), .ZN(n559) );
  OAI221_X1 U767 ( .B1(n2058), .B2(n97), .C1(n2026), .C2(n94), .A(n1748), .ZN(
        n1747) );
  AOI22_X1 U768 ( .A1(n91), .A2(\REGISTERS[19][0] ), .B1(n88), .B2(
        \REGISTERS[18][0] ), .ZN(n1748) );
  OAI221_X1 U769 ( .B1(n1802), .B2(n49), .C1(n506), .C2(n46), .A(n1766), .ZN(
        n1765) );
  AOI22_X1 U770 ( .A1(n43), .A2(\REGISTERS[3][0] ), .B1(n40), .B2(
        \REGISTERS[2][0] ), .ZN(n1766) );
  OAI221_X1 U771 ( .B1(n2057), .B2(n97), .C1(n2025), .C2(n94), .A(n1730), .ZN(
        n1729) );
  AOI22_X1 U772 ( .A1(n91), .A2(\REGISTERS[19][1] ), .B1(n88), .B2(
        \REGISTERS[18][1] ), .ZN(n1730) );
  OAI221_X1 U773 ( .B1(n1801), .B2(n49), .C1(n505), .C2(n46), .A(n1738), .ZN(
        n1737) );
  AOI22_X1 U774 ( .A1(n43), .A2(\REGISTERS[3][1] ), .B1(n40), .B2(
        \REGISTERS[2][1] ), .ZN(n1738) );
  OAI221_X1 U775 ( .B1(n2056), .B2(n97), .C1(n2024), .C2(n94), .A(n1712), .ZN(
        n1711) );
  AOI22_X1 U776 ( .A1(n91), .A2(\REGISTERS[19][2] ), .B1(n88), .B2(
        \REGISTERS[18][2] ), .ZN(n1712) );
  OAI221_X1 U777 ( .B1(n1800), .B2(n49), .C1(n504), .C2(n46), .A(n1720), .ZN(
        n1719) );
  AOI22_X1 U778 ( .A1(n43), .A2(\REGISTERS[3][2] ), .B1(n40), .B2(
        \REGISTERS[2][2] ), .ZN(n1720) );
  OAI221_X1 U779 ( .B1(n2055), .B2(n97), .C1(n2023), .C2(n94), .A(n1694), .ZN(
        n1693) );
  AOI22_X1 U780 ( .A1(n91), .A2(\REGISTERS[19][3] ), .B1(n88), .B2(
        \REGISTERS[18][3] ), .ZN(n1694) );
  OAI221_X1 U781 ( .B1(n1799), .B2(n49), .C1(n503), .C2(n46), .A(n1702), .ZN(
        n1701) );
  AOI22_X1 U782 ( .A1(n43), .A2(\REGISTERS[3][3] ), .B1(n40), .B2(
        \REGISTERS[2][3] ), .ZN(n1702) );
  OAI221_X1 U783 ( .B1(n2054), .B2(n97), .C1(n2022), .C2(n94), .A(n1676), .ZN(
        n1675) );
  AOI22_X1 U784 ( .A1(n91), .A2(\REGISTERS[19][4] ), .B1(n88), .B2(
        \REGISTERS[18][4] ), .ZN(n1676) );
  OAI221_X1 U785 ( .B1(n1798), .B2(n49), .C1(n502), .C2(n46), .A(n1684), .ZN(
        n1683) );
  AOI22_X1 U786 ( .A1(n43), .A2(\REGISTERS[3][4] ), .B1(n40), .B2(
        \REGISTERS[2][4] ), .ZN(n1684) );
  OAI221_X1 U787 ( .B1(n2053), .B2(n97), .C1(n2021), .C2(n94), .A(n1658), .ZN(
        n1657) );
  AOI22_X1 U788 ( .A1(n91), .A2(\REGISTERS[19][5] ), .B1(n88), .B2(
        \REGISTERS[18][5] ), .ZN(n1658) );
  OAI221_X1 U789 ( .B1(n1797), .B2(n49), .C1(n501), .C2(n46), .A(n1666), .ZN(
        n1665) );
  AOI22_X1 U790 ( .A1(n43), .A2(\REGISTERS[3][5] ), .B1(n40), .B2(
        \REGISTERS[2][5] ), .ZN(n1666) );
  OAI221_X1 U791 ( .B1(n2052), .B2(n97), .C1(n2020), .C2(n94), .A(n1640), .ZN(
        n1639) );
  AOI22_X1 U792 ( .A1(n91), .A2(\REGISTERS[19][6] ), .B1(n88), .B2(
        \REGISTERS[18][6] ), .ZN(n1640) );
  OAI221_X1 U793 ( .B1(n1796), .B2(n49), .C1(n500), .C2(n46), .A(n1648), .ZN(
        n1647) );
  AOI22_X1 U794 ( .A1(n43), .A2(\REGISTERS[3][6] ), .B1(n40), .B2(
        \REGISTERS[2][6] ), .ZN(n1648) );
  OAI221_X1 U795 ( .B1(n2051), .B2(n97), .C1(n2019), .C2(n94), .A(n1622), .ZN(
        n1621) );
  AOI22_X1 U796 ( .A1(n91), .A2(\REGISTERS[19][7] ), .B1(n88), .B2(
        \REGISTERS[18][7] ), .ZN(n1622) );
  OAI221_X1 U797 ( .B1(n1795), .B2(n49), .C1(n499), .C2(n46), .A(n1630), .ZN(
        n1629) );
  AOI22_X1 U798 ( .A1(n43), .A2(\REGISTERS[3][7] ), .B1(n40), .B2(
        \REGISTERS[2][7] ), .ZN(n1630) );
  OAI221_X1 U799 ( .B1(n2050), .B2(n97), .C1(n2018), .C2(n94), .A(n1604), .ZN(
        n1603) );
  AOI22_X1 U800 ( .A1(n91), .A2(\REGISTERS[19][8] ), .B1(n88), .B2(
        \REGISTERS[18][8] ), .ZN(n1604) );
  OAI221_X1 U801 ( .B1(n1794), .B2(n49), .C1(n498), .C2(n46), .A(n1612), .ZN(
        n1611) );
  AOI22_X1 U802 ( .A1(n43), .A2(\REGISTERS[3][8] ), .B1(n40), .B2(
        \REGISTERS[2][8] ), .ZN(n1612) );
  OAI221_X1 U803 ( .B1(n2049), .B2(n97), .C1(n2017), .C2(n94), .A(n1586), .ZN(
        n1585) );
  AOI22_X1 U804 ( .A1(n91), .A2(\REGISTERS[19][9] ), .B1(n88), .B2(
        \REGISTERS[18][9] ), .ZN(n1586) );
  OAI221_X1 U805 ( .B1(n1793), .B2(n49), .C1(n497), .C2(n46), .A(n1594), .ZN(
        n1593) );
  AOI22_X1 U806 ( .A1(n43), .A2(\REGISTERS[3][9] ), .B1(n40), .B2(
        \REGISTERS[2][9] ), .ZN(n1594) );
  OAI221_X1 U807 ( .B1(n2048), .B2(n97), .C1(n2016), .C2(n94), .A(n1568), .ZN(
        n1567) );
  AOI22_X1 U808 ( .A1(n91), .A2(\REGISTERS[19][10] ), .B1(n88), .B2(
        \REGISTERS[18][10] ), .ZN(n1568) );
  OAI221_X1 U809 ( .B1(n1792), .B2(n49), .C1(n496), .C2(n46), .A(n1576), .ZN(
        n1575) );
  AOI22_X1 U810 ( .A1(n43), .A2(\REGISTERS[3][10] ), .B1(n40), .B2(
        \REGISTERS[2][10] ), .ZN(n1576) );
  OAI221_X1 U811 ( .B1(n2036), .B2(n99), .C1(n2004), .C2(n96), .A(n1352), .ZN(
        n1351) );
  AOI22_X1 U812 ( .A1(n93), .A2(\REGISTERS[19][22] ), .B1(n90), .B2(
        \REGISTERS[18][22] ), .ZN(n1352) );
  OAI221_X1 U813 ( .B1(n516), .B2(n51), .C1(n484), .C2(n48), .A(n1360), .ZN(
        n1359) );
  AOI22_X1 U814 ( .A1(n45), .A2(\REGISTERS[3][22] ), .B1(n42), .B2(
        \REGISTERS[2][22] ), .ZN(n1360) );
  OAI221_X1 U815 ( .B1(n2035), .B2(n99), .C1(n2003), .C2(n96), .A(n1334), .ZN(
        n1333) );
  AOI22_X1 U816 ( .A1(n93), .A2(\REGISTERS[19][23] ), .B1(n90), .B2(
        \REGISTERS[18][23] ), .ZN(n1334) );
  OAI221_X1 U817 ( .B1(n515), .B2(n51), .C1(n483), .C2(n48), .A(n1342), .ZN(
        n1341) );
  AOI22_X1 U818 ( .A1(n45), .A2(\REGISTERS[3][23] ), .B1(n42), .B2(
        \REGISTERS[2][23] ), .ZN(n1342) );
  OAI221_X1 U819 ( .B1(n2034), .B2(n99), .C1(n2002), .C2(n96), .A(n1316), .ZN(
        n1315) );
  AOI22_X1 U820 ( .A1(n93), .A2(\REGISTERS[19][24] ), .B1(n90), .B2(
        \REGISTERS[18][24] ), .ZN(n1316) );
  OAI221_X1 U821 ( .B1(n514), .B2(n51), .C1(n482), .C2(n48), .A(n1324), .ZN(
        n1323) );
  AOI22_X1 U822 ( .A1(n45), .A2(\REGISTERS[3][24] ), .B1(n42), .B2(
        \REGISTERS[2][24] ), .ZN(n1324) );
  OAI221_X1 U823 ( .B1(n2033), .B2(n99), .C1(n2001), .C2(n96), .A(n1298), .ZN(
        n1297) );
  AOI22_X1 U824 ( .A1(n93), .A2(\REGISTERS[19][25] ), .B1(n90), .B2(
        \REGISTERS[18][25] ), .ZN(n1298) );
  OAI221_X1 U825 ( .B1(n513), .B2(n51), .C1(n481), .C2(n48), .A(n1306), .ZN(
        n1305) );
  AOI22_X1 U826 ( .A1(n45), .A2(\REGISTERS[3][25] ), .B1(n42), .B2(
        \REGISTERS[2][25] ), .ZN(n1306) );
  OAI221_X1 U827 ( .B1(n2032), .B2(n99), .C1(n2000), .C2(n96), .A(n1280), .ZN(
        n1279) );
  AOI22_X1 U828 ( .A1(n93), .A2(\REGISTERS[19][26] ), .B1(n90), .B2(
        \REGISTERS[18][26] ), .ZN(n1280) );
  OAI221_X1 U829 ( .B1(n512), .B2(n51), .C1(n480), .C2(n48), .A(n1288), .ZN(
        n1287) );
  AOI22_X1 U830 ( .A1(n45), .A2(\REGISTERS[3][26] ), .B1(n42), .B2(
        \REGISTERS[2][26] ), .ZN(n1288) );
  OAI221_X1 U831 ( .B1(n2031), .B2(n99), .C1(n1999), .C2(n96), .A(n1262), .ZN(
        n1261) );
  AOI22_X1 U832 ( .A1(n93), .A2(\REGISTERS[19][27] ), .B1(n90), .B2(
        \REGISTERS[18][27] ), .ZN(n1262) );
  OAI221_X1 U833 ( .B1(n511), .B2(n51), .C1(n479), .C2(n48), .A(n1270), .ZN(
        n1269) );
  AOI22_X1 U834 ( .A1(n45), .A2(\REGISTERS[3][27] ), .B1(n42), .B2(
        \REGISTERS[2][27] ), .ZN(n1270) );
  OAI221_X1 U835 ( .B1(n2030), .B2(n99), .C1(n1998), .C2(n96), .A(n1244), .ZN(
        n1243) );
  AOI22_X1 U836 ( .A1(n93), .A2(\REGISTERS[19][28] ), .B1(n90), .B2(
        \REGISTERS[18][28] ), .ZN(n1244) );
  OAI221_X1 U837 ( .B1(n510), .B2(n51), .C1(n478), .C2(n48), .A(n1252), .ZN(
        n1251) );
  AOI22_X1 U838 ( .A1(n45), .A2(\REGISTERS[3][28] ), .B1(n42), .B2(
        \REGISTERS[2][28] ), .ZN(n1252) );
  OAI221_X1 U839 ( .B1(n2029), .B2(n99), .C1(n1997), .C2(n96), .A(n1226), .ZN(
        n1225) );
  AOI22_X1 U840 ( .A1(n93), .A2(\REGISTERS[19][29] ), .B1(n90), .B2(
        \REGISTERS[18][29] ), .ZN(n1226) );
  OAI221_X1 U841 ( .B1(n509), .B2(n51), .C1(n477), .C2(n48), .A(n1234), .ZN(
        n1233) );
  AOI22_X1 U842 ( .A1(n45), .A2(\REGISTERS[3][29] ), .B1(n42), .B2(
        \REGISTERS[2][29] ), .ZN(n1234) );
  OAI221_X1 U843 ( .B1(n2028), .B2(n99), .C1(n1996), .C2(n96), .A(n1208), .ZN(
        n1207) );
  AOI22_X1 U844 ( .A1(n93), .A2(\REGISTERS[19][30] ), .B1(n90), .B2(
        \REGISTERS[18][30] ), .ZN(n1208) );
  OAI221_X1 U845 ( .B1(n508), .B2(n51), .C1(n476), .C2(n48), .A(n1216), .ZN(
        n1215) );
  AOI22_X1 U846 ( .A1(n45), .A2(\REGISTERS[3][30] ), .B1(n42), .B2(
        \REGISTERS[2][30] ), .ZN(n1216) );
  OAI221_X1 U847 ( .B1(n2027), .B2(n99), .C1(n1995), .C2(n96), .A(n1160), .ZN(
        n1157) );
  AOI22_X1 U848 ( .A1(n93), .A2(\REGISTERS[19][31] ), .B1(n90), .B2(
        \REGISTERS[18][31] ), .ZN(n1160) );
  OAI221_X1 U849 ( .B1(n507), .B2(n51), .C1(n475), .C2(n48), .A(n1184), .ZN(
        n1181) );
  AOI22_X1 U850 ( .A1(n45), .A2(\REGISTERS[3][31] ), .B1(n42), .B2(
        \REGISTERS[2][31] ), .ZN(n1184) );
  OAI221_X1 U851 ( .B1(n183), .B2(n2098), .C1(n180), .C2(n2066), .A(n692), 
        .ZN(n689) );
  AOI22_X1 U852 ( .A1(\REGISTERS[23][24] ), .A2(n177), .B1(\REGISTERS[22][24] ), .B2(n174), .ZN(n692) );
  OAI221_X1 U853 ( .B1(n135), .B2(n1842), .C1(n132), .C2(n1810), .A(n700), 
        .ZN(n697) );
  AOI22_X1 U854 ( .A1(\REGISTERS[7][24] ), .A2(n129), .B1(\REGISTERS[6][24] ), 
        .B2(n126), .ZN(n700) );
  OAI221_X1 U855 ( .B1(n183), .B2(n2097), .C1(n180), .C2(n2065), .A(n674), 
        .ZN(n671) );
  AOI22_X1 U856 ( .A1(\REGISTERS[23][25] ), .A2(n177), .B1(\REGISTERS[22][25] ), .B2(n174), .ZN(n674) );
  OAI221_X1 U857 ( .B1(n135), .B2(n1841), .C1(n132), .C2(n1809), .A(n682), 
        .ZN(n679) );
  AOI22_X1 U858 ( .A1(\REGISTERS[7][25] ), .A2(n129), .B1(\REGISTERS[6][25] ), 
        .B2(n126), .ZN(n682) );
  OAI221_X1 U859 ( .B1(n183), .B2(n2096), .C1(n180), .C2(n2064), .A(n656), 
        .ZN(n653) );
  AOI22_X1 U860 ( .A1(\REGISTERS[23][26] ), .A2(n177), .B1(\REGISTERS[22][26] ), .B2(n174), .ZN(n656) );
  OAI221_X1 U861 ( .B1(n135), .B2(n1840), .C1(n132), .C2(n1808), .A(n664), 
        .ZN(n661) );
  AOI22_X1 U862 ( .A1(\REGISTERS[7][26] ), .A2(n129), .B1(\REGISTERS[6][26] ), 
        .B2(n126), .ZN(n664) );
  OAI221_X1 U863 ( .B1(n183), .B2(n2095), .C1(n180), .C2(n2063), .A(n638), 
        .ZN(n635) );
  AOI22_X1 U864 ( .A1(\REGISTERS[23][27] ), .A2(n177), .B1(\REGISTERS[22][27] ), .B2(n174), .ZN(n638) );
  OAI221_X1 U865 ( .B1(n135), .B2(n1839), .C1(n132), .C2(n1807), .A(n646), 
        .ZN(n643) );
  AOI22_X1 U866 ( .A1(\REGISTERS[7][27] ), .A2(n129), .B1(\REGISTERS[6][27] ), 
        .B2(n126), .ZN(n646) );
  OAI221_X1 U867 ( .B1(n183), .B2(n2094), .C1(n180), .C2(n2062), .A(n620), 
        .ZN(n617) );
  AOI22_X1 U868 ( .A1(\REGISTERS[23][28] ), .A2(n177), .B1(\REGISTERS[22][28] ), .B2(n174), .ZN(n620) );
  OAI221_X1 U869 ( .B1(n135), .B2(n1838), .C1(n132), .C2(n1806), .A(n628), 
        .ZN(n625) );
  AOI22_X1 U870 ( .A1(\REGISTERS[7][28] ), .A2(n129), .B1(\REGISTERS[6][28] ), 
        .B2(n126), .ZN(n628) );
  OAI221_X1 U871 ( .B1(n183), .B2(n2093), .C1(n180), .C2(n2061), .A(n602), 
        .ZN(n599) );
  AOI22_X1 U872 ( .A1(\REGISTERS[23][29] ), .A2(n177), .B1(\REGISTERS[22][29] ), .B2(n174), .ZN(n602) );
  OAI221_X1 U873 ( .B1(n135), .B2(n1837), .C1(n132), .C2(n1805), .A(n610), 
        .ZN(n607) );
  AOI22_X1 U874 ( .A1(\REGISTERS[7][29] ), .A2(n129), .B1(\REGISTERS[6][29] ), 
        .B2(n126), .ZN(n610) );
  OAI221_X1 U875 ( .B1(n183), .B2(n2092), .C1(n180), .C2(n2060), .A(n584), 
        .ZN(n581) );
  AOI22_X1 U876 ( .A1(\REGISTERS[23][30] ), .A2(n177), .B1(\REGISTERS[22][30] ), .B2(n174), .ZN(n584) );
  OAI221_X1 U877 ( .B1(n135), .B2(n1836), .C1(n132), .C2(n1804), .A(n592), 
        .ZN(n589) );
  AOI22_X1 U878 ( .A1(\REGISTERS[7][30] ), .A2(n129), .B1(\REGISTERS[6][30] ), 
        .B2(n126), .ZN(n592) );
  OAI221_X1 U879 ( .B1(n183), .B2(n2091), .C1(n180), .C2(n2059), .A(n540), 
        .ZN(n531) );
  AOI22_X1 U880 ( .A1(\REGISTERS[23][31] ), .A2(n177), .B1(\REGISTERS[22][31] ), .B2(n174), .ZN(n540) );
  OAI221_X1 U881 ( .B1(n135), .B2(n1835), .C1(n132), .C2(n1803), .A(n564), 
        .ZN(n555) );
  AOI22_X1 U882 ( .A1(\REGISTERS[7][31] ), .A2(n129), .B1(\REGISTERS[6][31] ), 
        .B2(n126), .ZN(n564) );
  OAI221_X1 U883 ( .B1(n193), .B2(n2058), .C1(n190), .C2(n2026), .A(n1123), 
        .ZN(n1122) );
  AOI22_X1 U884 ( .A1(\REGISTERS[19][0] ), .A2(n187), .B1(\REGISTERS[18][0] ), 
        .B2(n184), .ZN(n1123) );
  OAI221_X1 U885 ( .B1(n145), .B2(n1802), .C1(n142), .C2(n506), .A(n1141), 
        .ZN(n1140) );
  AOI22_X1 U886 ( .A1(\REGISTERS[3][0] ), .A2(n139), .B1(\REGISTERS[2][0] ), 
        .B2(n136), .ZN(n1141) );
  OAI221_X1 U887 ( .B1(n193), .B2(n2057), .C1(n190), .C2(n2025), .A(n1105), 
        .ZN(n1104) );
  AOI22_X1 U888 ( .A1(\REGISTERS[19][1] ), .A2(n187), .B1(\REGISTERS[18][1] ), 
        .B2(n184), .ZN(n1105) );
  OAI221_X1 U889 ( .B1(n145), .B2(n1801), .C1(n142), .C2(n505), .A(n1113), 
        .ZN(n1112) );
  AOI22_X1 U890 ( .A1(\REGISTERS[3][1] ), .A2(n139), .B1(\REGISTERS[2][1] ), 
        .B2(n136), .ZN(n1113) );
  OAI221_X1 U891 ( .B1(n193), .B2(n2056), .C1(n190), .C2(n2024), .A(n1087), 
        .ZN(n1086) );
  AOI22_X1 U892 ( .A1(\REGISTERS[19][2] ), .A2(n187), .B1(\REGISTERS[18][2] ), 
        .B2(n184), .ZN(n1087) );
  OAI221_X1 U893 ( .B1(n145), .B2(n1800), .C1(n142), .C2(n504), .A(n1095), 
        .ZN(n1094) );
  AOI22_X1 U894 ( .A1(\REGISTERS[3][2] ), .A2(n139), .B1(\REGISTERS[2][2] ), 
        .B2(n136), .ZN(n1095) );
  OAI221_X1 U895 ( .B1(n193), .B2(n2055), .C1(n190), .C2(n2023), .A(n1069), 
        .ZN(n1068) );
  AOI22_X1 U896 ( .A1(\REGISTERS[19][3] ), .A2(n187), .B1(\REGISTERS[18][3] ), 
        .B2(n184), .ZN(n1069) );
  OAI221_X1 U897 ( .B1(n145), .B2(n1799), .C1(n142), .C2(n503), .A(n1077), 
        .ZN(n1076) );
  AOI22_X1 U898 ( .A1(\REGISTERS[3][3] ), .A2(n139), .B1(\REGISTERS[2][3] ), 
        .B2(n136), .ZN(n1077) );
  OAI221_X1 U899 ( .B1(n193), .B2(n2054), .C1(n190), .C2(n2022), .A(n1051), 
        .ZN(n1050) );
  AOI22_X1 U900 ( .A1(\REGISTERS[19][4] ), .A2(n187), .B1(\REGISTERS[18][4] ), 
        .B2(n184), .ZN(n1051) );
  OAI221_X1 U901 ( .B1(n145), .B2(n1798), .C1(n142), .C2(n502), .A(n1059), 
        .ZN(n1058) );
  AOI22_X1 U902 ( .A1(\REGISTERS[3][4] ), .A2(n139), .B1(\REGISTERS[2][4] ), 
        .B2(n136), .ZN(n1059) );
  OAI221_X1 U903 ( .B1(n193), .B2(n2053), .C1(n190), .C2(n2021), .A(n1033), 
        .ZN(n1032) );
  AOI22_X1 U904 ( .A1(\REGISTERS[19][5] ), .A2(n187), .B1(\REGISTERS[18][5] ), 
        .B2(n184), .ZN(n1033) );
  OAI221_X1 U905 ( .B1(n145), .B2(n1797), .C1(n142), .C2(n501), .A(n1041), 
        .ZN(n1040) );
  AOI22_X1 U906 ( .A1(\REGISTERS[3][5] ), .A2(n139), .B1(\REGISTERS[2][5] ), 
        .B2(n136), .ZN(n1041) );
  OAI221_X1 U907 ( .B1(n193), .B2(n2052), .C1(n190), .C2(n2020), .A(n1015), 
        .ZN(n1014) );
  AOI22_X1 U908 ( .A1(\REGISTERS[19][6] ), .A2(n187), .B1(\REGISTERS[18][6] ), 
        .B2(n184), .ZN(n1015) );
  OAI221_X1 U909 ( .B1(n145), .B2(n1796), .C1(n142), .C2(n500), .A(n1023), 
        .ZN(n1022) );
  AOI22_X1 U910 ( .A1(\REGISTERS[3][6] ), .A2(n139), .B1(\REGISTERS[2][6] ), 
        .B2(n136), .ZN(n1023) );
  OAI221_X1 U911 ( .B1(n193), .B2(n2051), .C1(n190), .C2(n2019), .A(n997), 
        .ZN(n996) );
  AOI22_X1 U912 ( .A1(\REGISTERS[19][7] ), .A2(n187), .B1(\REGISTERS[18][7] ), 
        .B2(n184), .ZN(n997) );
  OAI221_X1 U913 ( .B1(n145), .B2(n1795), .C1(n142), .C2(n499), .A(n1005), 
        .ZN(n1004) );
  AOI22_X1 U914 ( .A1(\REGISTERS[3][7] ), .A2(n139), .B1(\REGISTERS[2][7] ), 
        .B2(n136), .ZN(n1005) );
  OAI221_X1 U915 ( .B1(n193), .B2(n2050), .C1(n190), .C2(n2018), .A(n979), 
        .ZN(n978) );
  AOI22_X1 U916 ( .A1(\REGISTERS[19][8] ), .A2(n187), .B1(\REGISTERS[18][8] ), 
        .B2(n184), .ZN(n979) );
  OAI221_X1 U917 ( .B1(n145), .B2(n1794), .C1(n142), .C2(n498), .A(n987), .ZN(
        n986) );
  AOI22_X1 U918 ( .A1(\REGISTERS[3][8] ), .A2(n139), .B1(\REGISTERS[2][8] ), 
        .B2(n136), .ZN(n987) );
  OAI221_X1 U919 ( .B1(n193), .B2(n2049), .C1(n190), .C2(n2017), .A(n961), 
        .ZN(n960) );
  AOI22_X1 U920 ( .A1(\REGISTERS[19][9] ), .A2(n187), .B1(\REGISTERS[18][9] ), 
        .B2(n184), .ZN(n961) );
  OAI221_X1 U921 ( .B1(n145), .B2(n1793), .C1(n142), .C2(n497), .A(n969), .ZN(
        n968) );
  AOI22_X1 U922 ( .A1(\REGISTERS[3][9] ), .A2(n139), .B1(\REGISTERS[2][9] ), 
        .B2(n136), .ZN(n969) );
  OAI221_X1 U923 ( .B1(n193), .B2(n2048), .C1(n190), .C2(n2016), .A(n943), 
        .ZN(n942) );
  AOI22_X1 U924 ( .A1(\REGISTERS[19][10] ), .A2(n187), .B1(\REGISTERS[18][10] ), .B2(n184), .ZN(n943) );
  OAI221_X1 U925 ( .B1(n145), .B2(n1792), .C1(n142), .C2(n496), .A(n951), .ZN(
        n950) );
  AOI22_X1 U926 ( .A1(\REGISTERS[3][10] ), .A2(n139), .B1(\REGISTERS[2][10] ), 
        .B2(n136), .ZN(n951) );
  OAI221_X1 U927 ( .B1(n193), .B2(n2047), .C1(n191), .C2(n2015), .A(n925), 
        .ZN(n924) );
  AOI22_X1 U928 ( .A1(\REGISTERS[19][11] ), .A2(n187), .B1(\REGISTERS[18][11] ), .B2(n184), .ZN(n925) );
  OAI221_X1 U929 ( .B1(n145), .B2(n1791), .C1(n143), .C2(n495), .A(n933), .ZN(
        n932) );
  AOI22_X1 U930 ( .A1(\REGISTERS[3][11] ), .A2(n139), .B1(\REGISTERS[2][11] ), 
        .B2(n136), .ZN(n933) );
  OAI221_X1 U931 ( .B1(n194), .B2(n2046), .C1(n191), .C2(n2014), .A(n907), 
        .ZN(n906) );
  AOI22_X1 U932 ( .A1(\REGISTERS[19][12] ), .A2(n188), .B1(\REGISTERS[18][12] ), .B2(n185), .ZN(n907) );
  OAI221_X1 U933 ( .B1(n146), .B2(n526), .C1(n143), .C2(n494), .A(n915), .ZN(
        n914) );
  AOI22_X1 U934 ( .A1(\REGISTERS[3][12] ), .A2(n140), .B1(\REGISTERS[2][12] ), 
        .B2(n137), .ZN(n915) );
  OAI221_X1 U935 ( .B1(n194), .B2(n2045), .C1(n191), .C2(n2013), .A(n889), 
        .ZN(n888) );
  AOI22_X1 U936 ( .A1(\REGISTERS[19][13] ), .A2(n188), .B1(\REGISTERS[18][13] ), .B2(n185), .ZN(n889) );
  OAI221_X1 U937 ( .B1(n146), .B2(n525), .C1(n143), .C2(n493), .A(n897), .ZN(
        n896) );
  AOI22_X1 U938 ( .A1(\REGISTERS[3][13] ), .A2(n140), .B1(\REGISTERS[2][13] ), 
        .B2(n137), .ZN(n897) );
  OAI221_X1 U939 ( .B1(n194), .B2(n2044), .C1(n191), .C2(n2012), .A(n871), 
        .ZN(n870) );
  AOI22_X1 U940 ( .A1(\REGISTERS[19][14] ), .A2(n188), .B1(\REGISTERS[18][14] ), .B2(n185), .ZN(n871) );
  OAI221_X1 U941 ( .B1(n146), .B2(n524), .C1(n143), .C2(n492), .A(n879), .ZN(
        n878) );
  AOI22_X1 U942 ( .A1(\REGISTERS[3][14] ), .A2(n140), .B1(\REGISTERS[2][14] ), 
        .B2(n137), .ZN(n879) );
  OAI221_X1 U943 ( .B1(n194), .B2(n2043), .C1(n191), .C2(n2011), .A(n853), 
        .ZN(n852) );
  AOI22_X1 U944 ( .A1(\REGISTERS[19][15] ), .A2(n188), .B1(\REGISTERS[18][15] ), .B2(n185), .ZN(n853) );
  OAI221_X1 U945 ( .B1(n146), .B2(n523), .C1(n143), .C2(n491), .A(n861), .ZN(
        n860) );
  AOI22_X1 U946 ( .A1(\REGISTERS[3][15] ), .A2(n140), .B1(\REGISTERS[2][15] ), 
        .B2(n137), .ZN(n861) );
  OAI221_X1 U947 ( .B1(n194), .B2(n2042), .C1(n191), .C2(n2010), .A(n835), 
        .ZN(n834) );
  AOI22_X1 U948 ( .A1(\REGISTERS[19][16] ), .A2(n188), .B1(\REGISTERS[18][16] ), .B2(n185), .ZN(n835) );
  OAI221_X1 U949 ( .B1(n146), .B2(n522), .C1(n143), .C2(n490), .A(n843), .ZN(
        n842) );
  AOI22_X1 U950 ( .A1(\REGISTERS[3][16] ), .A2(n140), .B1(\REGISTERS[2][16] ), 
        .B2(n137), .ZN(n843) );
  OAI221_X1 U951 ( .B1(n194), .B2(n2041), .C1(n191), .C2(n2009), .A(n817), 
        .ZN(n816) );
  AOI22_X1 U952 ( .A1(\REGISTERS[19][17] ), .A2(n188), .B1(\REGISTERS[18][17] ), .B2(n185), .ZN(n817) );
  OAI221_X1 U953 ( .B1(n146), .B2(n521), .C1(n143), .C2(n489), .A(n825), .ZN(
        n824) );
  AOI22_X1 U954 ( .A1(\REGISTERS[3][17] ), .A2(n140), .B1(\REGISTERS[2][17] ), 
        .B2(n137), .ZN(n825) );
  OAI221_X1 U955 ( .B1(n194), .B2(n2040), .C1(n191), .C2(n2008), .A(n799), 
        .ZN(n798) );
  AOI22_X1 U956 ( .A1(\REGISTERS[19][18] ), .A2(n188), .B1(\REGISTERS[18][18] ), .B2(n185), .ZN(n799) );
  OAI221_X1 U957 ( .B1(n146), .B2(n520), .C1(n143), .C2(n488), .A(n807), .ZN(
        n806) );
  AOI22_X1 U958 ( .A1(\REGISTERS[3][18] ), .A2(n140), .B1(\REGISTERS[2][18] ), 
        .B2(n137), .ZN(n807) );
  OAI221_X1 U959 ( .B1(n194), .B2(n2039), .C1(n191), .C2(n2007), .A(n781), 
        .ZN(n780) );
  AOI22_X1 U960 ( .A1(\REGISTERS[19][19] ), .A2(n188), .B1(\REGISTERS[18][19] ), .B2(n185), .ZN(n781) );
  OAI221_X1 U961 ( .B1(n146), .B2(n519), .C1(n143), .C2(n487), .A(n789), .ZN(
        n788) );
  AOI22_X1 U962 ( .A1(\REGISTERS[3][19] ), .A2(n140), .B1(\REGISTERS[2][19] ), 
        .B2(n137), .ZN(n789) );
  OAI221_X1 U963 ( .B1(n194), .B2(n2038), .C1(n191), .C2(n2006), .A(n763), 
        .ZN(n762) );
  AOI22_X1 U964 ( .A1(\REGISTERS[19][20] ), .A2(n188), .B1(\REGISTERS[18][20] ), .B2(n185), .ZN(n763) );
  OAI221_X1 U965 ( .B1(n146), .B2(n518), .C1(n143), .C2(n486), .A(n771), .ZN(
        n770) );
  AOI22_X1 U966 ( .A1(\REGISTERS[3][20] ), .A2(n140), .B1(\REGISTERS[2][20] ), 
        .B2(n137), .ZN(n771) );
  OAI221_X1 U967 ( .B1(n194), .B2(n2037), .C1(n191), .C2(n2005), .A(n745), 
        .ZN(n744) );
  AOI22_X1 U968 ( .A1(\REGISTERS[19][21] ), .A2(n188), .B1(\REGISTERS[18][21] ), .B2(n185), .ZN(n745) );
  OAI221_X1 U969 ( .B1(n146), .B2(n517), .C1(n143), .C2(n485), .A(n753), .ZN(
        n752) );
  AOI22_X1 U970 ( .A1(\REGISTERS[3][21] ), .A2(n140), .B1(\REGISTERS[2][21] ), 
        .B2(n137), .ZN(n753) );
  OAI221_X1 U971 ( .B1(n194), .B2(n2036), .C1(n192), .C2(n2004), .A(n727), 
        .ZN(n726) );
  AOI22_X1 U972 ( .A1(\REGISTERS[19][22] ), .A2(n188), .B1(\REGISTERS[18][22] ), .B2(n185), .ZN(n727) );
  OAI221_X1 U973 ( .B1(n146), .B2(n516), .C1(n144), .C2(n484), .A(n735), .ZN(
        n734) );
  AOI22_X1 U974 ( .A1(\REGISTERS[3][22] ), .A2(n140), .B1(\REGISTERS[2][22] ), 
        .B2(n137), .ZN(n735) );
  OAI221_X1 U975 ( .B1(n194), .B2(n2035), .C1(n192), .C2(n2003), .A(n709), 
        .ZN(n708) );
  AOI22_X1 U976 ( .A1(\REGISTERS[19][23] ), .A2(n188), .B1(\REGISTERS[18][23] ), .B2(n185), .ZN(n709) );
  OAI221_X1 U977 ( .B1(n146), .B2(n515), .C1(n144), .C2(n483), .A(n717), .ZN(
        n716) );
  AOI22_X1 U978 ( .A1(\REGISTERS[3][23] ), .A2(n140), .B1(\REGISTERS[2][23] ), 
        .B2(n137), .ZN(n717) );
  OAI221_X1 U979 ( .B1(n2047), .B2(n98), .C1(n2015), .C2(n95), .A(n1550), .ZN(
        n1549) );
  AOI22_X1 U980 ( .A1(n92), .A2(\REGISTERS[19][11] ), .B1(n89), .B2(
        \REGISTERS[18][11] ), .ZN(n1550) );
  OAI221_X1 U981 ( .B1(n1791), .B2(n50), .C1(n495), .C2(n47), .A(n1558), .ZN(
        n1557) );
  AOI22_X1 U982 ( .A1(n44), .A2(\REGISTERS[3][11] ), .B1(n41), .B2(
        \REGISTERS[2][11] ), .ZN(n1558) );
  OAI221_X1 U983 ( .B1(n2046), .B2(n98), .C1(n2014), .C2(n95), .A(n1532), .ZN(
        n1531) );
  AOI22_X1 U984 ( .A1(n92), .A2(\REGISTERS[19][12] ), .B1(n89), .B2(
        \REGISTERS[18][12] ), .ZN(n1532) );
  OAI221_X1 U985 ( .B1(n526), .B2(n50), .C1(n494), .C2(n47), .A(n1540), .ZN(
        n1539) );
  AOI22_X1 U986 ( .A1(n44), .A2(\REGISTERS[3][12] ), .B1(n41), .B2(
        \REGISTERS[2][12] ), .ZN(n1540) );
  OAI221_X1 U987 ( .B1(n2045), .B2(n98), .C1(n2013), .C2(n95), .A(n1514), .ZN(
        n1513) );
  AOI22_X1 U988 ( .A1(n92), .A2(\REGISTERS[19][13] ), .B1(n89), .B2(
        \REGISTERS[18][13] ), .ZN(n1514) );
  OAI221_X1 U989 ( .B1(n525), .B2(n50), .C1(n493), .C2(n47), .A(n1522), .ZN(
        n1521) );
  AOI22_X1 U990 ( .A1(n44), .A2(\REGISTERS[3][13] ), .B1(n41), .B2(
        \REGISTERS[2][13] ), .ZN(n1522) );
  OAI221_X1 U991 ( .B1(n2044), .B2(n98), .C1(n2012), .C2(n95), .A(n1496), .ZN(
        n1495) );
  AOI22_X1 U992 ( .A1(n92), .A2(\REGISTERS[19][14] ), .B1(n89), .B2(
        \REGISTERS[18][14] ), .ZN(n1496) );
  OAI221_X1 U993 ( .B1(n524), .B2(n50), .C1(n492), .C2(n47), .A(n1504), .ZN(
        n1503) );
  AOI22_X1 U994 ( .A1(n44), .A2(\REGISTERS[3][14] ), .B1(n41), .B2(
        \REGISTERS[2][14] ), .ZN(n1504) );
  OAI221_X1 U995 ( .B1(n2043), .B2(n98), .C1(n2011), .C2(n95), .A(n1478), .ZN(
        n1477) );
  AOI22_X1 U996 ( .A1(n92), .A2(\REGISTERS[19][15] ), .B1(n89), .B2(
        \REGISTERS[18][15] ), .ZN(n1478) );
  OAI221_X1 U997 ( .B1(n523), .B2(n50), .C1(n491), .C2(n47), .A(n1486), .ZN(
        n1485) );
  AOI22_X1 U998 ( .A1(n44), .A2(\REGISTERS[3][15] ), .B1(n41), .B2(
        \REGISTERS[2][15] ), .ZN(n1486) );
  OAI221_X1 U999 ( .B1(n2042), .B2(n98), .C1(n2010), .C2(n95), .A(n1460), .ZN(
        n1459) );
  AOI22_X1 U1000 ( .A1(n92), .A2(\REGISTERS[19][16] ), .B1(n89), .B2(
        \REGISTERS[18][16] ), .ZN(n1460) );
  OAI221_X1 U1001 ( .B1(n522), .B2(n50), .C1(n490), .C2(n47), .A(n1468), .ZN(
        n1467) );
  AOI22_X1 U1002 ( .A1(n44), .A2(\REGISTERS[3][16] ), .B1(n41), .B2(
        \REGISTERS[2][16] ), .ZN(n1468) );
  OAI221_X1 U1003 ( .B1(n2041), .B2(n98), .C1(n2009), .C2(n95), .A(n1442), 
        .ZN(n1441) );
  AOI22_X1 U1004 ( .A1(n92), .A2(\REGISTERS[19][17] ), .B1(n89), .B2(
        \REGISTERS[18][17] ), .ZN(n1442) );
  OAI221_X1 U1005 ( .B1(n521), .B2(n50), .C1(n489), .C2(n47), .A(n1450), .ZN(
        n1449) );
  AOI22_X1 U1006 ( .A1(n44), .A2(\REGISTERS[3][17] ), .B1(n41), .B2(
        \REGISTERS[2][17] ), .ZN(n1450) );
  OAI221_X1 U1007 ( .B1(n2040), .B2(n98), .C1(n2008), .C2(n95), .A(n1424), 
        .ZN(n1423) );
  AOI22_X1 U1008 ( .A1(n92), .A2(\REGISTERS[19][18] ), .B1(n89), .B2(
        \REGISTERS[18][18] ), .ZN(n1424) );
  OAI221_X1 U1009 ( .B1(n520), .B2(n50), .C1(n488), .C2(n47), .A(n1432), .ZN(
        n1431) );
  AOI22_X1 U1010 ( .A1(n44), .A2(\REGISTERS[3][18] ), .B1(n41), .B2(
        \REGISTERS[2][18] ), .ZN(n1432) );
  OAI221_X1 U1011 ( .B1(n2039), .B2(n98), .C1(n2007), .C2(n95), .A(n1406), 
        .ZN(n1405) );
  AOI22_X1 U1012 ( .A1(n92), .A2(\REGISTERS[19][19] ), .B1(n89), .B2(
        \REGISTERS[18][19] ), .ZN(n1406) );
  OAI221_X1 U1013 ( .B1(n519), .B2(n50), .C1(n487), .C2(n47), .A(n1414), .ZN(
        n1413) );
  AOI22_X1 U1014 ( .A1(n44), .A2(\REGISTERS[3][19] ), .B1(n41), .B2(
        \REGISTERS[2][19] ), .ZN(n1414) );
  OAI221_X1 U1015 ( .B1(n2038), .B2(n98), .C1(n2006), .C2(n95), .A(n1388), 
        .ZN(n1387) );
  AOI22_X1 U1016 ( .A1(n92), .A2(\REGISTERS[19][20] ), .B1(n89), .B2(
        \REGISTERS[18][20] ), .ZN(n1388) );
  OAI221_X1 U1017 ( .B1(n518), .B2(n50), .C1(n486), .C2(n47), .A(n1396), .ZN(
        n1395) );
  AOI22_X1 U1018 ( .A1(n44), .A2(\REGISTERS[3][20] ), .B1(n41), .B2(
        \REGISTERS[2][20] ), .ZN(n1396) );
  OAI221_X1 U1019 ( .B1(n2037), .B2(n98), .C1(n2005), .C2(n95), .A(n1370), 
        .ZN(n1369) );
  AOI22_X1 U1020 ( .A1(n92), .A2(\REGISTERS[19][21] ), .B1(n89), .B2(
        \REGISTERS[18][21] ), .ZN(n1370) );
  OAI221_X1 U1021 ( .B1(n517), .B2(n50), .C1(n485), .C2(n47), .A(n1378), .ZN(
        n1377) );
  AOI22_X1 U1022 ( .A1(n44), .A2(\REGISTERS[3][21] ), .B1(n41), .B2(
        \REGISTERS[2][21] ), .ZN(n1378) );
  OAI221_X1 U1023 ( .B1(n2122), .B2(n85), .C1(n2090), .C2(n82), .A(n1753), 
        .ZN(n1746) );
  AOI22_X1 U1024 ( .A1(n79), .A2(\REGISTERS[23][0] ), .B1(n76), .B2(
        \REGISTERS[22][0] ), .ZN(n1753) );
  OAI221_X1 U1025 ( .B1(n1866), .B2(n37), .C1(n1834), .C2(n34), .A(n1769), 
        .ZN(n1764) );
  AOI22_X1 U1026 ( .A1(n31), .A2(\REGISTERS[7][0] ), .B1(n28), .B2(
        \REGISTERS[6][0] ), .ZN(n1769) );
  OAI221_X1 U1027 ( .B1(n2121), .B2(n85), .C1(n2089), .C2(n82), .A(n1731), 
        .ZN(n1728) );
  AOI22_X1 U1028 ( .A1(n79), .A2(\REGISTERS[23][1] ), .B1(n76), .B2(
        \REGISTERS[22][1] ), .ZN(n1731) );
  OAI221_X1 U1029 ( .B1(n1865), .B2(n37), .C1(n1833), .C2(n34), .A(n1739), 
        .ZN(n1736) );
  AOI22_X1 U1030 ( .A1(n31), .A2(\REGISTERS[7][1] ), .B1(n28), .B2(
        \REGISTERS[6][1] ), .ZN(n1739) );
  OAI221_X1 U1031 ( .B1(n2120), .B2(n85), .C1(n2088), .C2(n82), .A(n1713), 
        .ZN(n1710) );
  AOI22_X1 U1032 ( .A1(n79), .A2(\REGISTERS[23][2] ), .B1(n76), .B2(
        \REGISTERS[22][2] ), .ZN(n1713) );
  OAI221_X1 U1033 ( .B1(n1864), .B2(n37), .C1(n1832), .C2(n34), .A(n1721), 
        .ZN(n1718) );
  AOI22_X1 U1034 ( .A1(n31), .A2(\REGISTERS[7][2] ), .B1(n28), .B2(
        \REGISTERS[6][2] ), .ZN(n1721) );
  OAI221_X1 U1035 ( .B1(n2119), .B2(n85), .C1(n2087), .C2(n82), .A(n1695), 
        .ZN(n1692) );
  AOI22_X1 U1036 ( .A1(n79), .A2(\REGISTERS[23][3] ), .B1(n76), .B2(
        \REGISTERS[22][3] ), .ZN(n1695) );
  OAI221_X1 U1037 ( .B1(n1863), .B2(n37), .C1(n1831), .C2(n34), .A(n1703), 
        .ZN(n1700) );
  AOI22_X1 U1038 ( .A1(n31), .A2(\REGISTERS[7][3] ), .B1(n28), .B2(
        \REGISTERS[6][3] ), .ZN(n1703) );
  OAI221_X1 U1039 ( .B1(n2118), .B2(n85), .C1(n2086), .C2(n82), .A(n1677), 
        .ZN(n1674) );
  AOI22_X1 U1040 ( .A1(n79), .A2(\REGISTERS[23][4] ), .B1(n76), .B2(
        \REGISTERS[22][4] ), .ZN(n1677) );
  OAI221_X1 U1041 ( .B1(n1862), .B2(n37), .C1(n1830), .C2(n34), .A(n1685), 
        .ZN(n1682) );
  AOI22_X1 U1042 ( .A1(n31), .A2(\REGISTERS[7][4] ), .B1(n28), .B2(
        \REGISTERS[6][4] ), .ZN(n1685) );
  OAI221_X1 U1043 ( .B1(n2117), .B2(n85), .C1(n2085), .C2(n82), .A(n1659), 
        .ZN(n1656) );
  AOI22_X1 U1044 ( .A1(n79), .A2(\REGISTERS[23][5] ), .B1(n76), .B2(
        \REGISTERS[22][5] ), .ZN(n1659) );
  OAI221_X1 U1045 ( .B1(n1861), .B2(n37), .C1(n1829), .C2(n34), .A(n1667), 
        .ZN(n1664) );
  AOI22_X1 U1046 ( .A1(n31), .A2(\REGISTERS[7][5] ), .B1(n28), .B2(
        \REGISTERS[6][5] ), .ZN(n1667) );
  OAI221_X1 U1047 ( .B1(n2116), .B2(n85), .C1(n2084), .C2(n82), .A(n1641), 
        .ZN(n1638) );
  AOI22_X1 U1048 ( .A1(n79), .A2(\REGISTERS[23][6] ), .B1(n76), .B2(
        \REGISTERS[22][6] ), .ZN(n1641) );
  OAI221_X1 U1049 ( .B1(n1860), .B2(n37), .C1(n1828), .C2(n34), .A(n1649), 
        .ZN(n1646) );
  AOI22_X1 U1050 ( .A1(n31), .A2(\REGISTERS[7][6] ), .B1(n28), .B2(
        \REGISTERS[6][6] ), .ZN(n1649) );
  OAI221_X1 U1051 ( .B1(n2115), .B2(n85), .C1(n2083), .C2(n82), .A(n1623), 
        .ZN(n1620) );
  AOI22_X1 U1052 ( .A1(n79), .A2(\REGISTERS[23][7] ), .B1(n76), .B2(
        \REGISTERS[22][7] ), .ZN(n1623) );
  OAI221_X1 U1053 ( .B1(n1859), .B2(n37), .C1(n1827), .C2(n34), .A(n1631), 
        .ZN(n1628) );
  AOI22_X1 U1054 ( .A1(n31), .A2(\REGISTERS[7][7] ), .B1(n28), .B2(
        \REGISTERS[6][7] ), .ZN(n1631) );
  OAI221_X1 U1055 ( .B1(n2114), .B2(n85), .C1(n2082), .C2(n82), .A(n1605), 
        .ZN(n1602) );
  AOI22_X1 U1056 ( .A1(n79), .A2(\REGISTERS[23][8] ), .B1(n76), .B2(
        \REGISTERS[22][8] ), .ZN(n1605) );
  OAI221_X1 U1057 ( .B1(n1858), .B2(n37), .C1(n1826), .C2(n34), .A(n1613), 
        .ZN(n1610) );
  AOI22_X1 U1058 ( .A1(n31), .A2(\REGISTERS[7][8] ), .B1(n28), .B2(
        \REGISTERS[6][8] ), .ZN(n1613) );
  OAI221_X1 U1059 ( .B1(n2113), .B2(n85), .C1(n2081), .C2(n82), .A(n1587), 
        .ZN(n1584) );
  AOI22_X1 U1060 ( .A1(n79), .A2(\REGISTERS[23][9] ), .B1(n76), .B2(
        \REGISTERS[22][9] ), .ZN(n1587) );
  OAI221_X1 U1061 ( .B1(n1857), .B2(n37), .C1(n1825), .C2(n34), .A(n1595), 
        .ZN(n1592) );
  AOI22_X1 U1062 ( .A1(n31), .A2(\REGISTERS[7][9] ), .B1(n28), .B2(
        \REGISTERS[6][9] ), .ZN(n1595) );
  OAI221_X1 U1063 ( .B1(n2112), .B2(n85), .C1(n2080), .C2(n82), .A(n1569), 
        .ZN(n1566) );
  AOI22_X1 U1064 ( .A1(n79), .A2(\REGISTERS[23][10] ), .B1(n76), .B2(
        \REGISTERS[22][10] ), .ZN(n1569) );
  OAI221_X1 U1065 ( .B1(n1856), .B2(n37), .C1(n1824), .C2(n34), .A(n1577), 
        .ZN(n1574) );
  AOI22_X1 U1066 ( .A1(n31), .A2(\REGISTERS[7][10] ), .B1(n28), .B2(
        \REGISTERS[6][10] ), .ZN(n1577) );
  OAI221_X1 U1067 ( .B1(n2100), .B2(n87), .C1(n2068), .C2(n84), .A(n1353), 
        .ZN(n1350) );
  AOI22_X1 U1068 ( .A1(n81), .A2(\REGISTERS[23][22] ), .B1(n78), .B2(
        \REGISTERS[22][22] ), .ZN(n1353) );
  OAI221_X1 U1069 ( .B1(n1844), .B2(n39), .C1(n1812), .C2(n36), .A(n1361), 
        .ZN(n1358) );
  AOI22_X1 U1070 ( .A1(n33), .A2(\REGISTERS[7][22] ), .B1(n30), .B2(
        \REGISTERS[6][22] ), .ZN(n1361) );
  OAI221_X1 U1071 ( .B1(n2099), .B2(n87), .C1(n2067), .C2(n84), .A(n1335), 
        .ZN(n1332) );
  AOI22_X1 U1072 ( .A1(n81), .A2(\REGISTERS[23][23] ), .B1(n78), .B2(
        \REGISTERS[22][23] ), .ZN(n1335) );
  OAI221_X1 U1073 ( .B1(n1843), .B2(n39), .C1(n1811), .C2(n36), .A(n1343), 
        .ZN(n1340) );
  AOI22_X1 U1074 ( .A1(n33), .A2(\REGISTERS[7][23] ), .B1(n30), .B2(
        \REGISTERS[6][23] ), .ZN(n1343) );
  OAI221_X1 U1075 ( .B1(n2098), .B2(n87), .C1(n2066), .C2(n84), .A(n1317), 
        .ZN(n1314) );
  AOI22_X1 U1076 ( .A1(n81), .A2(\REGISTERS[23][24] ), .B1(n78), .B2(
        \REGISTERS[22][24] ), .ZN(n1317) );
  OAI221_X1 U1077 ( .B1(n1842), .B2(n39), .C1(n1810), .C2(n36), .A(n1325), 
        .ZN(n1322) );
  AOI22_X1 U1078 ( .A1(n33), .A2(\REGISTERS[7][24] ), .B1(n30), .B2(
        \REGISTERS[6][24] ), .ZN(n1325) );
  OAI221_X1 U1079 ( .B1(n2097), .B2(n87), .C1(n2065), .C2(n84), .A(n1299), 
        .ZN(n1296) );
  AOI22_X1 U1080 ( .A1(n81), .A2(\REGISTERS[23][25] ), .B1(n78), .B2(
        \REGISTERS[22][25] ), .ZN(n1299) );
  OAI221_X1 U1081 ( .B1(n1841), .B2(n39), .C1(n1809), .C2(n36), .A(n1307), 
        .ZN(n1304) );
  AOI22_X1 U1082 ( .A1(n33), .A2(\REGISTERS[7][25] ), .B1(n30), .B2(
        \REGISTERS[6][25] ), .ZN(n1307) );
  OAI221_X1 U1083 ( .B1(n2096), .B2(n87), .C1(n2064), .C2(n84), .A(n1281), 
        .ZN(n1278) );
  AOI22_X1 U1084 ( .A1(n81), .A2(\REGISTERS[23][26] ), .B1(n78), .B2(
        \REGISTERS[22][26] ), .ZN(n1281) );
  OAI221_X1 U1085 ( .B1(n1840), .B2(n39), .C1(n1808), .C2(n36), .A(n1289), 
        .ZN(n1286) );
  AOI22_X1 U1086 ( .A1(n33), .A2(\REGISTERS[7][26] ), .B1(n30), .B2(
        \REGISTERS[6][26] ), .ZN(n1289) );
  OAI221_X1 U1087 ( .B1(n2095), .B2(n87), .C1(n2063), .C2(n84), .A(n1263), 
        .ZN(n1260) );
  AOI22_X1 U1088 ( .A1(n81), .A2(\REGISTERS[23][27] ), .B1(n78), .B2(
        \REGISTERS[22][27] ), .ZN(n1263) );
  OAI221_X1 U1089 ( .B1(n1839), .B2(n39), .C1(n1807), .C2(n36), .A(n1271), 
        .ZN(n1268) );
  AOI22_X1 U1090 ( .A1(n33), .A2(\REGISTERS[7][27] ), .B1(n30), .B2(
        \REGISTERS[6][27] ), .ZN(n1271) );
  OAI221_X1 U1091 ( .B1(n2094), .B2(n87), .C1(n2062), .C2(n84), .A(n1245), 
        .ZN(n1242) );
  AOI22_X1 U1092 ( .A1(n81), .A2(\REGISTERS[23][28] ), .B1(n78), .B2(
        \REGISTERS[22][28] ), .ZN(n1245) );
  OAI221_X1 U1093 ( .B1(n1838), .B2(n39), .C1(n1806), .C2(n36), .A(n1253), 
        .ZN(n1250) );
  AOI22_X1 U1094 ( .A1(n33), .A2(\REGISTERS[7][28] ), .B1(n30), .B2(
        \REGISTERS[6][28] ), .ZN(n1253) );
  OAI221_X1 U1095 ( .B1(n2093), .B2(n87), .C1(n2061), .C2(n84), .A(n1227), 
        .ZN(n1224) );
  AOI22_X1 U1096 ( .A1(n81), .A2(\REGISTERS[23][29] ), .B1(n78), .B2(
        \REGISTERS[22][29] ), .ZN(n1227) );
  OAI221_X1 U1097 ( .B1(n1837), .B2(n39), .C1(n1805), .C2(n36), .A(n1235), 
        .ZN(n1232) );
  AOI22_X1 U1098 ( .A1(n33), .A2(\REGISTERS[7][29] ), .B1(n30), .B2(
        \REGISTERS[6][29] ), .ZN(n1235) );
  OAI221_X1 U1099 ( .B1(n2092), .B2(n87), .C1(n2060), .C2(n84), .A(n1209), 
        .ZN(n1206) );
  AOI22_X1 U1100 ( .A1(n81), .A2(\REGISTERS[23][30] ), .B1(n78), .B2(
        \REGISTERS[22][30] ), .ZN(n1209) );
  OAI221_X1 U1101 ( .B1(n1836), .B2(n39), .C1(n1804), .C2(n36), .A(n1217), 
        .ZN(n1214) );
  AOI22_X1 U1102 ( .A1(n33), .A2(\REGISTERS[7][30] ), .B1(n30), .B2(
        \REGISTERS[6][30] ), .ZN(n1217) );
  OAI221_X1 U1103 ( .B1(n2091), .B2(n87), .C1(n2059), .C2(n84), .A(n1165), 
        .ZN(n1156) );
  AOI22_X1 U1104 ( .A1(n81), .A2(\REGISTERS[23][31] ), .B1(n78), .B2(
        \REGISTERS[22][31] ), .ZN(n1165) );
  OAI221_X1 U1105 ( .B1(n1835), .B2(n39), .C1(n1803), .C2(n36), .A(n1189), 
        .ZN(n1180) );
  AOI22_X1 U1106 ( .A1(n33), .A2(\REGISTERS[7][31] ), .B1(n30), .B2(
        \REGISTERS[6][31] ), .ZN(n1189) );
  OAI221_X1 U1107 ( .B1(n181), .B2(n2122), .C1(n178), .C2(n2090), .A(n1128), 
        .ZN(n1121) );
  AOI22_X1 U1108 ( .A1(\REGISTERS[23][0] ), .A2(n175), .B1(\REGISTERS[22][0] ), 
        .B2(n172), .ZN(n1128) );
  OAI221_X1 U1109 ( .B1(n133), .B2(n1866), .C1(n130), .C2(n1834), .A(n1144), 
        .ZN(n1139) );
  AOI22_X1 U1110 ( .A1(\REGISTERS[7][0] ), .A2(n127), .B1(\REGISTERS[6][0] ), 
        .B2(n124), .ZN(n1144) );
  OAI221_X1 U1111 ( .B1(n181), .B2(n2121), .C1(n178), .C2(n2089), .A(n1106), 
        .ZN(n1103) );
  AOI22_X1 U1112 ( .A1(\REGISTERS[23][1] ), .A2(n175), .B1(\REGISTERS[22][1] ), 
        .B2(n172), .ZN(n1106) );
  OAI221_X1 U1113 ( .B1(n133), .B2(n1865), .C1(n130), .C2(n1833), .A(n1114), 
        .ZN(n1111) );
  AOI22_X1 U1114 ( .A1(\REGISTERS[7][1] ), .A2(n127), .B1(\REGISTERS[6][1] ), 
        .B2(n124), .ZN(n1114) );
  OAI221_X1 U1115 ( .B1(n181), .B2(n2120), .C1(n178), .C2(n2088), .A(n1088), 
        .ZN(n1085) );
  AOI22_X1 U1116 ( .A1(\REGISTERS[23][2] ), .A2(n175), .B1(\REGISTERS[22][2] ), 
        .B2(n172), .ZN(n1088) );
  OAI221_X1 U1117 ( .B1(n133), .B2(n1864), .C1(n130), .C2(n1832), .A(n1096), 
        .ZN(n1093) );
  AOI22_X1 U1118 ( .A1(\REGISTERS[7][2] ), .A2(n127), .B1(\REGISTERS[6][2] ), 
        .B2(n124), .ZN(n1096) );
  OAI221_X1 U1119 ( .B1(n181), .B2(n2119), .C1(n178), .C2(n2087), .A(n1070), 
        .ZN(n1067) );
  AOI22_X1 U1120 ( .A1(\REGISTERS[23][3] ), .A2(n175), .B1(\REGISTERS[22][3] ), 
        .B2(n172), .ZN(n1070) );
  OAI221_X1 U1121 ( .B1(n133), .B2(n1863), .C1(n130), .C2(n1831), .A(n1078), 
        .ZN(n1075) );
  AOI22_X1 U1122 ( .A1(\REGISTERS[7][3] ), .A2(n127), .B1(\REGISTERS[6][3] ), 
        .B2(n124), .ZN(n1078) );
  OAI221_X1 U1123 ( .B1(n181), .B2(n2118), .C1(n178), .C2(n2086), .A(n1052), 
        .ZN(n1049) );
  AOI22_X1 U1124 ( .A1(\REGISTERS[23][4] ), .A2(n175), .B1(\REGISTERS[22][4] ), 
        .B2(n172), .ZN(n1052) );
  OAI221_X1 U1125 ( .B1(n133), .B2(n1862), .C1(n130), .C2(n1830), .A(n1060), 
        .ZN(n1057) );
  AOI22_X1 U1126 ( .A1(\REGISTERS[7][4] ), .A2(n127), .B1(\REGISTERS[6][4] ), 
        .B2(n124), .ZN(n1060) );
  OAI221_X1 U1127 ( .B1(n181), .B2(n2117), .C1(n178), .C2(n2085), .A(n1034), 
        .ZN(n1031) );
  AOI22_X1 U1128 ( .A1(\REGISTERS[23][5] ), .A2(n175), .B1(\REGISTERS[22][5] ), 
        .B2(n172), .ZN(n1034) );
  OAI221_X1 U1129 ( .B1(n133), .B2(n1861), .C1(n130), .C2(n1829), .A(n1042), 
        .ZN(n1039) );
  AOI22_X1 U1130 ( .A1(\REGISTERS[7][5] ), .A2(n127), .B1(\REGISTERS[6][5] ), 
        .B2(n124), .ZN(n1042) );
  OAI221_X1 U1131 ( .B1(n181), .B2(n2116), .C1(n178), .C2(n2084), .A(n1016), 
        .ZN(n1013) );
  AOI22_X1 U1132 ( .A1(\REGISTERS[23][6] ), .A2(n175), .B1(\REGISTERS[22][6] ), 
        .B2(n172), .ZN(n1016) );
  OAI221_X1 U1133 ( .B1(n133), .B2(n1860), .C1(n130), .C2(n1828), .A(n1024), 
        .ZN(n1021) );
  AOI22_X1 U1134 ( .A1(\REGISTERS[7][6] ), .A2(n127), .B1(\REGISTERS[6][6] ), 
        .B2(n124), .ZN(n1024) );
  OAI221_X1 U1135 ( .B1(n181), .B2(n2115), .C1(n178), .C2(n2083), .A(n998), 
        .ZN(n995) );
  AOI22_X1 U1136 ( .A1(\REGISTERS[23][7] ), .A2(n175), .B1(\REGISTERS[22][7] ), 
        .B2(n172), .ZN(n998) );
  OAI221_X1 U1137 ( .B1(n133), .B2(n1859), .C1(n130), .C2(n1827), .A(n1006), 
        .ZN(n1003) );
  AOI22_X1 U1138 ( .A1(\REGISTERS[7][7] ), .A2(n127), .B1(\REGISTERS[6][7] ), 
        .B2(n124), .ZN(n1006) );
  OAI221_X1 U1139 ( .B1(n181), .B2(n2114), .C1(n178), .C2(n2082), .A(n980), 
        .ZN(n977) );
  AOI22_X1 U1140 ( .A1(\REGISTERS[23][8] ), .A2(n175), .B1(\REGISTERS[22][8] ), 
        .B2(n172), .ZN(n980) );
  OAI221_X1 U1141 ( .B1(n133), .B2(n1858), .C1(n130), .C2(n1826), .A(n988), 
        .ZN(n985) );
  AOI22_X1 U1142 ( .A1(\REGISTERS[7][8] ), .A2(n127), .B1(\REGISTERS[6][8] ), 
        .B2(n124), .ZN(n988) );
  OAI221_X1 U1143 ( .B1(n181), .B2(n2113), .C1(n178), .C2(n2081), .A(n962), 
        .ZN(n959) );
  AOI22_X1 U1144 ( .A1(\REGISTERS[23][9] ), .A2(n175), .B1(\REGISTERS[22][9] ), 
        .B2(n172), .ZN(n962) );
  OAI221_X1 U1145 ( .B1(n133), .B2(n1857), .C1(n130), .C2(n1825), .A(n970), 
        .ZN(n967) );
  AOI22_X1 U1146 ( .A1(\REGISTERS[7][9] ), .A2(n127), .B1(\REGISTERS[6][9] ), 
        .B2(n124), .ZN(n970) );
  OAI221_X1 U1147 ( .B1(n181), .B2(n2112), .C1(n178), .C2(n2080), .A(n944), 
        .ZN(n941) );
  AOI22_X1 U1148 ( .A1(\REGISTERS[23][10] ), .A2(n175), .B1(
        \REGISTERS[22][10] ), .B2(n172), .ZN(n944) );
  OAI221_X1 U1149 ( .B1(n133), .B2(n1856), .C1(n130), .C2(n1824), .A(n952), 
        .ZN(n949) );
  AOI22_X1 U1150 ( .A1(\REGISTERS[7][10] ), .A2(n127), .B1(\REGISTERS[6][10] ), 
        .B2(n124), .ZN(n952) );
  OAI221_X1 U1151 ( .B1(n181), .B2(n2111), .C1(n179), .C2(n2079), .A(n926), 
        .ZN(n923) );
  AOI22_X1 U1152 ( .A1(\REGISTERS[23][11] ), .A2(n175), .B1(
        \REGISTERS[22][11] ), .B2(n172), .ZN(n926) );
  OAI221_X1 U1153 ( .B1(n133), .B2(n1855), .C1(n131), .C2(n1823), .A(n934), 
        .ZN(n931) );
  AOI22_X1 U1154 ( .A1(\REGISTERS[7][11] ), .A2(n127), .B1(\REGISTERS[6][11] ), 
        .B2(n124), .ZN(n934) );
  OAI221_X1 U1155 ( .B1(n182), .B2(n2110), .C1(n179), .C2(n2078), .A(n908), 
        .ZN(n905) );
  AOI22_X1 U1156 ( .A1(\REGISTERS[23][12] ), .A2(n176), .B1(
        \REGISTERS[22][12] ), .B2(n173), .ZN(n908) );
  OAI221_X1 U1157 ( .B1(n134), .B2(n1854), .C1(n131), .C2(n1822), .A(n916), 
        .ZN(n913) );
  AOI22_X1 U1158 ( .A1(\REGISTERS[7][12] ), .A2(n128), .B1(\REGISTERS[6][12] ), 
        .B2(n125), .ZN(n916) );
  OAI221_X1 U1159 ( .B1(n182), .B2(n2109), .C1(n179), .C2(n2077), .A(n890), 
        .ZN(n887) );
  AOI22_X1 U1160 ( .A1(\REGISTERS[23][13] ), .A2(n176), .B1(
        \REGISTERS[22][13] ), .B2(n173), .ZN(n890) );
  OAI221_X1 U1161 ( .B1(n134), .B2(n1853), .C1(n131), .C2(n1821), .A(n898), 
        .ZN(n895) );
  AOI22_X1 U1162 ( .A1(\REGISTERS[7][13] ), .A2(n128), .B1(\REGISTERS[6][13] ), 
        .B2(n125), .ZN(n898) );
  OAI221_X1 U1163 ( .B1(n182), .B2(n2108), .C1(n179), .C2(n2076), .A(n872), 
        .ZN(n869) );
  AOI22_X1 U1164 ( .A1(\REGISTERS[23][14] ), .A2(n176), .B1(
        \REGISTERS[22][14] ), .B2(n173), .ZN(n872) );
  OAI221_X1 U1165 ( .B1(n134), .B2(n1852), .C1(n131), .C2(n1820), .A(n880), 
        .ZN(n877) );
  AOI22_X1 U1166 ( .A1(\REGISTERS[7][14] ), .A2(n128), .B1(\REGISTERS[6][14] ), 
        .B2(n125), .ZN(n880) );
  OAI221_X1 U1167 ( .B1(n182), .B2(n2107), .C1(n179), .C2(n2075), .A(n854), 
        .ZN(n851) );
  AOI22_X1 U1168 ( .A1(\REGISTERS[23][15] ), .A2(n176), .B1(
        \REGISTERS[22][15] ), .B2(n173), .ZN(n854) );
  OAI221_X1 U1169 ( .B1(n134), .B2(n1851), .C1(n131), .C2(n1819), .A(n862), 
        .ZN(n859) );
  AOI22_X1 U1170 ( .A1(\REGISTERS[7][15] ), .A2(n128), .B1(\REGISTERS[6][15] ), 
        .B2(n125), .ZN(n862) );
  OAI221_X1 U1171 ( .B1(n182), .B2(n2106), .C1(n179), .C2(n2074), .A(n836), 
        .ZN(n833) );
  AOI22_X1 U1172 ( .A1(\REGISTERS[23][16] ), .A2(n176), .B1(
        \REGISTERS[22][16] ), .B2(n173), .ZN(n836) );
  OAI221_X1 U1173 ( .B1(n134), .B2(n1850), .C1(n131), .C2(n1818), .A(n844), 
        .ZN(n841) );
  AOI22_X1 U1174 ( .A1(\REGISTERS[7][16] ), .A2(n128), .B1(\REGISTERS[6][16] ), 
        .B2(n125), .ZN(n844) );
  OAI221_X1 U1175 ( .B1(n182), .B2(n2105), .C1(n179), .C2(n2073), .A(n818), 
        .ZN(n815) );
  AOI22_X1 U1176 ( .A1(\REGISTERS[23][17] ), .A2(n176), .B1(
        \REGISTERS[22][17] ), .B2(n173), .ZN(n818) );
  OAI221_X1 U1177 ( .B1(n134), .B2(n1849), .C1(n131), .C2(n1817), .A(n826), 
        .ZN(n823) );
  AOI22_X1 U1178 ( .A1(\REGISTERS[7][17] ), .A2(n128), .B1(\REGISTERS[6][17] ), 
        .B2(n125), .ZN(n826) );
  OAI221_X1 U1179 ( .B1(n182), .B2(n2104), .C1(n179), .C2(n2072), .A(n800), 
        .ZN(n797) );
  AOI22_X1 U1180 ( .A1(\REGISTERS[23][18] ), .A2(n176), .B1(
        \REGISTERS[22][18] ), .B2(n173), .ZN(n800) );
  OAI221_X1 U1181 ( .B1(n134), .B2(n1848), .C1(n131), .C2(n1816), .A(n808), 
        .ZN(n805) );
  AOI22_X1 U1182 ( .A1(\REGISTERS[7][18] ), .A2(n128), .B1(\REGISTERS[6][18] ), 
        .B2(n125), .ZN(n808) );
  OAI221_X1 U1183 ( .B1(n182), .B2(n2103), .C1(n179), .C2(n2071), .A(n782), 
        .ZN(n779) );
  AOI22_X1 U1184 ( .A1(\REGISTERS[23][19] ), .A2(n176), .B1(
        \REGISTERS[22][19] ), .B2(n173), .ZN(n782) );
  OAI221_X1 U1185 ( .B1(n134), .B2(n1847), .C1(n131), .C2(n1815), .A(n790), 
        .ZN(n787) );
  AOI22_X1 U1186 ( .A1(\REGISTERS[7][19] ), .A2(n128), .B1(\REGISTERS[6][19] ), 
        .B2(n125), .ZN(n790) );
  OAI221_X1 U1187 ( .B1(n182), .B2(n2102), .C1(n179), .C2(n2070), .A(n764), 
        .ZN(n761) );
  AOI22_X1 U1188 ( .A1(\REGISTERS[23][20] ), .A2(n176), .B1(
        \REGISTERS[22][20] ), .B2(n173), .ZN(n764) );
  OAI221_X1 U1189 ( .B1(n134), .B2(n1846), .C1(n131), .C2(n1814), .A(n772), 
        .ZN(n769) );
  AOI22_X1 U1190 ( .A1(\REGISTERS[7][20] ), .A2(n128), .B1(\REGISTERS[6][20] ), 
        .B2(n125), .ZN(n772) );
  OAI221_X1 U1191 ( .B1(n182), .B2(n2101), .C1(n179), .C2(n2069), .A(n746), 
        .ZN(n743) );
  AOI22_X1 U1192 ( .A1(\REGISTERS[23][21] ), .A2(n176), .B1(
        \REGISTERS[22][21] ), .B2(n173), .ZN(n746) );
  OAI221_X1 U1193 ( .B1(n134), .B2(n1845), .C1(n131), .C2(n1813), .A(n754), 
        .ZN(n751) );
  AOI22_X1 U1194 ( .A1(\REGISTERS[7][21] ), .A2(n128), .B1(\REGISTERS[6][21] ), 
        .B2(n125), .ZN(n754) );
  OAI221_X1 U1195 ( .B1(n182), .B2(n2100), .C1(n180), .C2(n2068), .A(n728), 
        .ZN(n725) );
  AOI22_X1 U1196 ( .A1(\REGISTERS[23][22] ), .A2(n176), .B1(
        \REGISTERS[22][22] ), .B2(n173), .ZN(n728) );
  OAI221_X1 U1197 ( .B1(n134), .B2(n1844), .C1(n132), .C2(n1812), .A(n736), 
        .ZN(n733) );
  AOI22_X1 U1198 ( .A1(\REGISTERS[7][22] ), .A2(n128), .B1(\REGISTERS[6][22] ), 
        .B2(n125), .ZN(n736) );
  OAI221_X1 U1199 ( .B1(n182), .B2(n2099), .C1(n180), .C2(n2067), .A(n710), 
        .ZN(n707) );
  AOI22_X1 U1200 ( .A1(\REGISTERS[23][23] ), .A2(n176), .B1(
        \REGISTERS[22][23] ), .B2(n173), .ZN(n710) );
  OAI221_X1 U1201 ( .B1(n134), .B2(n1843), .C1(n132), .C2(n1811), .A(n718), 
        .ZN(n715) );
  AOI22_X1 U1202 ( .A1(\REGISTERS[7][23] ), .A2(n128), .B1(\REGISTERS[6][23] ), 
        .B2(n125), .ZN(n718) );
  OAI221_X1 U1203 ( .B1(n2111), .B2(n86), .C1(n2079), .C2(n83), .A(n1551), 
        .ZN(n1548) );
  AOI22_X1 U1204 ( .A1(n80), .A2(\REGISTERS[23][11] ), .B1(n77), .B2(
        \REGISTERS[22][11] ), .ZN(n1551) );
  OAI221_X1 U1205 ( .B1(n1855), .B2(n38), .C1(n1823), .C2(n35), .A(n1559), 
        .ZN(n1556) );
  AOI22_X1 U1206 ( .A1(n32), .A2(\REGISTERS[7][11] ), .B1(n29), .B2(
        \REGISTERS[6][11] ), .ZN(n1559) );
  OAI221_X1 U1207 ( .B1(n2110), .B2(n86), .C1(n2078), .C2(n83), .A(n1533), 
        .ZN(n1530) );
  AOI22_X1 U1208 ( .A1(n80), .A2(\REGISTERS[23][12] ), .B1(n77), .B2(
        \REGISTERS[22][12] ), .ZN(n1533) );
  OAI221_X1 U1209 ( .B1(n1854), .B2(n38), .C1(n1822), .C2(n35), .A(n1541), 
        .ZN(n1538) );
  AOI22_X1 U1210 ( .A1(n32), .A2(\REGISTERS[7][12] ), .B1(n29), .B2(
        \REGISTERS[6][12] ), .ZN(n1541) );
  OAI221_X1 U1211 ( .B1(n2109), .B2(n86), .C1(n2077), .C2(n83), .A(n1515), 
        .ZN(n1512) );
  AOI22_X1 U1212 ( .A1(n80), .A2(\REGISTERS[23][13] ), .B1(n77), .B2(
        \REGISTERS[22][13] ), .ZN(n1515) );
  OAI221_X1 U1213 ( .B1(n1853), .B2(n38), .C1(n1821), .C2(n35), .A(n1523), 
        .ZN(n1520) );
  AOI22_X1 U1214 ( .A1(n32), .A2(\REGISTERS[7][13] ), .B1(n29), .B2(
        \REGISTERS[6][13] ), .ZN(n1523) );
  OAI221_X1 U1215 ( .B1(n2108), .B2(n86), .C1(n2076), .C2(n83), .A(n1497), 
        .ZN(n1494) );
  AOI22_X1 U1216 ( .A1(n80), .A2(\REGISTERS[23][14] ), .B1(n77), .B2(
        \REGISTERS[22][14] ), .ZN(n1497) );
  OAI221_X1 U1217 ( .B1(n1852), .B2(n38), .C1(n1820), .C2(n35), .A(n1505), 
        .ZN(n1502) );
  AOI22_X1 U1218 ( .A1(n32), .A2(\REGISTERS[7][14] ), .B1(n29), .B2(
        \REGISTERS[6][14] ), .ZN(n1505) );
  OAI221_X1 U1219 ( .B1(n2107), .B2(n86), .C1(n2075), .C2(n83), .A(n1479), 
        .ZN(n1476) );
  AOI22_X1 U1220 ( .A1(n80), .A2(\REGISTERS[23][15] ), .B1(n77), .B2(
        \REGISTERS[22][15] ), .ZN(n1479) );
  OAI221_X1 U1221 ( .B1(n1851), .B2(n38), .C1(n1819), .C2(n35), .A(n1487), 
        .ZN(n1484) );
  AOI22_X1 U1222 ( .A1(n32), .A2(\REGISTERS[7][15] ), .B1(n29), .B2(
        \REGISTERS[6][15] ), .ZN(n1487) );
  OAI221_X1 U1223 ( .B1(n2106), .B2(n86), .C1(n2074), .C2(n83), .A(n1461), 
        .ZN(n1458) );
  AOI22_X1 U1224 ( .A1(n80), .A2(\REGISTERS[23][16] ), .B1(n77), .B2(
        \REGISTERS[22][16] ), .ZN(n1461) );
  OAI221_X1 U1225 ( .B1(n1850), .B2(n38), .C1(n1818), .C2(n35), .A(n1469), 
        .ZN(n1466) );
  AOI22_X1 U1226 ( .A1(n32), .A2(\REGISTERS[7][16] ), .B1(n29), .B2(
        \REGISTERS[6][16] ), .ZN(n1469) );
  OAI221_X1 U1227 ( .B1(n2105), .B2(n86), .C1(n2073), .C2(n83), .A(n1443), 
        .ZN(n1440) );
  AOI22_X1 U1228 ( .A1(n80), .A2(\REGISTERS[23][17] ), .B1(n77), .B2(
        \REGISTERS[22][17] ), .ZN(n1443) );
  OAI221_X1 U1229 ( .B1(n1849), .B2(n38), .C1(n1817), .C2(n35), .A(n1451), 
        .ZN(n1448) );
  AOI22_X1 U1230 ( .A1(n32), .A2(\REGISTERS[7][17] ), .B1(n29), .B2(
        \REGISTERS[6][17] ), .ZN(n1451) );
  OAI221_X1 U1231 ( .B1(n2104), .B2(n86), .C1(n2072), .C2(n83), .A(n1425), 
        .ZN(n1422) );
  AOI22_X1 U1232 ( .A1(n80), .A2(\REGISTERS[23][18] ), .B1(n77), .B2(
        \REGISTERS[22][18] ), .ZN(n1425) );
  OAI221_X1 U1233 ( .B1(n1848), .B2(n38), .C1(n1816), .C2(n35), .A(n1433), 
        .ZN(n1430) );
  AOI22_X1 U1234 ( .A1(n32), .A2(\REGISTERS[7][18] ), .B1(n29), .B2(
        \REGISTERS[6][18] ), .ZN(n1433) );
  OAI221_X1 U1235 ( .B1(n2103), .B2(n86), .C1(n2071), .C2(n83), .A(n1407), 
        .ZN(n1404) );
  AOI22_X1 U1236 ( .A1(n80), .A2(\REGISTERS[23][19] ), .B1(n77), .B2(
        \REGISTERS[22][19] ), .ZN(n1407) );
  OAI221_X1 U1237 ( .B1(n1847), .B2(n38), .C1(n1815), .C2(n35), .A(n1415), 
        .ZN(n1412) );
  AOI22_X1 U1238 ( .A1(n32), .A2(\REGISTERS[7][19] ), .B1(n29), .B2(
        \REGISTERS[6][19] ), .ZN(n1415) );
  OAI221_X1 U1239 ( .B1(n2102), .B2(n86), .C1(n2070), .C2(n83), .A(n1389), 
        .ZN(n1386) );
  AOI22_X1 U1240 ( .A1(n80), .A2(\REGISTERS[23][20] ), .B1(n77), .B2(
        \REGISTERS[22][20] ), .ZN(n1389) );
  OAI221_X1 U1241 ( .B1(n1846), .B2(n38), .C1(n1814), .C2(n35), .A(n1397), 
        .ZN(n1394) );
  AOI22_X1 U1242 ( .A1(n32), .A2(\REGISTERS[7][20] ), .B1(n29), .B2(
        \REGISTERS[6][20] ), .ZN(n1397) );
  OAI221_X1 U1243 ( .B1(n2101), .B2(n86), .C1(n2069), .C2(n83), .A(n1371), 
        .ZN(n1368) );
  AOI22_X1 U1244 ( .A1(n80), .A2(\REGISTERS[23][21] ), .B1(n77), .B2(
        \REGISTERS[22][21] ), .ZN(n1371) );
  OAI221_X1 U1245 ( .B1(n1845), .B2(n38), .C1(n1813), .C2(n35), .A(n1379), 
        .ZN(n1376) );
  AOI22_X1 U1246 ( .A1(n32), .A2(\REGISTERS[7][21] ), .B1(n29), .B2(
        \REGISTERS[6][21] ), .ZN(n1379) );
  OAI221_X1 U1247 ( .B1(n171), .B2(n2162), .C1(n168), .C2(n2130), .A(n693), 
        .ZN(n688) );
  AOI22_X1 U1248 ( .A1(\REGISTERS[27][24] ), .A2(n165), .B1(
        \REGISTERS[26][24] ), .B2(n162), .ZN(n693) );
  OAI221_X1 U1249 ( .B1(n171), .B2(n2161), .C1(n168), .C2(n2129), .A(n675), 
        .ZN(n670) );
  AOI22_X1 U1250 ( .A1(\REGISTERS[27][25] ), .A2(n165), .B1(
        \REGISTERS[26][25] ), .B2(n162), .ZN(n675) );
  OAI221_X1 U1251 ( .B1(n171), .B2(n2160), .C1(n168), .C2(n2128), .A(n657), 
        .ZN(n652) );
  AOI22_X1 U1252 ( .A1(\REGISTERS[27][26] ), .A2(n165), .B1(
        \REGISTERS[26][26] ), .B2(n162), .ZN(n657) );
  OAI221_X1 U1253 ( .B1(n171), .B2(n2159), .C1(n168), .C2(n2127), .A(n639), 
        .ZN(n634) );
  AOI22_X1 U1254 ( .A1(\REGISTERS[27][27] ), .A2(n165), .B1(
        \REGISTERS[26][27] ), .B2(n162), .ZN(n639) );
  OAI221_X1 U1255 ( .B1(n171), .B2(n2158), .C1(n168), .C2(n2126), .A(n621), 
        .ZN(n616) );
  AOI22_X1 U1256 ( .A1(\REGISTERS[27][28] ), .A2(n165), .B1(
        \REGISTERS[26][28] ), .B2(n162), .ZN(n621) );
  OAI221_X1 U1257 ( .B1(n171), .B2(n2157), .C1(n168), .C2(n2125), .A(n603), 
        .ZN(n598) );
  AOI22_X1 U1258 ( .A1(\REGISTERS[27][29] ), .A2(n165), .B1(
        \REGISTERS[26][29] ), .B2(n162), .ZN(n603) );
  OAI221_X1 U1259 ( .B1(n171), .B2(n2156), .C1(n168), .C2(n2124), .A(n585), 
        .ZN(n580) );
  AOI22_X1 U1260 ( .A1(\REGISTERS[27][30] ), .A2(n165), .B1(
        \REGISTERS[26][30] ), .B2(n162), .ZN(n585) );
  OAI221_X1 U1261 ( .B1(n171), .B2(n2155), .C1(n168), .C2(n2123), .A(n545), 
        .ZN(n530) );
  AOI22_X1 U1262 ( .A1(\REGISTERS[27][31] ), .A2(n165), .B1(
        \REGISTERS[26][31] ), .B2(n162), .ZN(n545) );
  OAI221_X1 U1263 ( .B1(n123), .B2(n1906), .C1(n120), .C2(n1874), .A(n701), 
        .ZN(n696) );
  AOI22_X1 U1264 ( .A1(\REGISTERS[11][24] ), .A2(n117), .B1(
        \REGISTERS[10][24] ), .B2(n114), .ZN(n701) );
  OAI221_X1 U1265 ( .B1(n123), .B2(n1905), .C1(n120), .C2(n1873), .A(n683), 
        .ZN(n678) );
  AOI22_X1 U1266 ( .A1(\REGISTERS[11][25] ), .A2(n117), .B1(
        \REGISTERS[10][25] ), .B2(n114), .ZN(n683) );
  OAI221_X1 U1267 ( .B1(n123), .B2(n1904), .C1(n120), .C2(n1872), .A(n665), 
        .ZN(n660) );
  AOI22_X1 U1268 ( .A1(\REGISTERS[11][26] ), .A2(n117), .B1(
        \REGISTERS[10][26] ), .B2(n114), .ZN(n665) );
  OAI221_X1 U1269 ( .B1(n123), .B2(n1903), .C1(n120), .C2(n1871), .A(n647), 
        .ZN(n642) );
  AOI22_X1 U1270 ( .A1(\REGISTERS[11][27] ), .A2(n117), .B1(
        \REGISTERS[10][27] ), .B2(n114), .ZN(n647) );
  OAI221_X1 U1271 ( .B1(n123), .B2(n1902), .C1(n120), .C2(n1870), .A(n629), 
        .ZN(n624) );
  AOI22_X1 U1272 ( .A1(\REGISTERS[11][28] ), .A2(n117), .B1(
        \REGISTERS[10][28] ), .B2(n114), .ZN(n629) );
  OAI221_X1 U1273 ( .B1(n123), .B2(n1901), .C1(n120), .C2(n1869), .A(n611), 
        .ZN(n606) );
  AOI22_X1 U1274 ( .A1(\REGISTERS[11][29] ), .A2(n117), .B1(
        \REGISTERS[10][29] ), .B2(n114), .ZN(n611) );
  OAI221_X1 U1275 ( .B1(n123), .B2(n1900), .C1(n120), .C2(n1868), .A(n593), 
        .ZN(n588) );
  AOI22_X1 U1276 ( .A1(\REGISTERS[11][30] ), .A2(n117), .B1(
        \REGISTERS[10][30] ), .B2(n114), .ZN(n593) );
  OAI221_X1 U1277 ( .B1(n123), .B2(n1899), .C1(n120), .C2(n1867), .A(n569), 
        .ZN(n554) );
  AOI22_X1 U1278 ( .A1(\REGISTERS[11][31] ), .A2(n117), .B1(
        \REGISTERS[10][31] ), .B2(n114), .ZN(n569) );
  OAI221_X1 U1279 ( .B1(n2186), .B2(n73), .C1(n2154), .C2(n70), .A(n1757), 
        .ZN(n1745) );
  AOI22_X1 U1280 ( .A1(n67), .A2(\REGISTERS[27][0] ), .B1(n64), .B2(
        \REGISTERS[26][0] ), .ZN(n1757) );
  OAI221_X1 U1281 ( .B1(n1930), .B2(n25), .C1(n1898), .C2(n22), .A(n1771), 
        .ZN(n1763) );
  AOI22_X1 U1282 ( .A1(n19), .A2(\REGISTERS[11][0] ), .B1(n16), .B2(
        \REGISTERS[10][0] ), .ZN(n1771) );
  OAI221_X1 U1283 ( .B1(n2185), .B2(n73), .C1(n2153), .C2(n70), .A(n1732), 
        .ZN(n1727) );
  AOI22_X1 U1284 ( .A1(n67), .A2(\REGISTERS[27][1] ), .B1(n64), .B2(
        \REGISTERS[26][1] ), .ZN(n1732) );
  OAI221_X1 U1285 ( .B1(n1929), .B2(n25), .C1(n1897), .C2(n22), .A(n1740), 
        .ZN(n1735) );
  AOI22_X1 U1286 ( .A1(n19), .A2(\REGISTERS[11][1] ), .B1(n16), .B2(
        \REGISTERS[10][1] ), .ZN(n1740) );
  OAI221_X1 U1287 ( .B1(n2184), .B2(n73), .C1(n2152), .C2(n70), .A(n1714), 
        .ZN(n1709) );
  AOI22_X1 U1288 ( .A1(n67), .A2(\REGISTERS[27][2] ), .B1(n64), .B2(
        \REGISTERS[26][2] ), .ZN(n1714) );
  OAI221_X1 U1289 ( .B1(n1928), .B2(n25), .C1(n1896), .C2(n22), .A(n1722), 
        .ZN(n1717) );
  AOI22_X1 U1290 ( .A1(n19), .A2(\REGISTERS[11][2] ), .B1(n16), .B2(
        \REGISTERS[10][2] ), .ZN(n1722) );
  OAI221_X1 U1291 ( .B1(n2183), .B2(n73), .C1(n2151), .C2(n70), .A(n1696), 
        .ZN(n1691) );
  AOI22_X1 U1292 ( .A1(n67), .A2(\REGISTERS[27][3] ), .B1(n64), .B2(
        \REGISTERS[26][3] ), .ZN(n1696) );
  OAI221_X1 U1293 ( .B1(n1927), .B2(n25), .C1(n1895), .C2(n22), .A(n1704), 
        .ZN(n1699) );
  AOI22_X1 U1294 ( .A1(n19), .A2(\REGISTERS[11][3] ), .B1(n16), .B2(
        \REGISTERS[10][3] ), .ZN(n1704) );
  OAI221_X1 U1295 ( .B1(n2182), .B2(n73), .C1(n2150), .C2(n70), .A(n1678), 
        .ZN(n1673) );
  AOI22_X1 U1296 ( .A1(n67), .A2(\REGISTERS[27][4] ), .B1(n64), .B2(
        \REGISTERS[26][4] ), .ZN(n1678) );
  OAI221_X1 U1297 ( .B1(n1926), .B2(n25), .C1(n1894), .C2(n22), .A(n1686), 
        .ZN(n1681) );
  AOI22_X1 U1298 ( .A1(n19), .A2(\REGISTERS[11][4] ), .B1(n16), .B2(
        \REGISTERS[10][4] ), .ZN(n1686) );
  OAI221_X1 U1299 ( .B1(n2181), .B2(n73), .C1(n2149), .C2(n70), .A(n1660), 
        .ZN(n1655) );
  AOI22_X1 U1300 ( .A1(n67), .A2(\REGISTERS[27][5] ), .B1(n64), .B2(
        \REGISTERS[26][5] ), .ZN(n1660) );
  OAI221_X1 U1301 ( .B1(n1925), .B2(n25), .C1(n1893), .C2(n22), .A(n1668), 
        .ZN(n1663) );
  AOI22_X1 U1302 ( .A1(n19), .A2(\REGISTERS[11][5] ), .B1(n16), .B2(
        \REGISTERS[10][5] ), .ZN(n1668) );
  OAI221_X1 U1303 ( .B1(n2180), .B2(n73), .C1(n2148), .C2(n70), .A(n1642), 
        .ZN(n1637) );
  AOI22_X1 U1304 ( .A1(n67), .A2(\REGISTERS[27][6] ), .B1(n64), .B2(
        \REGISTERS[26][6] ), .ZN(n1642) );
  OAI221_X1 U1305 ( .B1(n1924), .B2(n25), .C1(n1892), .C2(n22), .A(n1650), 
        .ZN(n1645) );
  AOI22_X1 U1306 ( .A1(n19), .A2(\REGISTERS[11][6] ), .B1(n16), .B2(
        \REGISTERS[10][6] ), .ZN(n1650) );
  OAI221_X1 U1307 ( .B1(n2179), .B2(n73), .C1(n2147), .C2(n70), .A(n1624), 
        .ZN(n1619) );
  AOI22_X1 U1308 ( .A1(n67), .A2(\REGISTERS[27][7] ), .B1(n64), .B2(
        \REGISTERS[26][7] ), .ZN(n1624) );
  OAI221_X1 U1309 ( .B1(n1923), .B2(n25), .C1(n1891), .C2(n22), .A(n1632), 
        .ZN(n1627) );
  AOI22_X1 U1310 ( .A1(n19), .A2(\REGISTERS[11][7] ), .B1(n16), .B2(
        \REGISTERS[10][7] ), .ZN(n1632) );
  OAI221_X1 U1311 ( .B1(n2178), .B2(n73), .C1(n2146), .C2(n70), .A(n1606), 
        .ZN(n1601) );
  AOI22_X1 U1312 ( .A1(n67), .A2(\REGISTERS[27][8] ), .B1(n64), .B2(
        \REGISTERS[26][8] ), .ZN(n1606) );
  OAI221_X1 U1313 ( .B1(n1922), .B2(n25), .C1(n1890), .C2(n22), .A(n1614), 
        .ZN(n1609) );
  AOI22_X1 U1314 ( .A1(n19), .A2(\REGISTERS[11][8] ), .B1(n16), .B2(
        \REGISTERS[10][8] ), .ZN(n1614) );
  OAI221_X1 U1315 ( .B1(n2177), .B2(n73), .C1(n2145), .C2(n70), .A(n1588), 
        .ZN(n1583) );
  AOI22_X1 U1316 ( .A1(n67), .A2(\REGISTERS[27][9] ), .B1(n64), .B2(
        \REGISTERS[26][9] ), .ZN(n1588) );
  OAI221_X1 U1317 ( .B1(n1921), .B2(n25), .C1(n1889), .C2(n22), .A(n1596), 
        .ZN(n1591) );
  AOI22_X1 U1318 ( .A1(n19), .A2(\REGISTERS[11][9] ), .B1(n16), .B2(
        \REGISTERS[10][9] ), .ZN(n1596) );
  OAI221_X1 U1319 ( .B1(n2176), .B2(n73), .C1(n2144), .C2(n70), .A(n1570), 
        .ZN(n1565) );
  AOI22_X1 U1320 ( .A1(n67), .A2(\REGISTERS[27][10] ), .B1(n64), .B2(
        \REGISTERS[26][10] ), .ZN(n1570) );
  OAI221_X1 U1321 ( .B1(n1920), .B2(n25), .C1(n1888), .C2(n22), .A(n1578), 
        .ZN(n1573) );
  AOI22_X1 U1322 ( .A1(n19), .A2(\REGISTERS[11][10] ), .B1(n16), .B2(
        \REGISTERS[10][10] ), .ZN(n1578) );
  OAI221_X1 U1323 ( .B1(n159), .B2(n2226), .C1(n156), .C2(n2194), .A(n694), 
        .ZN(n687) );
  AOI22_X1 U1324 ( .A1(\REGISTERS[29][24] ), .A2(n153), .B1(
        \REGISTERS[28][24] ), .B2(n150), .ZN(n694) );
  OAI221_X1 U1325 ( .B1(n159), .B2(n2225), .C1(n156), .C2(n2193), .A(n676), 
        .ZN(n669) );
  AOI22_X1 U1326 ( .A1(\REGISTERS[29][25] ), .A2(n153), .B1(
        \REGISTERS[28][25] ), .B2(n150), .ZN(n676) );
  OAI221_X1 U1327 ( .B1(n159), .B2(n2224), .C1(n156), .C2(n2192), .A(n658), 
        .ZN(n651) );
  AOI22_X1 U1328 ( .A1(\REGISTERS[29][26] ), .A2(n153), .B1(
        \REGISTERS[28][26] ), .B2(n150), .ZN(n658) );
  OAI221_X1 U1329 ( .B1(n159), .B2(n2223), .C1(n156), .C2(n2191), .A(n640), 
        .ZN(n633) );
  AOI22_X1 U1330 ( .A1(\REGISTERS[29][27] ), .A2(n153), .B1(
        \REGISTERS[28][27] ), .B2(n150), .ZN(n640) );
  OAI221_X1 U1331 ( .B1(n159), .B2(n2222), .C1(n156), .C2(n2190), .A(n622), 
        .ZN(n615) );
  AOI22_X1 U1332 ( .A1(\REGISTERS[29][28] ), .A2(n153), .B1(
        \REGISTERS[28][28] ), .B2(n150), .ZN(n622) );
  OAI221_X1 U1333 ( .B1(n159), .B2(n2221), .C1(n156), .C2(n2189), .A(n604), 
        .ZN(n597) );
  AOI22_X1 U1334 ( .A1(\REGISTERS[29][29] ), .A2(n153), .B1(
        \REGISTERS[28][29] ), .B2(n150), .ZN(n604) );
  OAI221_X1 U1335 ( .B1(n159), .B2(n2220), .C1(n156), .C2(n2188), .A(n586), 
        .ZN(n579) );
  AOI22_X1 U1336 ( .A1(\REGISTERS[29][30] ), .A2(n153), .B1(
        \REGISTERS[28][30] ), .B2(n150), .ZN(n586) );
  OAI221_X1 U1337 ( .B1(n159), .B2(n2219), .C1(n156), .C2(n2187), .A(n550), 
        .ZN(n529) );
  AOI22_X1 U1338 ( .A1(\REGISTERS[29][31] ), .A2(n153), .B1(
        \REGISTERS[28][31] ), .B2(n150), .ZN(n550) );
  OAI221_X1 U1339 ( .B1(n2164), .B2(n75), .C1(n2132), .C2(n72), .A(n1354), 
        .ZN(n1349) );
  AOI22_X1 U1340 ( .A1(n69), .A2(\REGISTERS[27][22] ), .B1(n66), .B2(
        \REGISTERS[26][22] ), .ZN(n1354) );
  OAI221_X1 U1341 ( .B1(n1908), .B2(n27), .C1(n1876), .C2(n24), .A(n1362), 
        .ZN(n1357) );
  AOI22_X1 U1342 ( .A1(n21), .A2(\REGISTERS[11][22] ), .B1(n18), .B2(
        \REGISTERS[10][22] ), .ZN(n1362) );
  OAI221_X1 U1343 ( .B1(n2163), .B2(n75), .C1(n2131), .C2(n72), .A(n1336), 
        .ZN(n1331) );
  AOI22_X1 U1344 ( .A1(n69), .A2(\REGISTERS[27][23] ), .B1(n66), .B2(
        \REGISTERS[26][23] ), .ZN(n1336) );
  OAI221_X1 U1345 ( .B1(n1907), .B2(n27), .C1(n1875), .C2(n24), .A(n1344), 
        .ZN(n1339) );
  AOI22_X1 U1346 ( .A1(n21), .A2(\REGISTERS[11][23] ), .B1(n18), .B2(
        \REGISTERS[10][23] ), .ZN(n1344) );
  OAI221_X1 U1347 ( .B1(n2162), .B2(n75), .C1(n2130), .C2(n72), .A(n1318), 
        .ZN(n1313) );
  AOI22_X1 U1348 ( .A1(n69), .A2(\REGISTERS[27][24] ), .B1(n66), .B2(
        \REGISTERS[26][24] ), .ZN(n1318) );
  OAI221_X1 U1349 ( .B1(n1906), .B2(n27), .C1(n1874), .C2(n24), .A(n1326), 
        .ZN(n1321) );
  AOI22_X1 U1350 ( .A1(n21), .A2(\REGISTERS[11][24] ), .B1(n18), .B2(
        \REGISTERS[10][24] ), .ZN(n1326) );
  OAI221_X1 U1351 ( .B1(n2161), .B2(n75), .C1(n2129), .C2(n72), .A(n1300), 
        .ZN(n1295) );
  AOI22_X1 U1352 ( .A1(n69), .A2(\REGISTERS[27][25] ), .B1(n66), .B2(
        \REGISTERS[26][25] ), .ZN(n1300) );
  OAI221_X1 U1353 ( .B1(n1905), .B2(n27), .C1(n1873), .C2(n24), .A(n1308), 
        .ZN(n1303) );
  AOI22_X1 U1354 ( .A1(n21), .A2(\REGISTERS[11][25] ), .B1(n18), .B2(
        \REGISTERS[10][25] ), .ZN(n1308) );
  OAI221_X1 U1355 ( .B1(n2160), .B2(n75), .C1(n2128), .C2(n72), .A(n1282), 
        .ZN(n1277) );
  AOI22_X1 U1356 ( .A1(n69), .A2(\REGISTERS[27][26] ), .B1(n66), .B2(
        \REGISTERS[26][26] ), .ZN(n1282) );
  OAI221_X1 U1357 ( .B1(n1904), .B2(n27), .C1(n1872), .C2(n24), .A(n1290), 
        .ZN(n1285) );
  AOI22_X1 U1358 ( .A1(n21), .A2(\REGISTERS[11][26] ), .B1(n18), .B2(
        \REGISTERS[10][26] ), .ZN(n1290) );
  OAI221_X1 U1359 ( .B1(n2159), .B2(n75), .C1(n2127), .C2(n72), .A(n1264), 
        .ZN(n1259) );
  AOI22_X1 U1360 ( .A1(n69), .A2(\REGISTERS[27][27] ), .B1(n66), .B2(
        \REGISTERS[26][27] ), .ZN(n1264) );
  OAI221_X1 U1361 ( .B1(n1903), .B2(n27), .C1(n1871), .C2(n24), .A(n1272), 
        .ZN(n1267) );
  AOI22_X1 U1362 ( .A1(n21), .A2(\REGISTERS[11][27] ), .B1(n18), .B2(
        \REGISTERS[10][27] ), .ZN(n1272) );
  OAI221_X1 U1363 ( .B1(n2158), .B2(n75), .C1(n2126), .C2(n72), .A(n1246), 
        .ZN(n1241) );
  AOI22_X1 U1364 ( .A1(n69), .A2(\REGISTERS[27][28] ), .B1(n66), .B2(
        \REGISTERS[26][28] ), .ZN(n1246) );
  OAI221_X1 U1365 ( .B1(n1902), .B2(n27), .C1(n1870), .C2(n24), .A(n1254), 
        .ZN(n1249) );
  AOI22_X1 U1366 ( .A1(n21), .A2(\REGISTERS[11][28] ), .B1(n18), .B2(
        \REGISTERS[10][28] ), .ZN(n1254) );
  OAI221_X1 U1367 ( .B1(n2157), .B2(n75), .C1(n2125), .C2(n72), .A(n1228), 
        .ZN(n1223) );
  AOI22_X1 U1368 ( .A1(n69), .A2(\REGISTERS[27][29] ), .B1(n66), .B2(
        \REGISTERS[26][29] ), .ZN(n1228) );
  OAI221_X1 U1369 ( .B1(n1901), .B2(n27), .C1(n1869), .C2(n24), .A(n1236), 
        .ZN(n1231) );
  AOI22_X1 U1370 ( .A1(n21), .A2(\REGISTERS[11][29] ), .B1(n18), .B2(
        \REGISTERS[10][29] ), .ZN(n1236) );
  OAI221_X1 U1371 ( .B1(n2156), .B2(n75), .C1(n2124), .C2(n72), .A(n1210), 
        .ZN(n1205) );
  AOI22_X1 U1372 ( .A1(n69), .A2(\REGISTERS[27][30] ), .B1(n66), .B2(
        \REGISTERS[26][30] ), .ZN(n1210) );
  OAI221_X1 U1373 ( .B1(n1900), .B2(n27), .C1(n1868), .C2(n24), .A(n1218), 
        .ZN(n1213) );
  AOI22_X1 U1374 ( .A1(n21), .A2(\REGISTERS[11][30] ), .B1(n18), .B2(
        \REGISTERS[10][30] ), .ZN(n1218) );
  OAI221_X1 U1375 ( .B1(n2155), .B2(n75), .C1(n2123), .C2(n72), .A(n1170), 
        .ZN(n1155) );
  AOI22_X1 U1376 ( .A1(n69), .A2(\REGISTERS[27][31] ), .B1(n66), .B2(
        \REGISTERS[26][31] ), .ZN(n1170) );
  OAI221_X1 U1377 ( .B1(n1899), .B2(n27), .C1(n1867), .C2(n24), .A(n1194), 
        .ZN(n1179) );
  AOI22_X1 U1378 ( .A1(n21), .A2(\REGISTERS[11][31] ), .B1(n18), .B2(
        \REGISTERS[10][31] ), .ZN(n1194) );
  OAI221_X1 U1379 ( .B1(n2250), .B2(n61), .C1(n2218), .C2(n58), .A(n1760), 
        .ZN(n1744) );
  AOI22_X1 U1380 ( .A1(n55), .A2(\REGISTERS[29][0] ), .B1(n52), .B2(
        \REGISTERS[28][0] ), .ZN(n1760) );
  OAI221_X1 U1381 ( .B1(n2249), .B2(n61), .C1(n2217), .C2(n58), .A(n1733), 
        .ZN(n1726) );
  AOI22_X1 U1382 ( .A1(n55), .A2(\REGISTERS[29][1] ), .B1(n52), .B2(
        \REGISTERS[28][1] ), .ZN(n1733) );
  OAI221_X1 U1383 ( .B1(n2248), .B2(n61), .C1(n2216), .C2(n58), .A(n1715), 
        .ZN(n1708) );
  AOI22_X1 U1384 ( .A1(n55), .A2(\REGISTERS[29][2] ), .B1(n52), .B2(
        \REGISTERS[28][2] ), .ZN(n1715) );
  OAI221_X1 U1385 ( .B1(n2247), .B2(n61), .C1(n2215), .C2(n58), .A(n1697), 
        .ZN(n1690) );
  AOI22_X1 U1386 ( .A1(n55), .A2(\REGISTERS[29][3] ), .B1(n52), .B2(
        \REGISTERS[28][3] ), .ZN(n1697) );
  OAI221_X1 U1387 ( .B1(n2246), .B2(n61), .C1(n2214), .C2(n58), .A(n1679), 
        .ZN(n1672) );
  AOI22_X1 U1388 ( .A1(n55), .A2(\REGISTERS[29][4] ), .B1(n52), .B2(
        \REGISTERS[28][4] ), .ZN(n1679) );
  OAI221_X1 U1389 ( .B1(n2245), .B2(n61), .C1(n2213), .C2(n58), .A(n1661), 
        .ZN(n1654) );
  AOI22_X1 U1390 ( .A1(n55), .A2(\REGISTERS[29][5] ), .B1(n52), .B2(
        \REGISTERS[28][5] ), .ZN(n1661) );
  OAI221_X1 U1391 ( .B1(n2244), .B2(n61), .C1(n2212), .C2(n58), .A(n1643), 
        .ZN(n1636) );
  AOI22_X1 U1392 ( .A1(n55), .A2(\REGISTERS[29][6] ), .B1(n52), .B2(
        \REGISTERS[28][6] ), .ZN(n1643) );
  OAI221_X1 U1393 ( .B1(n2243), .B2(n61), .C1(n2211), .C2(n58), .A(n1625), 
        .ZN(n1618) );
  AOI22_X1 U1394 ( .A1(n55), .A2(\REGISTERS[29][7] ), .B1(n52), .B2(
        \REGISTERS[28][7] ), .ZN(n1625) );
  OAI221_X1 U1395 ( .B1(n2242), .B2(n61), .C1(n2210), .C2(n58), .A(n1607), 
        .ZN(n1600) );
  AOI22_X1 U1396 ( .A1(n55), .A2(\REGISTERS[29][8] ), .B1(n52), .B2(
        \REGISTERS[28][8] ), .ZN(n1607) );
  OAI221_X1 U1397 ( .B1(n2241), .B2(n61), .C1(n2209), .C2(n58), .A(n1589), 
        .ZN(n1582) );
  AOI22_X1 U1398 ( .A1(n55), .A2(\REGISTERS[29][9] ), .B1(n52), .B2(
        \REGISTERS[28][9] ), .ZN(n1589) );
  OAI221_X1 U1399 ( .B1(n2240), .B2(n61), .C1(n2208), .C2(n58), .A(n1571), 
        .ZN(n1564) );
  AOI22_X1 U1400 ( .A1(n55), .A2(\REGISTERS[29][10] ), .B1(n52), .B2(
        \REGISTERS[28][10] ), .ZN(n1571) );
  OAI221_X1 U1401 ( .B1(n2228), .B2(n63), .C1(n2196), .C2(n60), .A(n1355), 
        .ZN(n1348) );
  AOI22_X1 U1402 ( .A1(n57), .A2(\REGISTERS[29][22] ), .B1(n54), .B2(
        \REGISTERS[28][22] ), .ZN(n1355) );
  OAI221_X1 U1403 ( .B1(n2227), .B2(n63), .C1(n2195), .C2(n60), .A(n1337), 
        .ZN(n1330) );
  AOI22_X1 U1404 ( .A1(n57), .A2(\REGISTERS[29][23] ), .B1(n54), .B2(
        \REGISTERS[28][23] ), .ZN(n1337) );
  OAI221_X1 U1405 ( .B1(n2226), .B2(n63), .C1(n2194), .C2(n60), .A(n1319), 
        .ZN(n1312) );
  AOI22_X1 U1406 ( .A1(n57), .A2(\REGISTERS[29][24] ), .B1(n54), .B2(
        \REGISTERS[28][24] ), .ZN(n1319) );
  OAI221_X1 U1407 ( .B1(n2225), .B2(n63), .C1(n2193), .C2(n60), .A(n1301), 
        .ZN(n1294) );
  AOI22_X1 U1408 ( .A1(n57), .A2(\REGISTERS[29][25] ), .B1(n54), .B2(
        \REGISTERS[28][25] ), .ZN(n1301) );
  OAI221_X1 U1409 ( .B1(n2224), .B2(n63), .C1(n2192), .C2(n60), .A(n1283), 
        .ZN(n1276) );
  AOI22_X1 U1410 ( .A1(n57), .A2(\REGISTERS[29][26] ), .B1(n54), .B2(
        \REGISTERS[28][26] ), .ZN(n1283) );
  OAI221_X1 U1411 ( .B1(n2223), .B2(n63), .C1(n2191), .C2(n60), .A(n1265), 
        .ZN(n1258) );
  AOI22_X1 U1412 ( .A1(n57), .A2(\REGISTERS[29][27] ), .B1(n54), .B2(
        \REGISTERS[28][27] ), .ZN(n1265) );
  OAI221_X1 U1413 ( .B1(n2222), .B2(n63), .C1(n2190), .C2(n60), .A(n1247), 
        .ZN(n1240) );
  AOI22_X1 U1414 ( .A1(n57), .A2(\REGISTERS[29][28] ), .B1(n54), .B2(
        \REGISTERS[28][28] ), .ZN(n1247) );
  OAI221_X1 U1415 ( .B1(n2221), .B2(n63), .C1(n2189), .C2(n60), .A(n1229), 
        .ZN(n1222) );
  AOI22_X1 U1416 ( .A1(n57), .A2(\REGISTERS[29][29] ), .B1(n54), .B2(
        \REGISTERS[28][29] ), .ZN(n1229) );
  OAI221_X1 U1417 ( .B1(n2220), .B2(n63), .C1(n2188), .C2(n60), .A(n1211), 
        .ZN(n1204) );
  AOI22_X1 U1418 ( .A1(n57), .A2(\REGISTERS[29][30] ), .B1(n54), .B2(
        \REGISTERS[28][30] ), .ZN(n1211) );
  OAI221_X1 U1419 ( .B1(n2219), .B2(n63), .C1(n2187), .C2(n60), .A(n1175), 
        .ZN(n1154) );
  AOI22_X1 U1420 ( .A1(n57), .A2(\REGISTERS[29][31] ), .B1(n54), .B2(
        \REGISTERS[28][31] ), .ZN(n1175) );
  OAI221_X1 U1421 ( .B1(n169), .B2(n2186), .C1(n166), .C2(n2154), .A(n1132), 
        .ZN(n1120) );
  AOI22_X1 U1422 ( .A1(\REGISTERS[27][0] ), .A2(n163), .B1(\REGISTERS[26][0] ), 
        .B2(n160), .ZN(n1132) );
  OAI221_X1 U1423 ( .B1(n121), .B2(n1930), .C1(n118), .C2(n1898), .A(n1146), 
        .ZN(n1138) );
  AOI22_X1 U1424 ( .A1(\REGISTERS[11][0] ), .A2(n115), .B1(\REGISTERS[10][0] ), 
        .B2(n112), .ZN(n1146) );
  OAI221_X1 U1425 ( .B1(n169), .B2(n2185), .C1(n166), .C2(n2153), .A(n1107), 
        .ZN(n1102) );
  AOI22_X1 U1426 ( .A1(\REGISTERS[27][1] ), .A2(n163), .B1(\REGISTERS[26][1] ), 
        .B2(n160), .ZN(n1107) );
  OAI221_X1 U1427 ( .B1(n121), .B2(n1929), .C1(n118), .C2(n1897), .A(n1115), 
        .ZN(n1110) );
  AOI22_X1 U1428 ( .A1(\REGISTERS[11][1] ), .A2(n115), .B1(\REGISTERS[10][1] ), 
        .B2(n112), .ZN(n1115) );
  OAI221_X1 U1429 ( .B1(n169), .B2(n2184), .C1(n166), .C2(n2152), .A(n1089), 
        .ZN(n1084) );
  AOI22_X1 U1430 ( .A1(\REGISTERS[27][2] ), .A2(n163), .B1(\REGISTERS[26][2] ), 
        .B2(n160), .ZN(n1089) );
  OAI221_X1 U1431 ( .B1(n121), .B2(n1928), .C1(n118), .C2(n1896), .A(n1097), 
        .ZN(n1092) );
  AOI22_X1 U1432 ( .A1(\REGISTERS[11][2] ), .A2(n115), .B1(\REGISTERS[10][2] ), 
        .B2(n112), .ZN(n1097) );
  OAI221_X1 U1433 ( .B1(n169), .B2(n2183), .C1(n166), .C2(n2151), .A(n1071), 
        .ZN(n1066) );
  AOI22_X1 U1434 ( .A1(\REGISTERS[27][3] ), .A2(n163), .B1(\REGISTERS[26][3] ), 
        .B2(n160), .ZN(n1071) );
  OAI221_X1 U1435 ( .B1(n121), .B2(n1927), .C1(n118), .C2(n1895), .A(n1079), 
        .ZN(n1074) );
  AOI22_X1 U1436 ( .A1(\REGISTERS[11][3] ), .A2(n115), .B1(\REGISTERS[10][3] ), 
        .B2(n112), .ZN(n1079) );
  OAI221_X1 U1437 ( .B1(n169), .B2(n2182), .C1(n166), .C2(n2150), .A(n1053), 
        .ZN(n1048) );
  AOI22_X1 U1438 ( .A1(\REGISTERS[27][4] ), .A2(n163), .B1(\REGISTERS[26][4] ), 
        .B2(n160), .ZN(n1053) );
  OAI221_X1 U1439 ( .B1(n121), .B2(n1926), .C1(n118), .C2(n1894), .A(n1061), 
        .ZN(n1056) );
  AOI22_X1 U1440 ( .A1(\REGISTERS[11][4] ), .A2(n115), .B1(\REGISTERS[10][4] ), 
        .B2(n112), .ZN(n1061) );
  OAI221_X1 U1441 ( .B1(n169), .B2(n2181), .C1(n166), .C2(n2149), .A(n1035), 
        .ZN(n1030) );
  AOI22_X1 U1442 ( .A1(\REGISTERS[27][5] ), .A2(n163), .B1(\REGISTERS[26][5] ), 
        .B2(n160), .ZN(n1035) );
  OAI221_X1 U1443 ( .B1(n121), .B2(n1925), .C1(n118), .C2(n1893), .A(n1043), 
        .ZN(n1038) );
  AOI22_X1 U1444 ( .A1(\REGISTERS[11][5] ), .A2(n115), .B1(\REGISTERS[10][5] ), 
        .B2(n112), .ZN(n1043) );
  OAI221_X1 U1445 ( .B1(n169), .B2(n2180), .C1(n166), .C2(n2148), .A(n1017), 
        .ZN(n1012) );
  AOI22_X1 U1446 ( .A1(\REGISTERS[27][6] ), .A2(n163), .B1(\REGISTERS[26][6] ), 
        .B2(n160), .ZN(n1017) );
  OAI221_X1 U1447 ( .B1(n121), .B2(n1924), .C1(n118), .C2(n1892), .A(n1025), 
        .ZN(n1020) );
  AOI22_X1 U1448 ( .A1(\REGISTERS[11][6] ), .A2(n115), .B1(\REGISTERS[10][6] ), 
        .B2(n112), .ZN(n1025) );
  OAI221_X1 U1449 ( .B1(n169), .B2(n2179), .C1(n166), .C2(n2147), .A(n999), 
        .ZN(n994) );
  AOI22_X1 U1450 ( .A1(\REGISTERS[27][7] ), .A2(n163), .B1(\REGISTERS[26][7] ), 
        .B2(n160), .ZN(n999) );
  OAI221_X1 U1451 ( .B1(n121), .B2(n1923), .C1(n118), .C2(n1891), .A(n1007), 
        .ZN(n1002) );
  AOI22_X1 U1452 ( .A1(\REGISTERS[11][7] ), .A2(n115), .B1(\REGISTERS[10][7] ), 
        .B2(n112), .ZN(n1007) );
  OAI221_X1 U1453 ( .B1(n169), .B2(n2178), .C1(n166), .C2(n2146), .A(n981), 
        .ZN(n976) );
  AOI22_X1 U1454 ( .A1(\REGISTERS[27][8] ), .A2(n163), .B1(\REGISTERS[26][8] ), 
        .B2(n160), .ZN(n981) );
  OAI221_X1 U1455 ( .B1(n121), .B2(n1922), .C1(n118), .C2(n1890), .A(n989), 
        .ZN(n984) );
  AOI22_X1 U1456 ( .A1(\REGISTERS[11][8] ), .A2(n115), .B1(\REGISTERS[10][8] ), 
        .B2(n112), .ZN(n989) );
  OAI221_X1 U1457 ( .B1(n169), .B2(n2177), .C1(n166), .C2(n2145), .A(n963), 
        .ZN(n958) );
  AOI22_X1 U1458 ( .A1(\REGISTERS[27][9] ), .A2(n163), .B1(\REGISTERS[26][9] ), 
        .B2(n160), .ZN(n963) );
  OAI221_X1 U1459 ( .B1(n121), .B2(n1921), .C1(n118), .C2(n1889), .A(n971), 
        .ZN(n966) );
  AOI22_X1 U1460 ( .A1(\REGISTERS[11][9] ), .A2(n115), .B1(\REGISTERS[10][9] ), 
        .B2(n112), .ZN(n971) );
  OAI221_X1 U1461 ( .B1(n169), .B2(n2176), .C1(n166), .C2(n2144), .A(n945), 
        .ZN(n940) );
  AOI22_X1 U1462 ( .A1(\REGISTERS[27][10] ), .A2(n163), .B1(
        \REGISTERS[26][10] ), .B2(n160), .ZN(n945) );
  OAI221_X1 U1463 ( .B1(n121), .B2(n1920), .C1(n118), .C2(n1888), .A(n953), 
        .ZN(n948) );
  AOI22_X1 U1464 ( .A1(\REGISTERS[11][10] ), .A2(n115), .B1(
        \REGISTERS[10][10] ), .B2(n112), .ZN(n953) );
  OAI221_X1 U1465 ( .B1(n169), .B2(n2175), .C1(n167), .C2(n2143), .A(n927), 
        .ZN(n922) );
  AOI22_X1 U1466 ( .A1(\REGISTERS[27][11] ), .A2(n163), .B1(
        \REGISTERS[26][11] ), .B2(n160), .ZN(n927) );
  OAI221_X1 U1467 ( .B1(n121), .B2(n1919), .C1(n119), .C2(n1887), .A(n935), 
        .ZN(n930) );
  AOI22_X1 U1468 ( .A1(\REGISTERS[11][11] ), .A2(n115), .B1(
        \REGISTERS[10][11] ), .B2(n112), .ZN(n935) );
  OAI221_X1 U1469 ( .B1(n170), .B2(n2174), .C1(n167), .C2(n2142), .A(n909), 
        .ZN(n904) );
  AOI22_X1 U1470 ( .A1(\REGISTERS[27][12] ), .A2(n164), .B1(
        \REGISTERS[26][12] ), .B2(n161), .ZN(n909) );
  OAI221_X1 U1471 ( .B1(n122), .B2(n1918), .C1(n119), .C2(n1886), .A(n917), 
        .ZN(n912) );
  AOI22_X1 U1472 ( .A1(\REGISTERS[11][12] ), .A2(n116), .B1(
        \REGISTERS[10][12] ), .B2(n113), .ZN(n917) );
  OAI221_X1 U1473 ( .B1(n170), .B2(n2173), .C1(n167), .C2(n2141), .A(n891), 
        .ZN(n886) );
  AOI22_X1 U1474 ( .A1(\REGISTERS[27][13] ), .A2(n164), .B1(
        \REGISTERS[26][13] ), .B2(n161), .ZN(n891) );
  OAI221_X1 U1475 ( .B1(n122), .B2(n1917), .C1(n119), .C2(n1885), .A(n899), 
        .ZN(n894) );
  AOI22_X1 U1476 ( .A1(\REGISTERS[11][13] ), .A2(n116), .B1(
        \REGISTERS[10][13] ), .B2(n113), .ZN(n899) );
  OAI221_X1 U1477 ( .B1(n170), .B2(n2172), .C1(n167), .C2(n2140), .A(n873), 
        .ZN(n868) );
  AOI22_X1 U1478 ( .A1(\REGISTERS[27][14] ), .A2(n164), .B1(
        \REGISTERS[26][14] ), .B2(n161), .ZN(n873) );
  OAI221_X1 U1479 ( .B1(n122), .B2(n1916), .C1(n119), .C2(n1884), .A(n881), 
        .ZN(n876) );
  AOI22_X1 U1480 ( .A1(\REGISTERS[11][14] ), .A2(n116), .B1(
        \REGISTERS[10][14] ), .B2(n113), .ZN(n881) );
  OAI221_X1 U1481 ( .B1(n170), .B2(n2171), .C1(n167), .C2(n2139), .A(n855), 
        .ZN(n850) );
  AOI22_X1 U1482 ( .A1(\REGISTERS[27][15] ), .A2(n164), .B1(
        \REGISTERS[26][15] ), .B2(n161), .ZN(n855) );
  OAI221_X1 U1483 ( .B1(n122), .B2(n1915), .C1(n119), .C2(n1883), .A(n863), 
        .ZN(n858) );
  AOI22_X1 U1484 ( .A1(\REGISTERS[11][15] ), .A2(n116), .B1(
        \REGISTERS[10][15] ), .B2(n113), .ZN(n863) );
  OAI221_X1 U1485 ( .B1(n170), .B2(n2170), .C1(n167), .C2(n2138), .A(n837), 
        .ZN(n832) );
  AOI22_X1 U1486 ( .A1(\REGISTERS[27][16] ), .A2(n164), .B1(
        \REGISTERS[26][16] ), .B2(n161), .ZN(n837) );
  OAI221_X1 U1487 ( .B1(n122), .B2(n1914), .C1(n119), .C2(n1882), .A(n845), 
        .ZN(n840) );
  AOI22_X1 U1488 ( .A1(\REGISTERS[11][16] ), .A2(n116), .B1(
        \REGISTERS[10][16] ), .B2(n113), .ZN(n845) );
  OAI221_X1 U1489 ( .B1(n170), .B2(n2169), .C1(n167), .C2(n2137), .A(n819), 
        .ZN(n814) );
  AOI22_X1 U1490 ( .A1(\REGISTERS[27][17] ), .A2(n164), .B1(
        \REGISTERS[26][17] ), .B2(n161), .ZN(n819) );
  OAI221_X1 U1491 ( .B1(n122), .B2(n1913), .C1(n119), .C2(n1881), .A(n827), 
        .ZN(n822) );
  AOI22_X1 U1492 ( .A1(\REGISTERS[11][17] ), .A2(n116), .B1(
        \REGISTERS[10][17] ), .B2(n113), .ZN(n827) );
  OAI221_X1 U1493 ( .B1(n170), .B2(n2168), .C1(n167), .C2(n2136), .A(n801), 
        .ZN(n796) );
  AOI22_X1 U1494 ( .A1(\REGISTERS[27][18] ), .A2(n164), .B1(
        \REGISTERS[26][18] ), .B2(n161), .ZN(n801) );
  OAI221_X1 U1495 ( .B1(n122), .B2(n1912), .C1(n119), .C2(n1880), .A(n809), 
        .ZN(n804) );
  AOI22_X1 U1496 ( .A1(\REGISTERS[11][18] ), .A2(n116), .B1(
        \REGISTERS[10][18] ), .B2(n113), .ZN(n809) );
  OAI221_X1 U1497 ( .B1(n170), .B2(n2167), .C1(n167), .C2(n2135), .A(n783), 
        .ZN(n778) );
  AOI22_X1 U1498 ( .A1(\REGISTERS[27][19] ), .A2(n164), .B1(
        \REGISTERS[26][19] ), .B2(n161), .ZN(n783) );
  OAI221_X1 U1499 ( .B1(n122), .B2(n1911), .C1(n119), .C2(n1879), .A(n791), 
        .ZN(n786) );
  AOI22_X1 U1500 ( .A1(\REGISTERS[11][19] ), .A2(n116), .B1(
        \REGISTERS[10][19] ), .B2(n113), .ZN(n791) );
  OAI221_X1 U1501 ( .B1(n170), .B2(n2166), .C1(n167), .C2(n2134), .A(n765), 
        .ZN(n760) );
  AOI22_X1 U1502 ( .A1(\REGISTERS[27][20] ), .A2(n164), .B1(
        \REGISTERS[26][20] ), .B2(n161), .ZN(n765) );
  OAI221_X1 U1503 ( .B1(n122), .B2(n1910), .C1(n119), .C2(n1878), .A(n773), 
        .ZN(n768) );
  AOI22_X1 U1504 ( .A1(\REGISTERS[11][20] ), .A2(n116), .B1(
        \REGISTERS[10][20] ), .B2(n113), .ZN(n773) );
  OAI221_X1 U1505 ( .B1(n170), .B2(n2165), .C1(n167), .C2(n2133), .A(n747), 
        .ZN(n742) );
  AOI22_X1 U1506 ( .A1(\REGISTERS[27][21] ), .A2(n164), .B1(
        \REGISTERS[26][21] ), .B2(n161), .ZN(n747) );
  OAI221_X1 U1507 ( .B1(n122), .B2(n1909), .C1(n119), .C2(n1877), .A(n755), 
        .ZN(n750) );
  AOI22_X1 U1508 ( .A1(\REGISTERS[11][21] ), .A2(n116), .B1(
        \REGISTERS[10][21] ), .B2(n113), .ZN(n755) );
  OAI221_X1 U1509 ( .B1(n170), .B2(n2164), .C1(n168), .C2(n2132), .A(n729), 
        .ZN(n724) );
  AOI22_X1 U1510 ( .A1(\REGISTERS[27][22] ), .A2(n164), .B1(
        \REGISTERS[26][22] ), .B2(n161), .ZN(n729) );
  OAI221_X1 U1511 ( .B1(n122), .B2(n1908), .C1(n120), .C2(n1876), .A(n737), 
        .ZN(n732) );
  AOI22_X1 U1512 ( .A1(\REGISTERS[11][22] ), .A2(n116), .B1(
        \REGISTERS[10][22] ), .B2(n113), .ZN(n737) );
  OAI221_X1 U1513 ( .B1(n170), .B2(n2163), .C1(n168), .C2(n2131), .A(n711), 
        .ZN(n706) );
  AOI22_X1 U1514 ( .A1(\REGISTERS[27][23] ), .A2(n164), .B1(
        \REGISTERS[26][23] ), .B2(n161), .ZN(n711) );
  OAI221_X1 U1515 ( .B1(n122), .B2(n1907), .C1(n120), .C2(n1875), .A(n719), 
        .ZN(n714) );
  AOI22_X1 U1516 ( .A1(\REGISTERS[11][23] ), .A2(n116), .B1(
        \REGISTERS[10][23] ), .B2(n113), .ZN(n719) );
  OAI221_X1 U1517 ( .B1(n2175), .B2(n74), .C1(n2143), .C2(n71), .A(n1552), 
        .ZN(n1547) );
  AOI22_X1 U1518 ( .A1(n68), .A2(\REGISTERS[27][11] ), .B1(n65), .B2(
        \REGISTERS[26][11] ), .ZN(n1552) );
  OAI221_X1 U1519 ( .B1(n1919), .B2(n26), .C1(n1887), .C2(n23), .A(n1560), 
        .ZN(n1555) );
  AOI22_X1 U1520 ( .A1(n20), .A2(\REGISTERS[11][11] ), .B1(n17), .B2(
        \REGISTERS[10][11] ), .ZN(n1560) );
  OAI221_X1 U1521 ( .B1(n2174), .B2(n74), .C1(n2142), .C2(n71), .A(n1534), 
        .ZN(n1529) );
  AOI22_X1 U1522 ( .A1(n68), .A2(\REGISTERS[27][12] ), .B1(n65), .B2(
        \REGISTERS[26][12] ), .ZN(n1534) );
  OAI221_X1 U1523 ( .B1(n1918), .B2(n26), .C1(n1886), .C2(n23), .A(n1542), 
        .ZN(n1537) );
  AOI22_X1 U1524 ( .A1(n20), .A2(\REGISTERS[11][12] ), .B1(n17), .B2(
        \REGISTERS[10][12] ), .ZN(n1542) );
  OAI221_X1 U1525 ( .B1(n2173), .B2(n74), .C1(n2141), .C2(n71), .A(n1516), 
        .ZN(n1511) );
  AOI22_X1 U1526 ( .A1(n68), .A2(\REGISTERS[27][13] ), .B1(n65), .B2(
        \REGISTERS[26][13] ), .ZN(n1516) );
  OAI221_X1 U1527 ( .B1(n1917), .B2(n26), .C1(n1885), .C2(n23), .A(n1524), 
        .ZN(n1519) );
  AOI22_X1 U1528 ( .A1(n20), .A2(\REGISTERS[11][13] ), .B1(n17), .B2(
        \REGISTERS[10][13] ), .ZN(n1524) );
  OAI221_X1 U1529 ( .B1(n2172), .B2(n74), .C1(n2140), .C2(n71), .A(n1498), 
        .ZN(n1493) );
  AOI22_X1 U1530 ( .A1(n68), .A2(\REGISTERS[27][14] ), .B1(n65), .B2(
        \REGISTERS[26][14] ), .ZN(n1498) );
  OAI221_X1 U1531 ( .B1(n1916), .B2(n26), .C1(n1884), .C2(n23), .A(n1506), 
        .ZN(n1501) );
  AOI22_X1 U1532 ( .A1(n20), .A2(\REGISTERS[11][14] ), .B1(n17), .B2(
        \REGISTERS[10][14] ), .ZN(n1506) );
  OAI221_X1 U1533 ( .B1(n2171), .B2(n74), .C1(n2139), .C2(n71), .A(n1480), 
        .ZN(n1475) );
  AOI22_X1 U1534 ( .A1(n68), .A2(\REGISTERS[27][15] ), .B1(n65), .B2(
        \REGISTERS[26][15] ), .ZN(n1480) );
  OAI221_X1 U1535 ( .B1(n1915), .B2(n26), .C1(n1883), .C2(n23), .A(n1488), 
        .ZN(n1483) );
  AOI22_X1 U1536 ( .A1(n20), .A2(\REGISTERS[11][15] ), .B1(n17), .B2(
        \REGISTERS[10][15] ), .ZN(n1488) );
  OAI221_X1 U1537 ( .B1(n2170), .B2(n74), .C1(n2138), .C2(n71), .A(n1462), 
        .ZN(n1457) );
  AOI22_X1 U1538 ( .A1(n68), .A2(\REGISTERS[27][16] ), .B1(n65), .B2(
        \REGISTERS[26][16] ), .ZN(n1462) );
  OAI221_X1 U1539 ( .B1(n1914), .B2(n26), .C1(n1882), .C2(n23), .A(n1470), 
        .ZN(n1465) );
  AOI22_X1 U1540 ( .A1(n20), .A2(\REGISTERS[11][16] ), .B1(n17), .B2(
        \REGISTERS[10][16] ), .ZN(n1470) );
  OAI221_X1 U1541 ( .B1(n2169), .B2(n74), .C1(n2137), .C2(n71), .A(n1444), 
        .ZN(n1439) );
  AOI22_X1 U1542 ( .A1(n68), .A2(\REGISTERS[27][17] ), .B1(n65), .B2(
        \REGISTERS[26][17] ), .ZN(n1444) );
  OAI221_X1 U1543 ( .B1(n1913), .B2(n26), .C1(n1881), .C2(n23), .A(n1452), 
        .ZN(n1447) );
  AOI22_X1 U1544 ( .A1(n20), .A2(\REGISTERS[11][17] ), .B1(n17), .B2(
        \REGISTERS[10][17] ), .ZN(n1452) );
  OAI221_X1 U1545 ( .B1(n2168), .B2(n74), .C1(n2136), .C2(n71), .A(n1426), 
        .ZN(n1421) );
  AOI22_X1 U1546 ( .A1(n68), .A2(\REGISTERS[27][18] ), .B1(n65), .B2(
        \REGISTERS[26][18] ), .ZN(n1426) );
  OAI221_X1 U1547 ( .B1(n1912), .B2(n26), .C1(n1880), .C2(n23), .A(n1434), 
        .ZN(n1429) );
  AOI22_X1 U1548 ( .A1(n20), .A2(\REGISTERS[11][18] ), .B1(n17), .B2(
        \REGISTERS[10][18] ), .ZN(n1434) );
  OAI221_X1 U1549 ( .B1(n2167), .B2(n74), .C1(n2135), .C2(n71), .A(n1408), 
        .ZN(n1403) );
  AOI22_X1 U1550 ( .A1(n68), .A2(\REGISTERS[27][19] ), .B1(n65), .B2(
        \REGISTERS[26][19] ), .ZN(n1408) );
  OAI221_X1 U1551 ( .B1(n1911), .B2(n26), .C1(n1879), .C2(n23), .A(n1416), 
        .ZN(n1411) );
  AOI22_X1 U1552 ( .A1(n20), .A2(\REGISTERS[11][19] ), .B1(n17), .B2(
        \REGISTERS[10][19] ), .ZN(n1416) );
  OAI221_X1 U1553 ( .B1(n2166), .B2(n74), .C1(n2134), .C2(n71), .A(n1390), 
        .ZN(n1385) );
  AOI22_X1 U1554 ( .A1(n68), .A2(\REGISTERS[27][20] ), .B1(n65), .B2(
        \REGISTERS[26][20] ), .ZN(n1390) );
  OAI221_X1 U1555 ( .B1(n1910), .B2(n26), .C1(n1878), .C2(n23), .A(n1398), 
        .ZN(n1393) );
  AOI22_X1 U1556 ( .A1(n20), .A2(\REGISTERS[11][20] ), .B1(n17), .B2(
        \REGISTERS[10][20] ), .ZN(n1398) );
  OAI221_X1 U1557 ( .B1(n2165), .B2(n74), .C1(n2133), .C2(n71), .A(n1372), 
        .ZN(n1367) );
  AOI22_X1 U1558 ( .A1(n68), .A2(\REGISTERS[27][21] ), .B1(n65), .B2(
        \REGISTERS[26][21] ), .ZN(n1372) );
  OAI221_X1 U1559 ( .B1(n1909), .B2(n26), .C1(n1877), .C2(n23), .A(n1380), 
        .ZN(n1375) );
  AOI22_X1 U1560 ( .A1(n20), .A2(\REGISTERS[11][21] ), .B1(n17), .B2(
        \REGISTERS[10][21] ), .ZN(n1380) );
  OAI221_X1 U1561 ( .B1(n157), .B2(n2250), .C1(n154), .C2(n2218), .A(n1135), 
        .ZN(n1119) );
  AOI22_X1 U1562 ( .A1(\REGISTERS[29][0] ), .A2(n151), .B1(\REGISTERS[28][0] ), 
        .B2(n148), .ZN(n1135) );
  OAI221_X1 U1563 ( .B1(n157), .B2(n2249), .C1(n154), .C2(n2217), .A(n1108), 
        .ZN(n1101) );
  AOI22_X1 U1564 ( .A1(\REGISTERS[29][1] ), .A2(n151), .B1(\REGISTERS[28][1] ), 
        .B2(n148), .ZN(n1108) );
  OAI221_X1 U1565 ( .B1(n157), .B2(n2248), .C1(n154), .C2(n2216), .A(n1090), 
        .ZN(n1083) );
  AOI22_X1 U1566 ( .A1(\REGISTERS[29][2] ), .A2(n151), .B1(\REGISTERS[28][2] ), 
        .B2(n148), .ZN(n1090) );
  OAI221_X1 U1567 ( .B1(n157), .B2(n2247), .C1(n154), .C2(n2215), .A(n1072), 
        .ZN(n1065) );
  AOI22_X1 U1568 ( .A1(\REGISTERS[29][3] ), .A2(n151), .B1(\REGISTERS[28][3] ), 
        .B2(n148), .ZN(n1072) );
  OAI221_X1 U1569 ( .B1(n157), .B2(n2246), .C1(n154), .C2(n2214), .A(n1054), 
        .ZN(n1047) );
  AOI22_X1 U1570 ( .A1(\REGISTERS[29][4] ), .A2(n151), .B1(\REGISTERS[28][4] ), 
        .B2(n148), .ZN(n1054) );
  OAI221_X1 U1571 ( .B1(n157), .B2(n2245), .C1(n154), .C2(n2213), .A(n1036), 
        .ZN(n1029) );
  AOI22_X1 U1572 ( .A1(\REGISTERS[29][5] ), .A2(n151), .B1(\REGISTERS[28][5] ), 
        .B2(n148), .ZN(n1036) );
  OAI221_X1 U1573 ( .B1(n157), .B2(n2244), .C1(n154), .C2(n2212), .A(n1018), 
        .ZN(n1011) );
  AOI22_X1 U1574 ( .A1(\REGISTERS[29][6] ), .A2(n151), .B1(\REGISTERS[28][6] ), 
        .B2(n148), .ZN(n1018) );
  OAI221_X1 U1575 ( .B1(n157), .B2(n2243), .C1(n154), .C2(n2211), .A(n1000), 
        .ZN(n993) );
  AOI22_X1 U1576 ( .A1(\REGISTERS[29][7] ), .A2(n151), .B1(\REGISTERS[28][7] ), 
        .B2(n148), .ZN(n1000) );
  OAI221_X1 U1577 ( .B1(n157), .B2(n2242), .C1(n154), .C2(n2210), .A(n982), 
        .ZN(n975) );
  AOI22_X1 U1578 ( .A1(\REGISTERS[29][8] ), .A2(n151), .B1(\REGISTERS[28][8] ), 
        .B2(n148), .ZN(n982) );
  OAI221_X1 U1579 ( .B1(n157), .B2(n2241), .C1(n154), .C2(n2209), .A(n964), 
        .ZN(n957) );
  AOI22_X1 U1580 ( .A1(\REGISTERS[29][9] ), .A2(n151), .B1(\REGISTERS[28][9] ), 
        .B2(n148), .ZN(n964) );
  OAI221_X1 U1581 ( .B1(n157), .B2(n2240), .C1(n154), .C2(n2208), .A(n946), 
        .ZN(n939) );
  AOI22_X1 U1582 ( .A1(\REGISTERS[29][10] ), .A2(n151), .B1(
        \REGISTERS[28][10] ), .B2(n148), .ZN(n946) );
  OAI221_X1 U1583 ( .B1(n157), .B2(n2239), .C1(n155), .C2(n2207), .A(n928), 
        .ZN(n921) );
  AOI22_X1 U1584 ( .A1(\REGISTERS[29][11] ), .A2(n151), .B1(
        \REGISTERS[28][11] ), .B2(n148), .ZN(n928) );
  OAI221_X1 U1585 ( .B1(n158), .B2(n2238), .C1(n155), .C2(n2206), .A(n910), 
        .ZN(n903) );
  AOI22_X1 U1586 ( .A1(\REGISTERS[29][12] ), .A2(n152), .B1(
        \REGISTERS[28][12] ), .B2(n149), .ZN(n910) );
  OAI221_X1 U1587 ( .B1(n158), .B2(n2237), .C1(n155), .C2(n2205), .A(n892), 
        .ZN(n885) );
  AOI22_X1 U1588 ( .A1(\REGISTERS[29][13] ), .A2(n152), .B1(
        \REGISTERS[28][13] ), .B2(n149), .ZN(n892) );
  OAI221_X1 U1589 ( .B1(n158), .B2(n2236), .C1(n155), .C2(n2204), .A(n874), 
        .ZN(n867) );
  AOI22_X1 U1590 ( .A1(\REGISTERS[29][14] ), .A2(n152), .B1(
        \REGISTERS[28][14] ), .B2(n149), .ZN(n874) );
  OAI221_X1 U1591 ( .B1(n158), .B2(n2235), .C1(n155), .C2(n2203), .A(n856), 
        .ZN(n849) );
  AOI22_X1 U1592 ( .A1(\REGISTERS[29][15] ), .A2(n152), .B1(
        \REGISTERS[28][15] ), .B2(n149), .ZN(n856) );
  OAI221_X1 U1593 ( .B1(n158), .B2(n2234), .C1(n155), .C2(n2202), .A(n838), 
        .ZN(n831) );
  AOI22_X1 U1594 ( .A1(\REGISTERS[29][16] ), .A2(n152), .B1(
        \REGISTERS[28][16] ), .B2(n149), .ZN(n838) );
  OAI221_X1 U1595 ( .B1(n158), .B2(n2233), .C1(n155), .C2(n2201), .A(n820), 
        .ZN(n813) );
  AOI22_X1 U1596 ( .A1(\REGISTERS[29][17] ), .A2(n152), .B1(
        \REGISTERS[28][17] ), .B2(n149), .ZN(n820) );
  OAI221_X1 U1597 ( .B1(n158), .B2(n2232), .C1(n155), .C2(n2200), .A(n802), 
        .ZN(n795) );
  AOI22_X1 U1598 ( .A1(\REGISTERS[29][18] ), .A2(n152), .B1(
        \REGISTERS[28][18] ), .B2(n149), .ZN(n802) );
  OAI221_X1 U1599 ( .B1(n158), .B2(n2231), .C1(n155), .C2(n2199), .A(n784), 
        .ZN(n777) );
  AOI22_X1 U1600 ( .A1(\REGISTERS[29][19] ), .A2(n152), .B1(
        \REGISTERS[28][19] ), .B2(n149), .ZN(n784) );
  OAI221_X1 U1601 ( .B1(n158), .B2(n2230), .C1(n155), .C2(n2198), .A(n766), 
        .ZN(n759) );
  AOI22_X1 U1602 ( .A1(\REGISTERS[29][20] ), .A2(n152), .B1(
        \REGISTERS[28][20] ), .B2(n149), .ZN(n766) );
  OAI221_X1 U1603 ( .B1(n158), .B2(n2229), .C1(n155), .C2(n2197), .A(n748), 
        .ZN(n741) );
  AOI22_X1 U1604 ( .A1(\REGISTERS[29][21] ), .A2(n152), .B1(
        \REGISTERS[28][21] ), .B2(n149), .ZN(n748) );
  OAI221_X1 U1605 ( .B1(n158), .B2(n2228), .C1(n156), .C2(n2196), .A(n730), 
        .ZN(n723) );
  AOI22_X1 U1606 ( .A1(\REGISTERS[29][22] ), .A2(n152), .B1(
        \REGISTERS[28][22] ), .B2(n149), .ZN(n730) );
  OAI221_X1 U1607 ( .B1(n158), .B2(n2227), .C1(n156), .C2(n2195), .A(n712), 
        .ZN(n705) );
  AOI22_X1 U1608 ( .A1(\REGISTERS[29][23] ), .A2(n152), .B1(
        \REGISTERS[28][23] ), .B2(n149), .ZN(n712) );
  OAI221_X1 U1609 ( .B1(n2239), .B2(n62), .C1(n2207), .C2(n59), .A(n1553), 
        .ZN(n1546) );
  AOI22_X1 U1610 ( .A1(n56), .A2(\REGISTERS[29][11] ), .B1(n53), .B2(
        \REGISTERS[28][11] ), .ZN(n1553) );
  OAI221_X1 U1611 ( .B1(n2238), .B2(n62), .C1(n2206), .C2(n59), .A(n1535), 
        .ZN(n1528) );
  AOI22_X1 U1612 ( .A1(n56), .A2(\REGISTERS[29][12] ), .B1(n53), .B2(
        \REGISTERS[28][12] ), .ZN(n1535) );
  OAI221_X1 U1613 ( .B1(n2237), .B2(n62), .C1(n2205), .C2(n59), .A(n1517), 
        .ZN(n1510) );
  AOI22_X1 U1614 ( .A1(n56), .A2(\REGISTERS[29][13] ), .B1(n53), .B2(
        \REGISTERS[28][13] ), .ZN(n1517) );
  OAI221_X1 U1615 ( .B1(n2236), .B2(n62), .C1(n2204), .C2(n59), .A(n1499), 
        .ZN(n1492) );
  AOI22_X1 U1616 ( .A1(n56), .A2(\REGISTERS[29][14] ), .B1(n53), .B2(
        \REGISTERS[28][14] ), .ZN(n1499) );
  OAI221_X1 U1617 ( .B1(n2235), .B2(n62), .C1(n2203), .C2(n59), .A(n1481), 
        .ZN(n1474) );
  AOI22_X1 U1618 ( .A1(n56), .A2(\REGISTERS[29][15] ), .B1(n53), .B2(
        \REGISTERS[28][15] ), .ZN(n1481) );
  OAI221_X1 U1619 ( .B1(n2234), .B2(n62), .C1(n2202), .C2(n59), .A(n1463), 
        .ZN(n1456) );
  AOI22_X1 U1620 ( .A1(n56), .A2(\REGISTERS[29][16] ), .B1(n53), .B2(
        \REGISTERS[28][16] ), .ZN(n1463) );
  OAI221_X1 U1621 ( .B1(n2233), .B2(n62), .C1(n2201), .C2(n59), .A(n1445), 
        .ZN(n1438) );
  AOI22_X1 U1622 ( .A1(n56), .A2(\REGISTERS[29][17] ), .B1(n53), .B2(
        \REGISTERS[28][17] ), .ZN(n1445) );
  OAI221_X1 U1623 ( .B1(n2232), .B2(n62), .C1(n2200), .C2(n59), .A(n1427), 
        .ZN(n1420) );
  AOI22_X1 U1624 ( .A1(n56), .A2(\REGISTERS[29][18] ), .B1(n53), .B2(
        \REGISTERS[28][18] ), .ZN(n1427) );
  OAI221_X1 U1625 ( .B1(n2231), .B2(n62), .C1(n2199), .C2(n59), .A(n1409), 
        .ZN(n1402) );
  AOI22_X1 U1626 ( .A1(n56), .A2(\REGISTERS[29][19] ), .B1(n53), .B2(
        \REGISTERS[28][19] ), .ZN(n1409) );
  OAI221_X1 U1627 ( .B1(n2230), .B2(n62), .C1(n2198), .C2(n59), .A(n1391), 
        .ZN(n1384) );
  AOI22_X1 U1628 ( .A1(n56), .A2(\REGISTERS[29][20] ), .B1(n53), .B2(
        \REGISTERS[28][20] ), .ZN(n1391) );
  OAI221_X1 U1629 ( .B1(n2229), .B2(n62), .C1(n2197), .C2(n59), .A(n1373), 
        .ZN(n1366) );
  AOI22_X1 U1630 ( .A1(n56), .A2(\REGISTERS[29][21] ), .B1(n53), .B2(
        \REGISTERS[28][21] ), .ZN(n1373) );
  AOI22_X1 U1631 ( .A1(\REGISTERS[15][24] ), .A2(n105), .B1(
        \REGISTERS[14][24] ), .B2(n102), .ZN(n702) );
  AOI22_X1 U1632 ( .A1(\REGISTERS[15][25] ), .A2(n105), .B1(
        \REGISTERS[14][25] ), .B2(n102), .ZN(n684) );
  AOI22_X1 U1633 ( .A1(\REGISTERS[15][26] ), .A2(n105), .B1(
        \REGISTERS[14][26] ), .B2(n102), .ZN(n666) );
  AOI22_X1 U1634 ( .A1(\REGISTERS[15][27] ), .A2(n105), .B1(
        \REGISTERS[14][27] ), .B2(n102), .ZN(n648) );
  AOI22_X1 U1635 ( .A1(\REGISTERS[15][28] ), .A2(n105), .B1(
        \REGISTERS[14][28] ), .B2(n102), .ZN(n630) );
  AOI22_X1 U1636 ( .A1(\REGISTERS[15][29] ), .A2(n105), .B1(
        \REGISTERS[14][29] ), .B2(n102), .ZN(n612) );
  AOI22_X1 U1637 ( .A1(\REGISTERS[15][30] ), .A2(n105), .B1(
        \REGISTERS[14][30] ), .B2(n102), .ZN(n594) );
  AOI22_X1 U1638 ( .A1(\REGISTERS[15][31] ), .A2(n105), .B1(
        \REGISTERS[14][31] ), .B2(n102), .ZN(n574) );
  AOI22_X1 U1639 ( .A1(\REGISTERS[15][0] ), .A2(n103), .B1(\REGISTERS[14][0] ), 
        .B2(n100), .ZN(n1149) );
  AOI22_X1 U1640 ( .A1(\REGISTERS[15][1] ), .A2(n103), .B1(\REGISTERS[14][1] ), 
        .B2(n100), .ZN(n1116) );
  AOI22_X1 U1641 ( .A1(\REGISTERS[15][2] ), .A2(n103), .B1(\REGISTERS[14][2] ), 
        .B2(n100), .ZN(n1098) );
  AOI22_X1 U1642 ( .A1(\REGISTERS[15][3] ), .A2(n103), .B1(\REGISTERS[14][3] ), 
        .B2(n100), .ZN(n1080) );
  AOI22_X1 U1643 ( .A1(\REGISTERS[15][4] ), .A2(n103), .B1(\REGISTERS[14][4] ), 
        .B2(n100), .ZN(n1062) );
  AOI22_X1 U1644 ( .A1(\REGISTERS[15][5] ), .A2(n103), .B1(\REGISTERS[14][5] ), 
        .B2(n100), .ZN(n1044) );
  AOI22_X1 U1645 ( .A1(\REGISTERS[15][6] ), .A2(n103), .B1(\REGISTERS[14][6] ), 
        .B2(n100), .ZN(n1026) );
  AOI22_X1 U1646 ( .A1(\REGISTERS[15][7] ), .A2(n103), .B1(\REGISTERS[14][7] ), 
        .B2(n100), .ZN(n1008) );
  AOI22_X1 U1647 ( .A1(\REGISTERS[15][8] ), .A2(n103), .B1(\REGISTERS[14][8] ), 
        .B2(n100), .ZN(n990) );
  AOI22_X1 U1648 ( .A1(\REGISTERS[15][9] ), .A2(n103), .B1(\REGISTERS[14][9] ), 
        .B2(n100), .ZN(n972) );
  AOI22_X1 U1649 ( .A1(\REGISTERS[15][10] ), .A2(n103), .B1(
        \REGISTERS[14][10] ), .B2(n100), .ZN(n954) );
  AOI22_X1 U1650 ( .A1(\REGISTERS[15][11] ), .A2(n103), .B1(
        \REGISTERS[14][11] ), .B2(n100), .ZN(n936) );
  AOI22_X1 U1651 ( .A1(\REGISTERS[15][12] ), .A2(n104), .B1(
        \REGISTERS[14][12] ), .B2(n101), .ZN(n918) );
  AOI22_X1 U1652 ( .A1(\REGISTERS[15][13] ), .A2(n104), .B1(
        \REGISTERS[14][13] ), .B2(n101), .ZN(n900) );
  AOI22_X1 U1653 ( .A1(\REGISTERS[15][14] ), .A2(n104), .B1(
        \REGISTERS[14][14] ), .B2(n101), .ZN(n882) );
  AOI22_X1 U1654 ( .A1(\REGISTERS[15][15] ), .A2(n104), .B1(
        \REGISTERS[14][15] ), .B2(n101), .ZN(n864) );
  AOI22_X1 U1655 ( .A1(\REGISTERS[15][16] ), .A2(n104), .B1(
        \REGISTERS[14][16] ), .B2(n101), .ZN(n846) );
  AOI22_X1 U1656 ( .A1(\REGISTERS[15][17] ), .A2(n104), .B1(
        \REGISTERS[14][17] ), .B2(n101), .ZN(n828) );
  AOI22_X1 U1657 ( .A1(\REGISTERS[15][18] ), .A2(n104), .B1(
        \REGISTERS[14][18] ), .B2(n101), .ZN(n810) );
  AOI22_X1 U1658 ( .A1(\REGISTERS[15][19] ), .A2(n104), .B1(
        \REGISTERS[14][19] ), .B2(n101), .ZN(n792) );
  AOI22_X1 U1659 ( .A1(\REGISTERS[15][20] ), .A2(n104), .B1(
        \REGISTERS[14][20] ), .B2(n101), .ZN(n774) );
  AOI22_X1 U1660 ( .A1(\REGISTERS[15][21] ), .A2(n104), .B1(
        \REGISTERS[14][21] ), .B2(n101), .ZN(n756) );
  AOI22_X1 U1661 ( .A1(\REGISTERS[15][22] ), .A2(n104), .B1(
        \REGISTERS[14][22] ), .B2(n101), .ZN(n738) );
  AOI22_X1 U1662 ( .A1(\REGISTERS[15][23] ), .A2(n104), .B1(
        \REGISTERS[14][23] ), .B2(n101), .ZN(n720) );
  AOI22_X1 U1663 ( .A1(n7), .A2(\REGISTERS[15][0] ), .B1(n4), .B2(
        \REGISTERS[14][0] ), .ZN(n1774) );
  AOI22_X1 U1664 ( .A1(n7), .A2(\REGISTERS[15][1] ), .B1(n4), .B2(
        \REGISTERS[14][1] ), .ZN(n1741) );
  AOI22_X1 U1665 ( .A1(n7), .A2(\REGISTERS[15][2] ), .B1(n4), .B2(
        \REGISTERS[14][2] ), .ZN(n1723) );
  AOI22_X1 U1666 ( .A1(n7), .A2(\REGISTERS[15][3] ), .B1(n4), .B2(
        \REGISTERS[14][3] ), .ZN(n1705) );
  AOI22_X1 U1667 ( .A1(n7), .A2(\REGISTERS[15][4] ), .B1(n4), .B2(
        \REGISTERS[14][4] ), .ZN(n1687) );
  AOI22_X1 U1668 ( .A1(n7), .A2(\REGISTERS[15][5] ), .B1(n4), .B2(
        \REGISTERS[14][5] ), .ZN(n1669) );
  AOI22_X1 U1669 ( .A1(n7), .A2(\REGISTERS[15][6] ), .B1(n4), .B2(
        \REGISTERS[14][6] ), .ZN(n1651) );
  AOI22_X1 U1670 ( .A1(n7), .A2(\REGISTERS[15][7] ), .B1(n4), .B2(
        \REGISTERS[14][7] ), .ZN(n1633) );
  AOI22_X1 U1671 ( .A1(n7), .A2(\REGISTERS[15][8] ), .B1(n4), .B2(
        \REGISTERS[14][8] ), .ZN(n1615) );
  AOI22_X1 U1672 ( .A1(n7), .A2(\REGISTERS[15][9] ), .B1(n4), .B2(
        \REGISTERS[14][9] ), .ZN(n1597) );
  AOI22_X1 U1673 ( .A1(n7), .A2(\REGISTERS[15][10] ), .B1(n4), .B2(
        \REGISTERS[14][10] ), .ZN(n1579) );
  AOI22_X1 U1674 ( .A1(n8), .A2(\REGISTERS[15][11] ), .B1(n5), .B2(
        \REGISTERS[14][11] ), .ZN(n1561) );
  AOI22_X1 U1675 ( .A1(n8), .A2(\REGISTERS[15][12] ), .B1(n5), .B2(
        \REGISTERS[14][12] ), .ZN(n1543) );
  AOI22_X1 U1676 ( .A1(n8), .A2(\REGISTERS[15][13] ), .B1(n5), .B2(
        \REGISTERS[14][13] ), .ZN(n1525) );
  AOI22_X1 U1677 ( .A1(n8), .A2(\REGISTERS[15][14] ), .B1(n5), .B2(
        \REGISTERS[14][14] ), .ZN(n1507) );
  AOI22_X1 U1678 ( .A1(n8), .A2(\REGISTERS[15][15] ), .B1(n5), .B2(
        \REGISTERS[14][15] ), .ZN(n1489) );
  AOI22_X1 U1679 ( .A1(n8), .A2(\REGISTERS[15][16] ), .B1(n5), .B2(
        \REGISTERS[14][16] ), .ZN(n1471) );
  AOI22_X1 U1680 ( .A1(n8), .A2(\REGISTERS[15][17] ), .B1(n5), .B2(
        \REGISTERS[14][17] ), .ZN(n1453) );
  AOI22_X1 U1681 ( .A1(n8), .A2(\REGISTERS[15][18] ), .B1(n5), .B2(
        \REGISTERS[14][18] ), .ZN(n1435) );
  AOI22_X1 U1682 ( .A1(n8), .A2(\REGISTERS[15][19] ), .B1(n5), .B2(
        \REGISTERS[14][19] ), .ZN(n1417) );
  AOI22_X1 U1683 ( .A1(n8), .A2(\REGISTERS[15][20] ), .B1(n5), .B2(
        \REGISTERS[14][20] ), .ZN(n1399) );
  AOI22_X1 U1684 ( .A1(n8), .A2(\REGISTERS[15][21] ), .B1(n5), .B2(
        \REGISTERS[14][21] ), .ZN(n1381) );
  AOI22_X1 U1685 ( .A1(n9), .A2(\REGISTERS[15][22] ), .B1(n6), .B2(
        \REGISTERS[14][22] ), .ZN(n1363) );
  AOI22_X1 U1686 ( .A1(n9), .A2(\REGISTERS[15][23] ), .B1(n6), .B2(
        \REGISTERS[14][23] ), .ZN(n1345) );
  AOI22_X1 U1687 ( .A1(n9), .A2(\REGISTERS[15][24] ), .B1(n6), .B2(
        \REGISTERS[14][24] ), .ZN(n1327) );
  AOI22_X1 U1688 ( .A1(n9), .A2(\REGISTERS[15][25] ), .B1(n6), .B2(
        \REGISTERS[14][25] ), .ZN(n1309) );
  AOI22_X1 U1689 ( .A1(n9), .A2(\REGISTERS[15][26] ), .B1(n6), .B2(
        \REGISTERS[14][26] ), .ZN(n1291) );
  AOI22_X1 U1690 ( .A1(n9), .A2(\REGISTERS[15][27] ), .B1(n6), .B2(
        \REGISTERS[14][27] ), .ZN(n1273) );
  AOI22_X1 U1691 ( .A1(n9), .A2(\REGISTERS[15][28] ), .B1(n6), .B2(
        \REGISTERS[14][28] ), .ZN(n1255) );
  AOI22_X1 U1692 ( .A1(n9), .A2(\REGISTERS[15][29] ), .B1(n6), .B2(
        \REGISTERS[14][29] ), .ZN(n1237) );
  AOI22_X1 U1693 ( .A1(n9), .A2(\REGISTERS[15][30] ), .B1(n6), .B2(
        \REGISTERS[14][30] ), .ZN(n1219) );
  AOI22_X1 U1694 ( .A1(n9), .A2(\REGISTERS[15][31] ), .B1(n6), .B2(
        \REGISTERS[14][31] ), .ZN(n1199) );
  INV_X1 U1695 ( .A(ADD_WR[0]), .ZN(n2259) );
  INV_X1 U1696 ( .A(ADD_WR[1]), .ZN(n2260) );
  INV_X1 U1697 ( .A(ADD_WR[2]), .ZN(n2261) );
  INV_X1 U1698 ( .A(ADD_WR[3]), .ZN(n2262) );
  INV_X1 U1699 ( .A(ADD_WR[4]), .ZN(n2263) );
  OR3_X1 U1700 ( .A1(ADD_WR[3]), .A2(ADD_WR[4]), .A3(n1786), .ZN(n1777) );
  INV_X1 U1701 ( .A(\REGISTERS[17][0] ), .ZN(n2058) );
  INV_X1 U1702 ( .A(\REGISTERS[21][0] ), .ZN(n2122) );
  INV_X1 U1703 ( .A(\REGISTERS[25][0] ), .ZN(n2186) );
  INV_X1 U1704 ( .A(\REGISTERS[31][0] ), .ZN(n2250) );
  INV_X1 U1705 ( .A(\REGISTERS[1][0] ), .ZN(n1802) );
  INV_X1 U1706 ( .A(\REGISTERS[5][0] ), .ZN(n1866) );
  INV_X1 U1707 ( .A(\REGISTERS[9][0] ), .ZN(n1930) );
  INV_X1 U1708 ( .A(\REGISTERS[13][0] ), .ZN(n1994) );
  INV_X1 U1709 ( .A(\REGISTERS[17][1] ), .ZN(n2057) );
  INV_X1 U1710 ( .A(\REGISTERS[21][1] ), .ZN(n2121) );
  INV_X1 U1711 ( .A(\REGISTERS[25][1] ), .ZN(n2185) );
  INV_X1 U1712 ( .A(\REGISTERS[31][1] ), .ZN(n2249) );
  INV_X1 U1713 ( .A(\REGISTERS[1][1] ), .ZN(n1801) );
  INV_X1 U1714 ( .A(\REGISTERS[5][1] ), .ZN(n1865) );
  INV_X1 U1715 ( .A(\REGISTERS[9][1] ), .ZN(n1929) );
  INV_X1 U1716 ( .A(\REGISTERS[13][1] ), .ZN(n1993) );
  INV_X1 U1717 ( .A(\REGISTERS[17][2] ), .ZN(n2056) );
  INV_X1 U1718 ( .A(\REGISTERS[21][2] ), .ZN(n2120) );
  INV_X1 U1719 ( .A(\REGISTERS[25][2] ), .ZN(n2184) );
  INV_X1 U1720 ( .A(\REGISTERS[31][2] ), .ZN(n2248) );
  INV_X1 U1721 ( .A(\REGISTERS[1][2] ), .ZN(n1800) );
  INV_X1 U1722 ( .A(\REGISTERS[5][2] ), .ZN(n1864) );
  INV_X1 U1723 ( .A(\REGISTERS[9][2] ), .ZN(n1928) );
  INV_X1 U1724 ( .A(\REGISTERS[13][2] ), .ZN(n1992) );
  INV_X1 U1725 ( .A(\REGISTERS[17][3] ), .ZN(n2055) );
  INV_X1 U1726 ( .A(\REGISTERS[21][3] ), .ZN(n2119) );
  INV_X1 U1727 ( .A(\REGISTERS[25][3] ), .ZN(n2183) );
  INV_X1 U1728 ( .A(\REGISTERS[31][3] ), .ZN(n2247) );
  INV_X1 U1729 ( .A(\REGISTERS[1][3] ), .ZN(n1799) );
  INV_X1 U1730 ( .A(\REGISTERS[5][3] ), .ZN(n1863) );
  INV_X1 U1731 ( .A(\REGISTERS[9][3] ), .ZN(n1927) );
  INV_X1 U1732 ( .A(\REGISTERS[13][3] ), .ZN(n1991) );
  INV_X1 U1733 ( .A(\REGISTERS[17][4] ), .ZN(n2054) );
  INV_X1 U1734 ( .A(\REGISTERS[21][4] ), .ZN(n2118) );
  INV_X1 U1735 ( .A(\REGISTERS[25][4] ), .ZN(n2182) );
  INV_X1 U1736 ( .A(\REGISTERS[31][4] ), .ZN(n2246) );
  INV_X1 U1737 ( .A(\REGISTERS[1][4] ), .ZN(n1798) );
  INV_X1 U1738 ( .A(\REGISTERS[5][4] ), .ZN(n1862) );
  INV_X1 U1739 ( .A(\REGISTERS[9][4] ), .ZN(n1926) );
  INV_X1 U1740 ( .A(\REGISTERS[13][4] ), .ZN(n1990) );
  INV_X1 U1741 ( .A(\REGISTERS[17][5] ), .ZN(n2053) );
  INV_X1 U1742 ( .A(\REGISTERS[21][5] ), .ZN(n2117) );
  INV_X1 U1743 ( .A(\REGISTERS[25][5] ), .ZN(n2181) );
  INV_X1 U1744 ( .A(\REGISTERS[31][5] ), .ZN(n2245) );
  INV_X1 U1745 ( .A(\REGISTERS[1][5] ), .ZN(n1797) );
  INV_X1 U1746 ( .A(\REGISTERS[5][5] ), .ZN(n1861) );
  INV_X1 U1747 ( .A(\REGISTERS[9][5] ), .ZN(n1925) );
  INV_X1 U1748 ( .A(\REGISTERS[13][5] ), .ZN(n1989) );
  INV_X1 U1749 ( .A(\REGISTERS[17][6] ), .ZN(n2052) );
  INV_X1 U1750 ( .A(\REGISTERS[21][6] ), .ZN(n2116) );
  INV_X1 U1751 ( .A(\REGISTERS[25][6] ), .ZN(n2180) );
  INV_X1 U1752 ( .A(\REGISTERS[31][6] ), .ZN(n2244) );
  INV_X1 U1753 ( .A(\REGISTERS[1][6] ), .ZN(n1796) );
  INV_X1 U1754 ( .A(\REGISTERS[5][6] ), .ZN(n1860) );
  INV_X1 U1755 ( .A(\REGISTERS[9][6] ), .ZN(n1924) );
  INV_X1 U1756 ( .A(\REGISTERS[13][6] ), .ZN(n1988) );
  INV_X1 U1757 ( .A(\REGISTERS[17][7] ), .ZN(n2051) );
  INV_X1 U1758 ( .A(\REGISTERS[21][7] ), .ZN(n2115) );
  INV_X1 U1759 ( .A(\REGISTERS[25][7] ), .ZN(n2179) );
  INV_X1 U1760 ( .A(\REGISTERS[31][7] ), .ZN(n2243) );
  INV_X1 U1761 ( .A(\REGISTERS[1][7] ), .ZN(n1795) );
  INV_X1 U1762 ( .A(\REGISTERS[5][7] ), .ZN(n1859) );
  INV_X1 U1763 ( .A(\REGISTERS[9][7] ), .ZN(n1923) );
  INV_X1 U1764 ( .A(\REGISTERS[13][7] ), .ZN(n1987) );
  INV_X1 U1765 ( .A(\REGISTERS[17][8] ), .ZN(n2050) );
  INV_X1 U1766 ( .A(\REGISTERS[21][8] ), .ZN(n2114) );
  INV_X1 U1767 ( .A(\REGISTERS[25][8] ), .ZN(n2178) );
  INV_X1 U1768 ( .A(\REGISTERS[31][8] ), .ZN(n2242) );
  INV_X1 U1769 ( .A(\REGISTERS[1][8] ), .ZN(n1794) );
  INV_X1 U1770 ( .A(\REGISTERS[5][8] ), .ZN(n1858) );
  INV_X1 U1771 ( .A(\REGISTERS[9][8] ), .ZN(n1922) );
  INV_X1 U1772 ( .A(\REGISTERS[13][8] ), .ZN(n1986) );
  INV_X1 U1773 ( .A(\REGISTERS[17][9] ), .ZN(n2049) );
  INV_X1 U1774 ( .A(\REGISTERS[21][9] ), .ZN(n2113) );
  INV_X1 U1775 ( .A(\REGISTERS[25][9] ), .ZN(n2177) );
  INV_X1 U1776 ( .A(\REGISTERS[31][9] ), .ZN(n2241) );
  INV_X1 U1777 ( .A(\REGISTERS[1][9] ), .ZN(n1793) );
  INV_X1 U1778 ( .A(\REGISTERS[5][9] ), .ZN(n1857) );
  INV_X1 U1779 ( .A(\REGISTERS[9][9] ), .ZN(n1921) );
  INV_X1 U1780 ( .A(\REGISTERS[13][9] ), .ZN(n1985) );
  INV_X1 U1781 ( .A(\REGISTERS[17][10] ), .ZN(n2048) );
  INV_X1 U1782 ( .A(\REGISTERS[21][10] ), .ZN(n2112) );
  INV_X1 U1783 ( .A(\REGISTERS[25][10] ), .ZN(n2176) );
  INV_X1 U1784 ( .A(\REGISTERS[31][10] ), .ZN(n2240) );
  INV_X1 U1785 ( .A(\REGISTERS[1][10] ), .ZN(n1792) );
  INV_X1 U1786 ( .A(\REGISTERS[5][10] ), .ZN(n1856) );
  INV_X1 U1787 ( .A(\REGISTERS[9][10] ), .ZN(n1920) );
  INV_X1 U1788 ( .A(\REGISTERS[13][10] ), .ZN(n1984) );
  INV_X1 U1789 ( .A(\REGISTERS[17][11] ), .ZN(n2047) );
  INV_X1 U1790 ( .A(\REGISTERS[21][11] ), .ZN(n2111) );
  INV_X1 U1791 ( .A(\REGISTERS[25][11] ), .ZN(n2175) );
  INV_X1 U1792 ( .A(\REGISTERS[31][11] ), .ZN(n2239) );
  INV_X1 U1793 ( .A(\REGISTERS[1][11] ), .ZN(n1791) );
  INV_X1 U1794 ( .A(\REGISTERS[5][11] ), .ZN(n1855) );
  INV_X1 U1795 ( .A(\REGISTERS[9][11] ), .ZN(n1919) );
  INV_X1 U1796 ( .A(\REGISTERS[13][11] ), .ZN(n1983) );
  INV_X1 U1797 ( .A(\REGISTERS[17][12] ), .ZN(n2046) );
  INV_X1 U1798 ( .A(\REGISTERS[21][12] ), .ZN(n2110) );
  INV_X1 U1799 ( .A(\REGISTERS[25][12] ), .ZN(n2174) );
  INV_X1 U1800 ( .A(\REGISTERS[31][12] ), .ZN(n2238) );
  INV_X1 U1801 ( .A(\REGISTERS[1][12] ), .ZN(n526) );
  INV_X1 U1802 ( .A(\REGISTERS[5][12] ), .ZN(n1854) );
  INV_X1 U1803 ( .A(\REGISTERS[9][12] ), .ZN(n1918) );
  INV_X1 U1804 ( .A(\REGISTERS[13][12] ), .ZN(n1982) );
  INV_X1 U1805 ( .A(\REGISTERS[17][13] ), .ZN(n2045) );
  INV_X1 U1806 ( .A(\REGISTERS[21][13] ), .ZN(n2109) );
  INV_X1 U1807 ( .A(\REGISTERS[25][13] ), .ZN(n2173) );
  INV_X1 U1808 ( .A(\REGISTERS[31][13] ), .ZN(n2237) );
  INV_X1 U1809 ( .A(\REGISTERS[1][13] ), .ZN(n525) );
  INV_X1 U1810 ( .A(\REGISTERS[5][13] ), .ZN(n1853) );
  INV_X1 U1811 ( .A(\REGISTERS[9][13] ), .ZN(n1917) );
  INV_X1 U1812 ( .A(\REGISTERS[13][13] ), .ZN(n1981) );
  INV_X1 U1813 ( .A(\REGISTERS[17][14] ), .ZN(n2044) );
  INV_X1 U1814 ( .A(\REGISTERS[21][14] ), .ZN(n2108) );
  INV_X1 U1815 ( .A(\REGISTERS[25][14] ), .ZN(n2172) );
  INV_X1 U1816 ( .A(\REGISTERS[31][14] ), .ZN(n2236) );
  INV_X1 U1817 ( .A(\REGISTERS[1][14] ), .ZN(n524) );
  INV_X1 U1818 ( .A(\REGISTERS[5][14] ), .ZN(n1852) );
  INV_X1 U1819 ( .A(\REGISTERS[9][14] ), .ZN(n1916) );
  INV_X1 U1820 ( .A(\REGISTERS[13][14] ), .ZN(n1980) );
  INV_X1 U1821 ( .A(\REGISTERS[17][15] ), .ZN(n2043) );
  INV_X1 U1822 ( .A(\REGISTERS[21][15] ), .ZN(n2107) );
  INV_X1 U1823 ( .A(\REGISTERS[25][15] ), .ZN(n2171) );
  INV_X1 U1824 ( .A(\REGISTERS[31][15] ), .ZN(n2235) );
  INV_X1 U1825 ( .A(\REGISTERS[1][15] ), .ZN(n523) );
  INV_X1 U1826 ( .A(\REGISTERS[5][15] ), .ZN(n1851) );
  INV_X1 U1827 ( .A(\REGISTERS[9][15] ), .ZN(n1915) );
  INV_X1 U1828 ( .A(\REGISTERS[13][15] ), .ZN(n1979) );
  INV_X1 U1829 ( .A(\REGISTERS[17][16] ), .ZN(n2042) );
  INV_X1 U1830 ( .A(\REGISTERS[21][16] ), .ZN(n2106) );
  INV_X1 U1831 ( .A(\REGISTERS[25][16] ), .ZN(n2170) );
  INV_X1 U1832 ( .A(\REGISTERS[31][16] ), .ZN(n2234) );
  INV_X1 U1833 ( .A(\REGISTERS[1][16] ), .ZN(n522) );
  INV_X1 U1834 ( .A(\REGISTERS[5][16] ), .ZN(n1850) );
  INV_X1 U1835 ( .A(\REGISTERS[9][16] ), .ZN(n1914) );
  INV_X1 U1836 ( .A(\REGISTERS[13][16] ), .ZN(n1978) );
  INV_X1 U1837 ( .A(\REGISTERS[17][17] ), .ZN(n2041) );
  INV_X1 U1838 ( .A(\REGISTERS[21][17] ), .ZN(n2105) );
  INV_X1 U1839 ( .A(\REGISTERS[25][17] ), .ZN(n2169) );
  INV_X1 U1840 ( .A(\REGISTERS[31][17] ), .ZN(n2233) );
  INV_X1 U1841 ( .A(\REGISTERS[1][17] ), .ZN(n521) );
  INV_X1 U1842 ( .A(\REGISTERS[5][17] ), .ZN(n1849) );
  INV_X1 U1843 ( .A(\REGISTERS[9][17] ), .ZN(n1913) );
  INV_X1 U1844 ( .A(\REGISTERS[13][17] ), .ZN(n1977) );
  INV_X1 U1845 ( .A(\REGISTERS[17][18] ), .ZN(n2040) );
  INV_X1 U1846 ( .A(\REGISTERS[21][18] ), .ZN(n2104) );
  INV_X1 U1847 ( .A(\REGISTERS[25][18] ), .ZN(n2168) );
  INV_X1 U1848 ( .A(\REGISTERS[31][18] ), .ZN(n2232) );
  INV_X1 U1849 ( .A(\REGISTERS[1][18] ), .ZN(n520) );
  INV_X1 U1850 ( .A(\REGISTERS[5][18] ), .ZN(n1848) );
  INV_X1 U1851 ( .A(\REGISTERS[9][18] ), .ZN(n1912) );
  INV_X1 U1852 ( .A(\REGISTERS[13][18] ), .ZN(n1976) );
  INV_X1 U1853 ( .A(\REGISTERS[17][19] ), .ZN(n2039) );
  INV_X1 U1854 ( .A(\REGISTERS[21][19] ), .ZN(n2103) );
  INV_X1 U1855 ( .A(\REGISTERS[25][19] ), .ZN(n2167) );
  INV_X1 U1856 ( .A(\REGISTERS[31][19] ), .ZN(n2231) );
  INV_X1 U1857 ( .A(\REGISTERS[1][19] ), .ZN(n519) );
  INV_X1 U1858 ( .A(\REGISTERS[5][19] ), .ZN(n1847) );
  INV_X1 U1859 ( .A(\REGISTERS[9][19] ), .ZN(n1911) );
  INV_X1 U1860 ( .A(\REGISTERS[13][19] ), .ZN(n1975) );
  INV_X1 U1861 ( .A(\REGISTERS[17][20] ), .ZN(n2038) );
  INV_X1 U1862 ( .A(\REGISTERS[21][20] ), .ZN(n2102) );
  INV_X1 U1863 ( .A(\REGISTERS[25][20] ), .ZN(n2166) );
  INV_X1 U1864 ( .A(\REGISTERS[31][20] ), .ZN(n2230) );
  INV_X1 U1865 ( .A(\REGISTERS[1][20] ), .ZN(n518) );
  INV_X1 U1866 ( .A(\REGISTERS[5][20] ), .ZN(n1846) );
  INV_X1 U1867 ( .A(\REGISTERS[9][20] ), .ZN(n1910) );
  INV_X1 U1868 ( .A(\REGISTERS[13][20] ), .ZN(n1974) );
  INV_X1 U1869 ( .A(\REGISTERS[17][21] ), .ZN(n2037) );
  INV_X1 U1870 ( .A(\REGISTERS[21][21] ), .ZN(n2101) );
  INV_X1 U1871 ( .A(\REGISTERS[25][21] ), .ZN(n2165) );
  INV_X1 U1872 ( .A(\REGISTERS[31][21] ), .ZN(n2229) );
  INV_X1 U1873 ( .A(\REGISTERS[1][21] ), .ZN(n517) );
  INV_X1 U1874 ( .A(\REGISTERS[5][21] ), .ZN(n1845) );
  INV_X1 U1875 ( .A(\REGISTERS[9][21] ), .ZN(n1909) );
  INV_X1 U1876 ( .A(\REGISTERS[13][21] ), .ZN(n1973) );
  INV_X1 U1877 ( .A(\REGISTERS[17][22] ), .ZN(n2036) );
  INV_X1 U1878 ( .A(\REGISTERS[21][22] ), .ZN(n2100) );
  INV_X1 U1879 ( .A(\REGISTERS[25][22] ), .ZN(n2164) );
  INV_X1 U1880 ( .A(\REGISTERS[31][22] ), .ZN(n2228) );
  INV_X1 U1881 ( .A(\REGISTERS[1][22] ), .ZN(n516) );
  INV_X1 U1882 ( .A(\REGISTERS[5][22] ), .ZN(n1844) );
  INV_X1 U1883 ( .A(\REGISTERS[9][22] ), .ZN(n1908) );
  INV_X1 U1884 ( .A(\REGISTERS[13][22] ), .ZN(n1972) );
  INV_X1 U1885 ( .A(\REGISTERS[17][23] ), .ZN(n2035) );
  INV_X1 U1886 ( .A(\REGISTERS[21][23] ), .ZN(n2099) );
  INV_X1 U1887 ( .A(\REGISTERS[25][23] ), .ZN(n2163) );
  INV_X1 U1888 ( .A(\REGISTERS[31][23] ), .ZN(n2227) );
  INV_X1 U1889 ( .A(\REGISTERS[1][23] ), .ZN(n515) );
  INV_X1 U1890 ( .A(\REGISTERS[5][23] ), .ZN(n1843) );
  INV_X1 U1891 ( .A(\REGISTERS[9][23] ), .ZN(n1907) );
  INV_X1 U1892 ( .A(\REGISTERS[13][23] ), .ZN(n1971) );
  INV_X1 U1893 ( .A(\REGISTERS[17][24] ), .ZN(n2034) );
  INV_X1 U1894 ( .A(\REGISTERS[21][24] ), .ZN(n2098) );
  INV_X1 U1895 ( .A(\REGISTERS[25][24] ), .ZN(n2162) );
  INV_X1 U1896 ( .A(\REGISTERS[31][24] ), .ZN(n2226) );
  INV_X1 U1897 ( .A(\REGISTERS[1][24] ), .ZN(n514) );
  INV_X1 U1898 ( .A(\REGISTERS[5][24] ), .ZN(n1842) );
  INV_X1 U1899 ( .A(\REGISTERS[9][24] ), .ZN(n1906) );
  INV_X1 U1900 ( .A(\REGISTERS[13][24] ), .ZN(n1970) );
  INV_X1 U1901 ( .A(\REGISTERS[17][25] ), .ZN(n2033) );
  INV_X1 U1902 ( .A(\REGISTERS[21][25] ), .ZN(n2097) );
  INV_X1 U1903 ( .A(\REGISTERS[25][25] ), .ZN(n2161) );
  INV_X1 U1904 ( .A(\REGISTERS[31][25] ), .ZN(n2225) );
  INV_X1 U1905 ( .A(\REGISTERS[1][25] ), .ZN(n513) );
  INV_X1 U1906 ( .A(\REGISTERS[5][25] ), .ZN(n1841) );
  INV_X1 U1907 ( .A(\REGISTERS[9][25] ), .ZN(n1905) );
  INV_X1 U1908 ( .A(\REGISTERS[13][25] ), .ZN(n1969) );
  INV_X1 U1909 ( .A(\REGISTERS[17][26] ), .ZN(n2032) );
  INV_X1 U1910 ( .A(\REGISTERS[21][26] ), .ZN(n2096) );
  INV_X1 U1923 ( .A(\REGISTERS[25][26] ), .ZN(n2160) );
  INV_X1 U1924 ( .A(\REGISTERS[31][26] ), .ZN(n2224) );
  INV_X1 U1925 ( .A(\REGISTERS[1][26] ), .ZN(n512) );
  INV_X1 U1926 ( .A(\REGISTERS[5][26] ), .ZN(n1840) );
  INV_X1 U1927 ( .A(\REGISTERS[9][26] ), .ZN(n1904) );
  INV_X1 U1928 ( .A(\REGISTERS[13][26] ), .ZN(n1968) );
  INV_X1 U1929 ( .A(\REGISTERS[17][27] ), .ZN(n2031) );
  INV_X1 U1930 ( .A(\REGISTERS[21][27] ), .ZN(n2095) );
  INV_X1 U1931 ( .A(\REGISTERS[25][27] ), .ZN(n2159) );
  INV_X1 U1932 ( .A(\REGISTERS[31][27] ), .ZN(n2223) );
  INV_X1 U1933 ( .A(\REGISTERS[1][27] ), .ZN(n511) );
  INV_X1 U1934 ( .A(\REGISTERS[5][27] ), .ZN(n1839) );
  INV_X1 U1935 ( .A(\REGISTERS[9][27] ), .ZN(n1903) );
  INV_X1 U1936 ( .A(\REGISTERS[13][27] ), .ZN(n1967) );
  INV_X1 U1937 ( .A(\REGISTERS[17][28] ), .ZN(n2030) );
  INV_X1 U1938 ( .A(\REGISTERS[21][28] ), .ZN(n2094) );
  INV_X1 U1939 ( .A(\REGISTERS[25][28] ), .ZN(n2158) );
  INV_X1 U1940 ( .A(\REGISTERS[31][28] ), .ZN(n2222) );
  INV_X1 U1941 ( .A(\REGISTERS[1][28] ), .ZN(n510) );
  INV_X1 U1942 ( .A(\REGISTERS[5][28] ), .ZN(n1838) );
  INV_X1 U1943 ( .A(\REGISTERS[9][28] ), .ZN(n1902) );
  INV_X1 U1944 ( .A(\REGISTERS[13][28] ), .ZN(n1966) );
  INV_X1 U1945 ( .A(\REGISTERS[17][29] ), .ZN(n2029) );
  INV_X1 U1946 ( .A(\REGISTERS[21][29] ), .ZN(n2093) );
  INV_X1 U1947 ( .A(\REGISTERS[25][29] ), .ZN(n2157) );
  INV_X1 U1948 ( .A(\REGISTERS[31][29] ), .ZN(n2221) );
  INV_X1 U1949 ( .A(\REGISTERS[1][29] ), .ZN(n509) );
  INV_X1 U1950 ( .A(\REGISTERS[5][29] ), .ZN(n1837) );
  INV_X1 U1951 ( .A(\REGISTERS[9][29] ), .ZN(n1901) );
  INV_X1 U1952 ( .A(\REGISTERS[13][29] ), .ZN(n1965) );
  INV_X1 U1953 ( .A(\REGISTERS[17][30] ), .ZN(n2028) );
  INV_X1 U1954 ( .A(\REGISTERS[21][30] ), .ZN(n2092) );
  INV_X1 U1955 ( .A(\REGISTERS[25][30] ), .ZN(n2156) );
  INV_X1 U1956 ( .A(\REGISTERS[31][30] ), .ZN(n2220) );
  INV_X1 U1957 ( .A(\REGISTERS[1][30] ), .ZN(n508) );
  INV_X1 U1958 ( .A(\REGISTERS[5][30] ), .ZN(n1836) );
  INV_X1 U1959 ( .A(\REGISTERS[9][30] ), .ZN(n1900) );
  INV_X1 U1960 ( .A(\REGISTERS[13][30] ), .ZN(n1964) );
  INV_X1 U1961 ( .A(\REGISTERS[17][31] ), .ZN(n2027) );
  INV_X1 U1962 ( .A(\REGISTERS[21][31] ), .ZN(n2091) );
  INV_X1 U1963 ( .A(\REGISTERS[25][31] ), .ZN(n2155) );
  INV_X1 U1964 ( .A(\REGISTERS[31][31] ), .ZN(n2219) );
  INV_X1 U1965 ( .A(\REGISTERS[1][31] ), .ZN(n507) );
  INV_X1 U1966 ( .A(\REGISTERS[5][31] ), .ZN(n1835) );
  INV_X1 U1967 ( .A(\REGISTERS[9][31] ), .ZN(n1899) );
  INV_X1 U1968 ( .A(\REGISTERS[13][31] ), .ZN(n1963) );
  INV_X1 U1969 ( .A(\REGISTERS[16][0] ), .ZN(n2026) );
  INV_X1 U1970 ( .A(\REGISTERS[20][0] ), .ZN(n2090) );
  INV_X1 U1971 ( .A(\REGISTERS[24][0] ), .ZN(n2154) );
  INV_X1 U1972 ( .A(\REGISTERS[30][0] ), .ZN(n2218) );
  INV_X1 U1973 ( .A(\REGISTERS[0][0] ), .ZN(n506) );
  INV_X1 U1974 ( .A(\REGISTERS[4][0] ), .ZN(n1834) );
  INV_X1 U1975 ( .A(\REGISTERS[8][0] ), .ZN(n1898) );
  INV_X1 U1976 ( .A(\REGISTERS[12][0] ), .ZN(n1962) );
  INV_X1 U1977 ( .A(\REGISTERS[16][1] ), .ZN(n2025) );
  INV_X1 U1978 ( .A(\REGISTERS[20][1] ), .ZN(n2089) );
  INV_X1 U1979 ( .A(\REGISTERS[24][1] ), .ZN(n2153) );
  INV_X1 U1980 ( .A(\REGISTERS[30][1] ), .ZN(n2217) );
  INV_X1 U1981 ( .A(\REGISTERS[0][1] ), .ZN(n505) );
  INV_X1 U1982 ( .A(\REGISTERS[4][1] ), .ZN(n1833) );
  INV_X1 U1983 ( .A(\REGISTERS[8][1] ), .ZN(n1897) );
  INV_X1 U1984 ( .A(\REGISTERS[12][1] ), .ZN(n1961) );
  INV_X1 U1985 ( .A(\REGISTERS[16][2] ), .ZN(n2024) );
  INV_X1 U1986 ( .A(\REGISTERS[20][2] ), .ZN(n2088) );
  INV_X1 U1987 ( .A(\REGISTERS[24][2] ), .ZN(n2152) );
  INV_X1 U1988 ( .A(\REGISTERS[30][2] ), .ZN(n2216) );
  INV_X1 U1989 ( .A(\REGISTERS[0][2] ), .ZN(n504) );
  INV_X1 U1990 ( .A(\REGISTERS[4][2] ), .ZN(n1832) );
  INV_X1 U1991 ( .A(\REGISTERS[8][2] ), .ZN(n1896) );
  INV_X1 U1992 ( .A(\REGISTERS[12][2] ), .ZN(n1960) );
  INV_X1 U1993 ( .A(\REGISTERS[16][3] ), .ZN(n2023) );
  INV_X1 U1994 ( .A(\REGISTERS[20][3] ), .ZN(n2087) );
  INV_X1 U1995 ( .A(\REGISTERS[24][3] ), .ZN(n2151) );
  INV_X1 U1996 ( .A(\REGISTERS[30][3] ), .ZN(n2215) );
  INV_X1 U1997 ( .A(\REGISTERS[0][3] ), .ZN(n503) );
  INV_X1 U1998 ( .A(\REGISTERS[4][3] ), .ZN(n1831) );
  INV_X1 U1999 ( .A(\REGISTERS[8][3] ), .ZN(n1895) );
  INV_X1 U2000 ( .A(\REGISTERS[12][3] ), .ZN(n1959) );
  INV_X1 U2001 ( .A(\REGISTERS[16][4] ), .ZN(n2022) );
  INV_X1 U2002 ( .A(\REGISTERS[20][4] ), .ZN(n2086) );
  INV_X1 U2003 ( .A(\REGISTERS[24][4] ), .ZN(n2150) );
  INV_X1 U2004 ( .A(\REGISTERS[30][4] ), .ZN(n2214) );
  INV_X1 U2005 ( .A(\REGISTERS[0][4] ), .ZN(n502) );
  INV_X1 U2006 ( .A(\REGISTERS[4][4] ), .ZN(n1830) );
  INV_X1 U2007 ( .A(\REGISTERS[8][4] ), .ZN(n1894) );
  INV_X1 U2008 ( .A(\REGISTERS[12][4] ), .ZN(n1958) );
  INV_X1 U2009 ( .A(\REGISTERS[16][5] ), .ZN(n2021) );
  INV_X1 U2010 ( .A(\REGISTERS[20][5] ), .ZN(n2085) );
  INV_X1 U2011 ( .A(\REGISTERS[24][5] ), .ZN(n2149) );
  INV_X1 U2012 ( .A(\REGISTERS[30][5] ), .ZN(n2213) );
  INV_X1 U2013 ( .A(\REGISTERS[0][5] ), .ZN(n501) );
  INV_X1 U2014 ( .A(\REGISTERS[4][5] ), .ZN(n1829) );
  INV_X1 U2015 ( .A(\REGISTERS[8][5] ), .ZN(n1893) );
  INV_X1 U2016 ( .A(\REGISTERS[12][5] ), .ZN(n1957) );
  INV_X1 U2017 ( .A(\REGISTERS[16][6] ), .ZN(n2020) );
  INV_X1 U2018 ( .A(\REGISTERS[20][6] ), .ZN(n2084) );
  INV_X1 U2019 ( .A(\REGISTERS[24][6] ), .ZN(n2148) );
  INV_X1 U2020 ( .A(\REGISTERS[30][6] ), .ZN(n2212) );
  INV_X1 U2021 ( .A(\REGISTERS[0][6] ), .ZN(n500) );
  INV_X1 U2022 ( .A(\REGISTERS[4][6] ), .ZN(n1828) );
  INV_X1 U2023 ( .A(\REGISTERS[8][6] ), .ZN(n1892) );
  INV_X1 U2024 ( .A(\REGISTERS[12][6] ), .ZN(n1956) );
  INV_X1 U2025 ( .A(\REGISTERS[16][7] ), .ZN(n2019) );
  INV_X1 U2026 ( .A(\REGISTERS[20][7] ), .ZN(n2083) );
  INV_X1 U2027 ( .A(\REGISTERS[24][7] ), .ZN(n2147) );
  INV_X1 U2028 ( .A(\REGISTERS[30][7] ), .ZN(n2211) );
  INV_X1 U2029 ( .A(\REGISTERS[0][7] ), .ZN(n499) );
  INV_X1 U2030 ( .A(\REGISTERS[4][7] ), .ZN(n1827) );
  INV_X1 U2031 ( .A(\REGISTERS[8][7] ), .ZN(n1891) );
  INV_X1 U2032 ( .A(\REGISTERS[12][7] ), .ZN(n1955) );
  INV_X1 U2033 ( .A(\REGISTERS[16][8] ), .ZN(n2018) );
  INV_X1 U2034 ( .A(\REGISTERS[20][8] ), .ZN(n2082) );
  INV_X1 U2035 ( .A(\REGISTERS[24][8] ), .ZN(n2146) );
  INV_X1 U2036 ( .A(\REGISTERS[30][8] ), .ZN(n2210) );
  INV_X1 U2037 ( .A(\REGISTERS[0][8] ), .ZN(n498) );
  INV_X1 U2038 ( .A(\REGISTERS[4][8] ), .ZN(n1826) );
  INV_X1 U2039 ( .A(\REGISTERS[8][8] ), .ZN(n1890) );
  INV_X1 U2040 ( .A(\REGISTERS[12][8] ), .ZN(n1954) );
  INV_X1 U2041 ( .A(\REGISTERS[16][9] ), .ZN(n2017) );
  INV_X1 U2042 ( .A(\REGISTERS[20][9] ), .ZN(n2081) );
  INV_X1 U2043 ( .A(\REGISTERS[24][9] ), .ZN(n2145) );
  INV_X1 U2044 ( .A(\REGISTERS[30][9] ), .ZN(n2209) );
  INV_X1 U2045 ( .A(\REGISTERS[0][9] ), .ZN(n497) );
  INV_X1 U2046 ( .A(\REGISTERS[4][9] ), .ZN(n1825) );
  INV_X1 U2047 ( .A(\REGISTERS[8][9] ), .ZN(n1889) );
  INV_X1 U2048 ( .A(\REGISTERS[12][9] ), .ZN(n1953) );
  INV_X1 U2049 ( .A(\REGISTERS[16][10] ), .ZN(n2016) );
  INV_X1 U2050 ( .A(\REGISTERS[20][10] ), .ZN(n2080) );
  INV_X1 U2051 ( .A(\REGISTERS[24][10] ), .ZN(n2144) );
  INV_X1 U2052 ( .A(\REGISTERS[30][10] ), .ZN(n2208) );
  INV_X1 U2053 ( .A(\REGISTERS[0][10] ), .ZN(n496) );
  INV_X1 U2054 ( .A(\REGISTERS[4][10] ), .ZN(n1824) );
  INV_X1 U2055 ( .A(\REGISTERS[8][10] ), .ZN(n1888) );
  INV_X1 U2056 ( .A(\REGISTERS[12][10] ), .ZN(n1952) );
  INV_X1 U2057 ( .A(\REGISTERS[16][11] ), .ZN(n2015) );
  INV_X1 U2058 ( .A(\REGISTERS[20][11] ), .ZN(n2079) );
  INV_X1 U2059 ( .A(\REGISTERS[24][11] ), .ZN(n2143) );
  INV_X1 U2060 ( .A(\REGISTERS[30][11] ), .ZN(n2207) );
  INV_X1 U2061 ( .A(\REGISTERS[0][11] ), .ZN(n495) );
  INV_X1 U2062 ( .A(\REGISTERS[4][11] ), .ZN(n1823) );
  INV_X1 U2063 ( .A(\REGISTERS[8][11] ), .ZN(n1887) );
  INV_X1 U2064 ( .A(\REGISTERS[12][11] ), .ZN(n1951) );
  INV_X1 U2065 ( .A(\REGISTERS[16][12] ), .ZN(n2014) );
  INV_X1 U2066 ( .A(\REGISTERS[20][12] ), .ZN(n2078) );
  INV_X1 U2067 ( .A(\REGISTERS[24][12] ), .ZN(n2142) );
  INV_X1 U2068 ( .A(\REGISTERS[30][12] ), .ZN(n2206) );
  INV_X1 U2069 ( .A(\REGISTERS[0][12] ), .ZN(n494) );
  INV_X1 U2070 ( .A(\REGISTERS[4][12] ), .ZN(n1822) );
  INV_X1 U2071 ( .A(\REGISTERS[8][12] ), .ZN(n1886) );
  INV_X1 U2072 ( .A(\REGISTERS[12][12] ), .ZN(n1950) );
  INV_X1 U2073 ( .A(\REGISTERS[16][13] ), .ZN(n2013) );
  INV_X1 U2074 ( .A(\REGISTERS[20][13] ), .ZN(n2077) );
  INV_X1 U2075 ( .A(\REGISTERS[24][13] ), .ZN(n2141) );
  INV_X1 U2076 ( .A(\REGISTERS[30][13] ), .ZN(n2205) );
  INV_X1 U2077 ( .A(\REGISTERS[0][13] ), .ZN(n493) );
  INV_X1 U2078 ( .A(\REGISTERS[4][13] ), .ZN(n1821) );
  INV_X1 U2079 ( .A(\REGISTERS[8][13] ), .ZN(n1885) );
  INV_X1 U2080 ( .A(\REGISTERS[12][13] ), .ZN(n1949) );
  INV_X1 U2081 ( .A(\REGISTERS[16][14] ), .ZN(n2012) );
  INV_X1 U2082 ( .A(\REGISTERS[20][14] ), .ZN(n2076) );
  INV_X1 U2083 ( .A(\REGISTERS[24][14] ), .ZN(n2140) );
  INV_X1 U2084 ( .A(\REGISTERS[30][14] ), .ZN(n2204) );
  INV_X1 U2085 ( .A(\REGISTERS[0][14] ), .ZN(n492) );
  INV_X1 U2086 ( .A(\REGISTERS[4][14] ), .ZN(n1820) );
  INV_X1 U2087 ( .A(\REGISTERS[8][14] ), .ZN(n1884) );
  INV_X1 U2088 ( .A(\REGISTERS[12][14] ), .ZN(n1948) );
  INV_X1 U2089 ( .A(\REGISTERS[16][15] ), .ZN(n2011) );
  INV_X1 U2090 ( .A(\REGISTERS[20][15] ), .ZN(n2075) );
  INV_X1 U2091 ( .A(\REGISTERS[24][15] ), .ZN(n2139) );
  INV_X1 U2092 ( .A(\REGISTERS[30][15] ), .ZN(n2203) );
  INV_X1 U2093 ( .A(\REGISTERS[0][15] ), .ZN(n491) );
  INV_X1 U2094 ( .A(\REGISTERS[4][15] ), .ZN(n1819) );
  INV_X1 U2095 ( .A(\REGISTERS[8][15] ), .ZN(n1883) );
  INV_X1 U2096 ( .A(\REGISTERS[12][15] ), .ZN(n1947) );
  INV_X1 U2097 ( .A(\REGISTERS[16][16] ), .ZN(n2010) );
  INV_X1 U2098 ( .A(\REGISTERS[20][16] ), .ZN(n2074) );
  INV_X1 U2099 ( .A(\REGISTERS[24][16] ), .ZN(n2138) );
  INV_X1 U2100 ( .A(\REGISTERS[30][16] ), .ZN(n2202) );
  INV_X1 U2101 ( .A(\REGISTERS[0][16] ), .ZN(n490) );
  INV_X1 U2102 ( .A(\REGISTERS[4][16] ), .ZN(n1818) );
  INV_X1 U2103 ( .A(\REGISTERS[8][16] ), .ZN(n1882) );
  INV_X1 U2104 ( .A(\REGISTERS[12][16] ), .ZN(n1946) );
  INV_X1 U2105 ( .A(\REGISTERS[16][17] ), .ZN(n2009) );
  INV_X1 U2106 ( .A(\REGISTERS[20][17] ), .ZN(n2073) );
  INV_X1 U2107 ( .A(\REGISTERS[24][17] ), .ZN(n2137) );
  INV_X1 U2108 ( .A(\REGISTERS[30][17] ), .ZN(n2201) );
  INV_X1 U2109 ( .A(\REGISTERS[0][17] ), .ZN(n489) );
  INV_X1 U2110 ( .A(\REGISTERS[4][17] ), .ZN(n1817) );
  INV_X1 U2111 ( .A(\REGISTERS[8][17] ), .ZN(n1881) );
  INV_X1 U2112 ( .A(\REGISTERS[12][17] ), .ZN(n1945) );
  INV_X1 U2113 ( .A(\REGISTERS[16][18] ), .ZN(n2008) );
  INV_X1 U2114 ( .A(\REGISTERS[20][18] ), .ZN(n2072) );
  INV_X1 U2115 ( .A(\REGISTERS[24][18] ), .ZN(n2136) );
  INV_X1 U2116 ( .A(\REGISTERS[30][18] ), .ZN(n2200) );
  INV_X1 U2117 ( .A(\REGISTERS[0][18] ), .ZN(n488) );
  INV_X1 U2118 ( .A(\REGISTERS[4][18] ), .ZN(n1816) );
  INV_X1 U2119 ( .A(\REGISTERS[8][18] ), .ZN(n1880) );
  INV_X1 U2120 ( .A(\REGISTERS[12][18] ), .ZN(n1944) );
  INV_X1 U2121 ( .A(\REGISTERS[16][19] ), .ZN(n2007) );
  INV_X1 U2122 ( .A(\REGISTERS[20][19] ), .ZN(n2071) );
  INV_X1 U2123 ( .A(\REGISTERS[24][19] ), .ZN(n2135) );
  INV_X1 U2124 ( .A(\REGISTERS[30][19] ), .ZN(n2199) );
  INV_X1 U2125 ( .A(\REGISTERS[0][19] ), .ZN(n487) );
  INV_X1 U2126 ( .A(\REGISTERS[4][19] ), .ZN(n1815) );
  INV_X1 U2127 ( .A(\REGISTERS[8][19] ), .ZN(n1879) );
  INV_X1 U2128 ( .A(\REGISTERS[12][19] ), .ZN(n1943) );
  INV_X1 U2129 ( .A(\REGISTERS[16][20] ), .ZN(n2006) );
  INV_X1 U2130 ( .A(\REGISTERS[20][20] ), .ZN(n2070) );
  INV_X1 U2131 ( .A(\REGISTERS[24][20] ), .ZN(n2134) );
  INV_X1 U2132 ( .A(\REGISTERS[30][20] ), .ZN(n2198) );
  INV_X1 U2133 ( .A(\REGISTERS[0][20] ), .ZN(n486) );
  INV_X1 U2134 ( .A(\REGISTERS[4][20] ), .ZN(n1814) );
  INV_X1 U2135 ( .A(\REGISTERS[8][20] ), .ZN(n1878) );
  INV_X1 U2136 ( .A(\REGISTERS[12][20] ), .ZN(n1942) );
  INV_X1 U2137 ( .A(\REGISTERS[16][21] ), .ZN(n2005) );
  INV_X1 U2138 ( .A(\REGISTERS[20][21] ), .ZN(n2069) );
  INV_X1 U2139 ( .A(\REGISTERS[24][21] ), .ZN(n2133) );
  INV_X1 U2140 ( .A(\REGISTERS[30][21] ), .ZN(n2197) );
  INV_X1 U2141 ( .A(\REGISTERS[0][21] ), .ZN(n485) );
  INV_X1 U2142 ( .A(\REGISTERS[4][21] ), .ZN(n1813) );
  INV_X1 U2143 ( .A(\REGISTERS[8][21] ), .ZN(n1877) );
  INV_X1 U2144 ( .A(\REGISTERS[12][21] ), .ZN(n1941) );
  INV_X1 U2145 ( .A(\REGISTERS[16][22] ), .ZN(n2004) );
  INV_X1 U2146 ( .A(\REGISTERS[20][22] ), .ZN(n2068) );
  INV_X1 U2147 ( .A(\REGISTERS[24][22] ), .ZN(n2132) );
  INV_X1 U2148 ( .A(\REGISTERS[30][22] ), .ZN(n2196) );
  INV_X1 U2149 ( .A(\REGISTERS[0][22] ), .ZN(n484) );
  INV_X1 U2150 ( .A(\REGISTERS[4][22] ), .ZN(n1812) );
  INV_X1 U2151 ( .A(\REGISTERS[8][22] ), .ZN(n1876) );
  INV_X1 U2152 ( .A(\REGISTERS[12][22] ), .ZN(n1940) );
  INV_X1 U2153 ( .A(\REGISTERS[16][23] ), .ZN(n2003) );
  INV_X1 U2154 ( .A(\REGISTERS[20][23] ), .ZN(n2067) );
  INV_X1 U2155 ( .A(\REGISTERS[24][23] ), .ZN(n2131) );
  INV_X1 U2156 ( .A(\REGISTERS[30][23] ), .ZN(n2195) );
  INV_X1 U2157 ( .A(\REGISTERS[0][23] ), .ZN(n483) );
  INV_X1 U2158 ( .A(\REGISTERS[4][23] ), .ZN(n1811) );
  INV_X1 U2159 ( .A(\REGISTERS[8][23] ), .ZN(n1875) );
  INV_X1 U2160 ( .A(\REGISTERS[12][23] ), .ZN(n1939) );
  INV_X1 U2161 ( .A(\REGISTERS[16][24] ), .ZN(n2002) );
  INV_X1 U2162 ( .A(\REGISTERS[20][24] ), .ZN(n2066) );
  INV_X1 U2163 ( .A(\REGISTERS[24][24] ), .ZN(n2130) );
  INV_X1 U2164 ( .A(\REGISTERS[30][24] ), .ZN(n2194) );
  INV_X1 U2165 ( .A(\REGISTERS[0][24] ), .ZN(n482) );
  INV_X1 U2166 ( .A(\REGISTERS[4][24] ), .ZN(n1810) );
  INV_X1 U2167 ( .A(\REGISTERS[8][24] ), .ZN(n1874) );
  INV_X1 U2168 ( .A(\REGISTERS[12][24] ), .ZN(n1938) );
  INV_X1 U2169 ( .A(\REGISTERS[16][25] ), .ZN(n2001) );
  INV_X1 U2170 ( .A(\REGISTERS[20][25] ), .ZN(n2065) );
  INV_X1 U2171 ( .A(\REGISTERS[24][25] ), .ZN(n2129) );
  INV_X1 U2172 ( .A(\REGISTERS[30][25] ), .ZN(n2193) );
  INV_X1 U2173 ( .A(\REGISTERS[0][25] ), .ZN(n481) );
  INV_X1 U2174 ( .A(\REGISTERS[4][25] ), .ZN(n1809) );
  INV_X1 U2175 ( .A(\REGISTERS[8][25] ), .ZN(n1873) );
  INV_X1 U2176 ( .A(\REGISTERS[12][25] ), .ZN(n1937) );
  INV_X1 U2177 ( .A(\REGISTERS[16][26] ), .ZN(n2000) );
  INV_X1 U2178 ( .A(\REGISTERS[20][26] ), .ZN(n2064) );
  INV_X1 U2179 ( .A(\REGISTERS[24][26] ), .ZN(n2128) );
  INV_X1 U2180 ( .A(\REGISTERS[30][26] ), .ZN(n2192) );
  INV_X1 U2181 ( .A(\REGISTERS[0][26] ), .ZN(n480) );
  INV_X1 U2182 ( .A(\REGISTERS[4][26] ), .ZN(n1808) );
  INV_X1 U2183 ( .A(\REGISTERS[8][26] ), .ZN(n1872) );
  INV_X1 U2184 ( .A(\REGISTERS[12][26] ), .ZN(n1936) );
  INV_X1 U2185 ( .A(\REGISTERS[16][27] ), .ZN(n1999) );
  INV_X1 U2186 ( .A(\REGISTERS[20][27] ), .ZN(n2063) );
  INV_X1 U2187 ( .A(\REGISTERS[24][27] ), .ZN(n2127) );
  INV_X1 U2188 ( .A(\REGISTERS[30][27] ), .ZN(n2191) );
  INV_X1 U2189 ( .A(\REGISTERS[0][27] ), .ZN(n479) );
  INV_X1 U2190 ( .A(\REGISTERS[4][27] ), .ZN(n1807) );
  INV_X1 U2191 ( .A(\REGISTERS[8][27] ), .ZN(n1871) );
  INV_X1 U2192 ( .A(\REGISTERS[12][27] ), .ZN(n1935) );
  INV_X1 U2193 ( .A(\REGISTERS[16][28] ), .ZN(n1998) );
  INV_X1 U2194 ( .A(\REGISTERS[20][28] ), .ZN(n2062) );
  INV_X1 U2195 ( .A(\REGISTERS[24][28] ), .ZN(n2126) );
  INV_X1 U2196 ( .A(\REGISTERS[30][28] ), .ZN(n2190) );
  INV_X1 U2197 ( .A(\REGISTERS[0][28] ), .ZN(n478) );
  INV_X1 U2198 ( .A(\REGISTERS[4][28] ), .ZN(n1806) );
  INV_X1 U2199 ( .A(\REGISTERS[8][28] ), .ZN(n1870) );
  INV_X1 U2200 ( .A(\REGISTERS[12][28] ), .ZN(n1934) );
  INV_X1 U2201 ( .A(\REGISTERS[16][29] ), .ZN(n1997) );
  INV_X1 U2202 ( .A(\REGISTERS[20][29] ), .ZN(n2061) );
  INV_X1 U2203 ( .A(\REGISTERS[24][29] ), .ZN(n2125) );
  INV_X1 U2204 ( .A(\REGISTERS[30][29] ), .ZN(n2189) );
  INV_X1 U2205 ( .A(\REGISTERS[0][29] ), .ZN(n477) );
  INV_X1 U2206 ( .A(\REGISTERS[4][29] ), .ZN(n1805) );
  INV_X1 U2207 ( .A(\REGISTERS[8][29] ), .ZN(n1869) );
  INV_X1 U2208 ( .A(\REGISTERS[12][29] ), .ZN(n1933) );
  INV_X1 U2209 ( .A(\REGISTERS[16][30] ), .ZN(n1996) );
  INV_X1 U2210 ( .A(\REGISTERS[20][30] ), .ZN(n2060) );
  INV_X1 U2211 ( .A(\REGISTERS[24][30] ), .ZN(n2124) );
  INV_X1 U2212 ( .A(\REGISTERS[30][30] ), .ZN(n2188) );
  INV_X1 U2213 ( .A(\REGISTERS[0][30] ), .ZN(n476) );
  INV_X1 U2214 ( .A(\REGISTERS[4][30] ), .ZN(n1804) );
  INV_X1 U2215 ( .A(\REGISTERS[8][30] ), .ZN(n1868) );
  INV_X1 U2216 ( .A(\REGISTERS[12][30] ), .ZN(n1932) );
  INV_X1 U2217 ( .A(\REGISTERS[16][31] ), .ZN(n1995) );
  INV_X1 U2218 ( .A(\REGISTERS[20][31] ), .ZN(n2059) );
  INV_X1 U2219 ( .A(\REGISTERS[24][31] ), .ZN(n2123) );
  INV_X1 U2220 ( .A(\REGISTERS[30][31] ), .ZN(n2187) );
  INV_X1 U2221 ( .A(\REGISTERS[0][31] ), .ZN(n475) );
  INV_X1 U2222 ( .A(\REGISTERS[4][31] ), .ZN(n1803) );
  INV_X1 U2223 ( .A(\REGISTERS[8][31] ), .ZN(n1867) );
  INV_X1 U2224 ( .A(\REGISTERS[12][31] ), .ZN(n1931) );
  INV_X1 U2225 ( .A(ADD_RD1[2]), .ZN(n2257) );
  NOR2_X1 U2226 ( .A1(n2256), .A2(ADD_RD1[2]), .ZN(n1750) );
  NOR2_X1 U2227 ( .A1(ADD_RD1[1]), .A2(ADD_RD1[2]), .ZN(n1752) );
  CLKBUF_X1 U2228 ( .A(N409), .Z(n196) );
  CLKBUF_X1 U2229 ( .A(N409), .Z(n197) );
  CLKBUF_X1 U2230 ( .A(N409), .Z(n198) );
  CLKBUF_X1 U2231 ( .A(N409), .Z(n199) );
  CLKBUF_X1 U2232 ( .A(N376), .Z(n200) );
  CLKBUF_X1 U2233 ( .A(N376), .Z(n201) );
  CLKBUF_X1 U2234 ( .A(N376), .Z(n202) );
  CLKBUF_X1 U2235 ( .A(N376), .Z(n203) );
  CLKBUF_X1 U2236 ( .A(N375), .Z(n204) );
  CLKBUF_X1 U2237 ( .A(N375), .Z(n205) );
  CLKBUF_X1 U2238 ( .A(N375), .Z(n206) );
  CLKBUF_X1 U2239 ( .A(N375), .Z(n207) );
  CLKBUF_X1 U2240 ( .A(N374), .Z(n208) );
  CLKBUF_X1 U2241 ( .A(N374), .Z(n209) );
  CLKBUF_X1 U2242 ( .A(N374), .Z(n210) );
  CLKBUF_X1 U2243 ( .A(N374), .Z(n211) );
  CLKBUF_X1 U2244 ( .A(N373), .Z(n212) );
  CLKBUF_X1 U2245 ( .A(N373), .Z(n213) );
  CLKBUF_X1 U2246 ( .A(N373), .Z(n214) );
  CLKBUF_X1 U2247 ( .A(N373), .Z(n215) );
  CLKBUF_X1 U2248 ( .A(N372), .Z(n216) );
  CLKBUF_X1 U2249 ( .A(N372), .Z(n217) );
  CLKBUF_X1 U2250 ( .A(N372), .Z(n218) );
  CLKBUF_X1 U2251 ( .A(N372), .Z(n219) );
  CLKBUF_X1 U2252 ( .A(N371), .Z(n220) );
  CLKBUF_X1 U2253 ( .A(N371), .Z(n221) );
  CLKBUF_X1 U2254 ( .A(N371), .Z(n222) );
  CLKBUF_X1 U2255 ( .A(N371), .Z(n223) );
  CLKBUF_X1 U2256 ( .A(N370), .Z(n224) );
  CLKBUF_X1 U2257 ( .A(N370), .Z(n225) );
  CLKBUF_X1 U2258 ( .A(N370), .Z(n226) );
  CLKBUF_X1 U2259 ( .A(N370), .Z(n227) );
  CLKBUF_X1 U2260 ( .A(N369), .Z(n228) );
  CLKBUF_X1 U2261 ( .A(N369), .Z(n229) );
  CLKBUF_X1 U2262 ( .A(N369), .Z(n230) );
  CLKBUF_X1 U2263 ( .A(N369), .Z(n231) );
  CLKBUF_X1 U2264 ( .A(N368), .Z(n232) );
  CLKBUF_X1 U2265 ( .A(N368), .Z(n233) );
  CLKBUF_X1 U2266 ( .A(N368), .Z(n234) );
  CLKBUF_X1 U2267 ( .A(N368), .Z(n235) );
  CLKBUF_X1 U2268 ( .A(N367), .Z(n236) );
  CLKBUF_X1 U2269 ( .A(N367), .Z(n237) );
  CLKBUF_X1 U2270 ( .A(N367), .Z(n238) );
  CLKBUF_X1 U2271 ( .A(N367), .Z(n239) );
  CLKBUF_X1 U2272 ( .A(N366), .Z(n240) );
  CLKBUF_X1 U2273 ( .A(N366), .Z(n241) );
  CLKBUF_X1 U2274 ( .A(N366), .Z(n242) );
  CLKBUF_X1 U2275 ( .A(N366), .Z(n243) );
  CLKBUF_X1 U2276 ( .A(N365), .Z(n244) );
  CLKBUF_X1 U2277 ( .A(N365), .Z(n245) );
  CLKBUF_X1 U2278 ( .A(N365), .Z(n246) );
  CLKBUF_X1 U2279 ( .A(N365), .Z(n247) );
  CLKBUF_X1 U2280 ( .A(N364), .Z(n248) );
  CLKBUF_X1 U2281 ( .A(N364), .Z(n249) );
  CLKBUF_X1 U2282 ( .A(N364), .Z(n250) );
  CLKBUF_X1 U2283 ( .A(N364), .Z(n251) );
  CLKBUF_X1 U2284 ( .A(N363), .Z(n252) );
  CLKBUF_X1 U2285 ( .A(N363), .Z(n253) );
  CLKBUF_X1 U2286 ( .A(N363), .Z(n254) );
  CLKBUF_X1 U2287 ( .A(N363), .Z(n255) );
  CLKBUF_X1 U2288 ( .A(N362), .Z(n256) );
  CLKBUF_X1 U2289 ( .A(N362), .Z(n257) );
  CLKBUF_X1 U2290 ( .A(N362), .Z(n258) );
  CLKBUF_X1 U2291 ( .A(N362), .Z(n259) );
  CLKBUF_X1 U2292 ( .A(N361), .Z(n260) );
  CLKBUF_X1 U2293 ( .A(N361), .Z(n261) );
  CLKBUF_X1 U2294 ( .A(N361), .Z(n262) );
  CLKBUF_X1 U2295 ( .A(N361), .Z(n263) );
  CLKBUF_X1 U2296 ( .A(N360), .Z(n264) );
  CLKBUF_X1 U2297 ( .A(N360), .Z(n265) );
  CLKBUF_X1 U2298 ( .A(N360), .Z(n266) );
  CLKBUF_X1 U2299 ( .A(N360), .Z(n267) );
  CLKBUF_X1 U2300 ( .A(N359), .Z(n268) );
  CLKBUF_X1 U2301 ( .A(N359), .Z(n269) );
  CLKBUF_X1 U2302 ( .A(N359), .Z(n270) );
  CLKBUF_X1 U2303 ( .A(N359), .Z(n271) );
  CLKBUF_X1 U2304 ( .A(N358), .Z(n272) );
  CLKBUF_X1 U2305 ( .A(N358), .Z(n273) );
  CLKBUF_X1 U2306 ( .A(N358), .Z(n274) );
  CLKBUF_X1 U2307 ( .A(N358), .Z(n275) );
  CLKBUF_X1 U2308 ( .A(N357), .Z(n276) );
  CLKBUF_X1 U2309 ( .A(N357), .Z(n277) );
  CLKBUF_X1 U2310 ( .A(N357), .Z(n278) );
  CLKBUF_X1 U2311 ( .A(N357), .Z(n279) );
  CLKBUF_X1 U2312 ( .A(N356), .Z(n280) );
  CLKBUF_X1 U2313 ( .A(N356), .Z(n281) );
  CLKBUF_X1 U2314 ( .A(N356), .Z(n282) );
  CLKBUF_X1 U2315 ( .A(N356), .Z(n283) );
  CLKBUF_X1 U2316 ( .A(N355), .Z(n284) );
  CLKBUF_X1 U2317 ( .A(N355), .Z(n285) );
  CLKBUF_X1 U2318 ( .A(N355), .Z(n286) );
  CLKBUF_X1 U2319 ( .A(N355), .Z(n287) );
  CLKBUF_X1 U2320 ( .A(N354), .Z(n288) );
  CLKBUF_X1 U2321 ( .A(N354), .Z(n289) );
  CLKBUF_X1 U2322 ( .A(N354), .Z(n290) );
  CLKBUF_X1 U2323 ( .A(N354), .Z(n291) );
  CLKBUF_X1 U2324 ( .A(N353), .Z(n292) );
  CLKBUF_X1 U2325 ( .A(N353), .Z(n293) );
  CLKBUF_X1 U2326 ( .A(N353), .Z(n294) );
  CLKBUF_X1 U2327 ( .A(N353), .Z(n295) );
  CLKBUF_X1 U2328 ( .A(N352), .Z(n296) );
  CLKBUF_X1 U2329 ( .A(N352), .Z(n297) );
  CLKBUF_X1 U2330 ( .A(N352), .Z(n298) );
  CLKBUF_X1 U2331 ( .A(N352), .Z(n299) );
  CLKBUF_X1 U2332 ( .A(N351), .Z(n300) );
  CLKBUF_X1 U2333 ( .A(N351), .Z(n301) );
  CLKBUF_X1 U2334 ( .A(N351), .Z(n302) );
  CLKBUF_X1 U2335 ( .A(N351), .Z(n303) );
  CLKBUF_X1 U2336 ( .A(N350), .Z(n304) );
  CLKBUF_X1 U2337 ( .A(N350), .Z(n305) );
  CLKBUF_X1 U2338 ( .A(N350), .Z(n306) );
  CLKBUF_X1 U2339 ( .A(N350), .Z(n307) );
  CLKBUF_X1 U2340 ( .A(N349), .Z(n308) );
  CLKBUF_X1 U2341 ( .A(N349), .Z(n309) );
  CLKBUF_X1 U2342 ( .A(N349), .Z(n310) );
  CLKBUF_X1 U2343 ( .A(N349), .Z(n311) );
  CLKBUF_X1 U2344 ( .A(N348), .Z(n312) );
  CLKBUF_X1 U2345 ( .A(N348), .Z(n313) );
  CLKBUF_X1 U2346 ( .A(N348), .Z(n314) );
  CLKBUF_X1 U2347 ( .A(N348), .Z(n315) );
  CLKBUF_X1 U2348 ( .A(N347), .Z(n316) );
  CLKBUF_X1 U2349 ( .A(N347), .Z(n317) );
  CLKBUF_X1 U2350 ( .A(N347), .Z(n318) );
  CLKBUF_X1 U2351 ( .A(N347), .Z(n319) );
  CLKBUF_X1 U2352 ( .A(N346), .Z(n320) );
  CLKBUF_X1 U2353 ( .A(N346), .Z(n321) );
  CLKBUF_X1 U2354 ( .A(N346), .Z(n322) );
  CLKBUF_X1 U2355 ( .A(N346), .Z(n323) );
  CLKBUF_X1 U2356 ( .A(N345), .Z(n324) );
  CLKBUF_X1 U2357 ( .A(N345), .Z(n325) );
  CLKBUF_X1 U2358 ( .A(N345), .Z(n326) );
  CLKBUF_X1 U2359 ( .A(N345), .Z(n327) );
  CLKBUF_X1 U2360 ( .A(N344), .Z(n331) );
  CLKBUF_X1 U2361 ( .A(N343), .Z(n335) );
  CLKBUF_X1 U2362 ( .A(N342), .Z(n339) );
  CLKBUF_X1 U2363 ( .A(N341), .Z(n343) );
  CLKBUF_X1 U2364 ( .A(N340), .Z(n347) );
  CLKBUF_X1 U2365 ( .A(N339), .Z(n351) );
  CLKBUF_X1 U2366 ( .A(N338), .Z(n355) );
  CLKBUF_X1 U2367 ( .A(N337), .Z(n359) );
  CLKBUF_X1 U2368 ( .A(N336), .Z(n363) );
  CLKBUF_X1 U2369 ( .A(N335), .Z(n367) );
  CLKBUF_X1 U2370 ( .A(N334), .Z(n371) );
  CLKBUF_X1 U2371 ( .A(N333), .Z(n375) );
  CLKBUF_X1 U2372 ( .A(N332), .Z(n379) );
  CLKBUF_X1 U2373 ( .A(N331), .Z(n383) );
  CLKBUF_X1 U2374 ( .A(N330), .Z(n387) );
  CLKBUF_X1 U2375 ( .A(N329), .Z(n391) );
  CLKBUF_X1 U2376 ( .A(N328), .Z(n395) );
  CLKBUF_X1 U2377 ( .A(N327), .Z(n399) );
  CLKBUF_X1 U2378 ( .A(N326), .Z(n403) );
  CLKBUF_X1 U2379 ( .A(N325), .Z(n407) );
  CLKBUF_X1 U2380 ( .A(N324), .Z(n411) );
  CLKBUF_X1 U2381 ( .A(N323), .Z(n415) );
  CLKBUF_X1 U2382 ( .A(N322), .Z(n419) );
  CLKBUF_X1 U2383 ( .A(N321), .Z(n423) );
  CLKBUF_X1 U2384 ( .A(N320), .Z(n427) );
  CLKBUF_X1 U2385 ( .A(N319), .Z(n431) );
  CLKBUF_X1 U2386 ( .A(N318), .Z(n435) );
  CLKBUF_X1 U2387 ( .A(N317), .Z(n439) );
  CLKBUF_X1 U2388 ( .A(N316), .Z(n443) );
  CLKBUF_X1 U2389 ( .A(N315), .Z(n447) );
  CLKBUF_X1 U2390 ( .A(N314), .Z(n451) );
  CLKBUF_X1 U2391 ( .A(N313), .Z(n455) );
  CLKBUF_X1 U2392 ( .A(N312), .Z(n456) );
  CLKBUF_X1 U2393 ( .A(N312), .Z(n457) );
  CLKBUF_X1 U2394 ( .A(N312), .Z(n458) );
  CLKBUF_X1 U2395 ( .A(N312), .Z(n459) );
endmodule


module DEC ( instr, RST, RFdata_in, RFWA, NPC_in, EXE_RD, Ld, ALU_regout, 
        MEM_RD, WB_RD, RD_inmul, flag_structHzd, flag_ismul, RF1, RF2, WF1, 
        EN1, opcode, func, IMM, RA, RB, RSA, RSB, RD, stall_NPC, PC_sel, 
        dec_flag, NPC_jump );
  input [31:0] instr;
  input [31:0] RFdata_in;
  input [4:0] RFWA;
  input [31:0] NPC_in;
  input [4:0] EXE_RD;
  input [31:0] ALU_regout;
  input [4:0] MEM_RD;
  input [4:0] WB_RD;
  input [4:0] RD_inmul;
  output [5:0] opcode;
  output [10:0] func;
  output [31:0] IMM;
  output [31:0] RA;
  output [31:0] RB;
  output [4:0] RSA;
  output [4:0] RSB;
  output [4:0] RD;
  output [31:0] stall_NPC;
  output [31:0] NPC_jump;
  input RST, Ld, flag_structHzd, flag_ismul, RF1, RF2, WF1, EN1;
  output PC_sel, dec_flag;
  wire   mux_select, n3, n4, n5, n6, n7, n1, n2, n8, n9;
  wire   [5:0] s_opcode;
  wire   [10:0] s_FUNC;
  wire   [4:0] s_RD;
  wire   [25:0] s_IMM26;
  wire   [31:0] adder_out;
  wire   [31:0] s_Rega_new;
  assign IMM[16] = IMM[31];
  assign IMM[17] = IMM[31];
  assign IMM[18] = IMM[31];
  assign IMM[19] = IMM[31];
  assign IMM[20] = IMM[31];
  assign IMM[21] = IMM[31];
  assign IMM[22] = IMM[31];
  assign IMM[23] = IMM[31];
  assign IMM[24] = IMM[31];
  assign IMM[25] = IMM[31];
  assign IMM[26] = IMM[31];
  assign IMM[27] = IMM[31];
  assign IMM[28] = IMM[31];
  assign IMM[29] = IMM[31];
  assign IMM[30] = IMM[31];

  dec_logic_WORD_size32_NREG32 decode_logic ( .instr(instr), .NPC_in(NPC_in), 
        .opcode(s_opcode), .RS1(RSA), .RS2(RSB), .RD(s_RD), .FUNC(s_FUNC), 
        .IMM(IMM[15:0]), .IMM26(s_IMM26) );
  P4_ADDER_NBIT32_0 jump_npc_adder ( .A({n1, n1, n1, n1, n1, n2, n2, 
        s_IMM26[24:0]}), .B(NPC_in), .Cin(1'b0), .S(adder_out) );
  jump_logic_WORD_size32_NREG32_reg_file_size32 jmp_logic ( .opcode(opcode), 
        .RSA(RSA), .WB_RD(WB_RD), .MEM_RD(MEM_RD), .Rega(RA), .ALU_out(
        ALU_regout), .MEM_out(RFdata_in), .Rega_new(s_Rega_new), .mux_s(
        mux_select), .flag(dec_flag) );
  MUX21_GENERIC_NBIT32_3 MUX ( .A(adder_out), .B(s_Rega_new), .SEL(mux_select), 
        .Y(NPC_jump) );
  stall_detection_unit_op_code_size6_func_size11_PC_reg_size32_reg_file_size32 SDU ( 
        .opcode(s_opcode), .RSA(RSA), .RSB(RSB), .RD(s_RD), .FUNC(s_FUNC), 
        .EXE_RD(EXE_RD), .NPC_in(NPC_in), .Ld(Ld), .RD_inmul(RD_inmul), 
        .flag_structHzd(flag_structHzd), .flag_ismul(flag_ismul), .opcode_out(
        opcode), .RD_out(RD), .FUNC_out(func), .NPC_out(stall_NPC), .PC_sel(
        PC_sel) );
  register_file_NBIT32_NREG32 REG_FILE ( .RESET(RST), .ENABLE(EN1), .RD1(RF1), 
        .RD2(RF2), .WR(WF1), .ADD_WR(RFWA), .ADD_RD1(RSA), .ADD_RD2(RSB), 
        .DATAIN(RFdata_in), .OUT1(RA), .OUT2(RB) );
  AND2_X1 U2 ( .A1(IMM[15]), .A2(n3), .ZN(IMM[31]) );
  NAND4_X1 U3 ( .A1(n4), .A2(s_opcode[3]), .A3(n5), .A4(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(n7), .A2(n8), .ZN(n5) );
  INV_X1 U5 ( .A(s_opcode[2]), .ZN(n8) );
  BUF_X2 U6 ( .A(s_IMM26[25]), .Z(n1) );
  BUF_X1 U7 ( .A(s_IMM26[25]), .Z(n2) );
  XNOR2_X1 U8 ( .A(s_opcode[4]), .B(s_opcode[5]), .ZN(n4) );
  OAI211_X1 U9 ( .C1(s_opcode[0]), .C2(s_opcode[4]), .A(s_opcode[1]), .B(
        s_opcode[2]), .ZN(n6) );
  OAI22_X1 U10 ( .A1(s_opcode[0]), .A2(s_opcode[4]), .B1(s_opcode[1]), .B2(n9), 
        .ZN(n7) );
  INV_X1 U11 ( .A(s_opcode[4]), .ZN(n9) );
endmodule


module forwarding_unit_WORD_size32_NREG32 ( RSA, RSB, ALU_outmem, WB_out, 
        MEM_RD, WB_RD, LD_EN, WB_EN, S1, S2, SEL1, SEL2, SEL3 );
  input [4:0] RSA;
  input [4:0] RSB;
  input [31:0] ALU_outmem;
  input [31:0] WB_out;
  input [4:0] MEM_RD;
  input [4:0] WB_RD;
  output [1:0] SEL1;
  output [1:0] SEL2;
  output [1:0] SEL3;
  input LD_EN, WB_EN, S1, S2;
  wire   N30, N31, N32, N49, N50, N51, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44;

  DLH_X1 \SEL1_reg[1]  ( .G(N30), .D(N32), .Q(SEL1[1]) );
  DLH_X1 \SEL1_reg[0]  ( .G(N30), .D(N31), .Q(SEL1[0]) );
  DLH_X1 \SEL2_reg[1]  ( .G(N49), .D(N51), .Q(SEL2[1]) );
  DLH_X1 \SEL2_reg[0]  ( .G(N49), .D(N50), .Q(SEL2[0]) );
  NAND2_X1 U3 ( .A1(SEL3[0]), .A2(n1), .ZN(SEL3[1]) );
  NAND3_X1 U4 ( .A1(n2), .A2(n3), .A3(WB_EN), .ZN(n1) );
  INV_X1 U5 ( .A(n4), .ZN(N50) );
  AOI21_X1 U6 ( .B1(SEL3[0]), .B2(n5), .A(S2), .ZN(n4) );
  INV_X1 U7 ( .A(n6), .ZN(n5) );
  OAI211_X1 U8 ( .C1(n7), .C2(n8), .A(SEL3[0]), .B(N51), .ZN(N49) );
  NOR2_X1 U9 ( .A1(n6), .A2(S2), .ZN(N51) );
  OAI21_X1 U10 ( .B1(n9), .B2(n2), .A(n3), .ZN(n6) );
  INV_X1 U11 ( .A(n7), .ZN(n2) );
  NAND3_X1 U12 ( .A1(n3), .A2(n10), .A3(n9), .ZN(SEL3[0]) );
  AND4_X1 U13 ( .A1(n11), .A2(n12), .A3(n13), .A4(n14), .ZN(n9) );
  NOR2_X1 U14 ( .A1(n15), .A2(n16), .ZN(n14) );
  XOR2_X1 U15 ( .A(RSB[4]), .B(MEM_RD[4]), .Z(n16) );
  XOR2_X1 U16 ( .A(RSB[3]), .B(MEM_RD[3]), .Z(n15) );
  XNOR2_X1 U17 ( .A(MEM_RD[1]), .B(RSB[1]), .ZN(n13) );
  XNOR2_X1 U18 ( .A(MEM_RD[2]), .B(RSB[2]), .ZN(n12) );
  XNOR2_X1 U19 ( .A(MEM_RD[0]), .B(RSB[0]), .ZN(n11) );
  INV_X1 U20 ( .A(LD_EN), .ZN(n10) );
  OR4_X1 U21 ( .A1(RSB[3]), .A2(RSB[4]), .A3(RSB[2]), .A4(n17), .ZN(n3) );
  OR2_X1 U22 ( .A1(RSB[1]), .A2(RSB[0]), .ZN(n17) );
  NAND4_X1 U23 ( .A1(n18), .A2(n19), .A3(n20), .A4(n21), .ZN(n7) );
  NOR2_X1 U24 ( .A1(n22), .A2(n23), .ZN(n21) );
  XOR2_X1 U25 ( .A(WB_RD[4]), .B(RSB[4]), .Z(n23) );
  XOR2_X1 U26 ( .A(WB_RD[3]), .B(RSB[3]), .Z(n22) );
  XNOR2_X1 U27 ( .A(RSB[1]), .B(WB_RD[1]), .ZN(n20) );
  XNOR2_X1 U28 ( .A(RSB[2]), .B(WB_RD[2]), .ZN(n19) );
  XNOR2_X1 U29 ( .A(RSB[0]), .B(WB_RD[0]), .ZN(n18) );
  AOI21_X1 U30 ( .B1(n24), .B2(n25), .A(n26), .ZN(N31) );
  INV_X1 U31 ( .A(n27), .ZN(n25) );
  NOR2_X1 U32 ( .A1(LD_EN), .A2(n28), .ZN(n24) );
  OAI221_X1 U33 ( .B1(LD_EN), .B2(n27), .C1(n8), .C2(n29), .A(N32), .ZN(N30)
         );
  NOR2_X1 U34 ( .A1(n26), .A2(n28), .ZN(N32) );
  INV_X1 U35 ( .A(n30), .ZN(n28) );
  AOI21_X1 U36 ( .B1(n27), .B2(n29), .A(n31), .ZN(n30) );
  NOR4_X1 U37 ( .A1(RSA[3]), .A2(RSA[4]), .A3(RSA[2]), .A4(n32), .ZN(n31) );
  OR2_X1 U38 ( .A1(RSA[1]), .A2(RSA[0]), .ZN(n32) );
  INV_X1 U39 ( .A(S1), .ZN(n26) );
  NAND4_X1 U40 ( .A1(n33), .A2(n34), .A3(n35), .A4(n36), .ZN(n29) );
  NOR2_X1 U41 ( .A1(n37), .A2(n38), .ZN(n36) );
  XOR2_X1 U42 ( .A(WB_RD[4]), .B(RSA[4]), .Z(n38) );
  XOR2_X1 U43 ( .A(WB_RD[3]), .B(RSA[3]), .Z(n37) );
  XNOR2_X1 U44 ( .A(RSA[1]), .B(WB_RD[1]), .ZN(n35) );
  XNOR2_X1 U45 ( .A(RSA[2]), .B(WB_RD[2]), .ZN(n34) );
  XNOR2_X1 U46 ( .A(RSA[0]), .B(WB_RD[0]), .ZN(n33) );
  INV_X1 U47 ( .A(WB_EN), .ZN(n8) );
  NAND4_X1 U48 ( .A1(n39), .A2(n40), .A3(n41), .A4(n42), .ZN(n27) );
  NOR2_X1 U49 ( .A1(n43), .A2(n44), .ZN(n42) );
  XOR2_X1 U50 ( .A(RSA[4]), .B(MEM_RD[4]), .Z(n44) );
  XOR2_X1 U51 ( .A(RSA[3]), .B(MEM_RD[3]), .Z(n43) );
  XNOR2_X1 U52 ( .A(MEM_RD[1]), .B(RSA[1]), .ZN(n41) );
  XNOR2_X1 U53 ( .A(MEM_RD[2]), .B(RSA[2]), .ZN(n40) );
  XNOR2_X1 U54 ( .A(MEM_RD[0]), .B(RSA[0]), .ZN(n39) );
endmodule


module MUX41_0 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n3, n4, n5, n6, n7, n1, n2;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n6) );
  OAI211_X4 U1 ( .C1(n3), .C2(n4), .A(n5), .B(n6), .ZN(Y) );
  NOR2_X1 U2 ( .A1(S[0]), .A2(n2), .ZN(n7) );
  NOR2_X1 U3 ( .A1(n1), .A2(S[1]), .ZN(n3) );
  NAND2_X1 U4 ( .A1(B), .A2(n3), .ZN(n5) );
  AOI22_X1 U5 ( .A1(D), .A2(S[0]), .B1(n7), .B2(C), .ZN(n4) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_167 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  OAI211_X4 U1 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NOR2_X1 U2 ( .A1(n1), .A2(n8), .ZN(n9) );
  NOR2_X1 U3 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  NAND2_X1 U4 ( .A1(B), .A2(n13), .ZN(n11) );
  AOI22_X1 U5 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_166 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  OAI211_X4 U1 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NOR2_X1 U2 ( .A1(n1), .A2(n8), .ZN(n9) );
  NOR2_X1 U3 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  NAND2_X1 U4 ( .A1(B), .A2(n13), .ZN(n11) );
  AOI22_X1 U5 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_165 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  OAI211_X4 U1 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NOR2_X1 U2 ( .A1(n1), .A2(n8), .ZN(n9) );
  NOR2_X1 U3 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  NAND2_X1 U4 ( .A1(B), .A2(n13), .ZN(n11) );
  AOI22_X1 U5 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_164 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  OAI211_X4 U1 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NOR2_X1 U2 ( .A1(n1), .A2(n8), .ZN(n9) );
  NOR2_X1 U3 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  NAND2_X1 U4 ( .A1(B), .A2(n13), .ZN(n11) );
  AOI22_X1 U5 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_163 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  OAI211_X4 U1 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NOR2_X1 U2 ( .A1(n1), .A2(n8), .ZN(n9) );
  NOR2_X1 U3 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  NAND2_X1 U4 ( .A1(B), .A2(n13), .ZN(n11) );
  AOI22_X1 U5 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_162 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  OAI211_X4 U1 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NOR2_X1 U2 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  NOR2_X1 U3 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U5 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_161 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  OAI211_X4 U1 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NOR2_X1 U2 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  NOR2_X1 U3 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U5 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_160 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  OAI211_X2 U1 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  NOR2_X1 U2 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  NOR2_X1 U3 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U5 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_159 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  OAI211_X2 U1 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  NOR2_X1 U2 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  NOR2_X1 U3 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U5 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_158 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  OAI211_X2 U1 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  NOR2_X1 U2 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  NOR2_X1 U3 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U5 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_157 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  OAI211_X2 U1 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  NOR2_X1 U2 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  NOR2_X1 U3 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U5 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_156 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  OAI211_X2 U1 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  NOR2_X1 U2 ( .A1(n1), .A2(n8), .ZN(n9) );
  NOR2_X1 U3 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  NAND2_X1 U4 ( .A1(B), .A2(n13), .ZN(n11) );
  AOI22_X1 U5 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_155 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  OAI211_X2 U1 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  NOR2_X1 U2 ( .A1(n1), .A2(n8), .ZN(n9) );
  NOR2_X1 U3 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  NAND2_X1 U4 ( .A1(B), .A2(n13), .ZN(n11) );
  AOI22_X1 U5 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_154 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  OAI211_X2 U1 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  NOR2_X1 U2 ( .A1(n1), .A2(n8), .ZN(n9) );
  NOR2_X1 U3 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  NAND2_X1 U4 ( .A1(B), .A2(n13), .ZN(n11) );
  AOI22_X1 U5 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_153 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  OAI211_X2 U1 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  NOR2_X1 U2 ( .A1(n1), .A2(n8), .ZN(n9) );
  NOR2_X1 U3 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  NAND2_X1 U4 ( .A1(B), .A2(n13), .ZN(n11) );
  AOI22_X1 U5 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_152 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  OAI211_X2 U1 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  NOR2_X1 U2 ( .A1(n1), .A2(n8), .ZN(n9) );
  NOR2_X1 U3 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  NAND2_X1 U4 ( .A1(B), .A2(n13), .ZN(n11) );
  AOI22_X1 U5 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_151 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  OAI211_X2 U1 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  NOR2_X1 U2 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  NOR2_X1 U3 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U5 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_150 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  OAI211_X2 U1 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  NOR2_X1 U2 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  NOR2_X1 U3 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U5 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_149 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  OAI211_X2 U1 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  NOR2_X1 U2 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  NOR2_X1 U3 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U5 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_148 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  OAI211_X2 U1 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  NOR2_X1 U2 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  NOR2_X1 U3 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U5 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_147 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  OAI211_X2 U1 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  NOR2_X1 U2 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  NOR2_X1 U3 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U5 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_146 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  OAI211_X2 U1 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  NOR2_X1 U2 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  NOR2_X1 U3 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U5 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_145 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  OAI211_X2 U1 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  NOR2_X1 U2 ( .A1(n1), .A2(n8), .ZN(n9) );
  NOR2_X1 U3 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  NAND2_X1 U4 ( .A1(B), .A2(n13), .ZN(n11) );
  AOI22_X1 U5 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_144 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  OAI211_X4 U1 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NOR2_X1 U2 ( .A1(n1), .A2(n8), .ZN(n9) );
  NOR2_X1 U3 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  NAND2_X1 U4 ( .A1(B), .A2(n13), .ZN(n11) );
  AOI22_X1 U5 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_143 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  OAI211_X4 U1 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NOR2_X1 U2 ( .A1(n1), .A2(n8), .ZN(n9) );
  NOR2_X1 U3 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  NAND2_X1 U4 ( .A1(B), .A2(n13), .ZN(n11) );
  AOI22_X1 U5 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_142 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  OAI211_X4 U1 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NOR2_X1 U2 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  NOR2_X1 U3 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U5 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_141 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  OAI211_X4 U1 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NOR2_X1 U2 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  NOR2_X1 U3 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U5 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_140 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  OAI211_X4 U1 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NOR2_X1 U2 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  NOR2_X1 U3 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U5 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_139 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  OAI211_X2 U1 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  NOR2_X1 U2 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  NOR2_X1 U3 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U5 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_138 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  OAI211_X2 U1 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  NOR2_X1 U2 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  NOR2_X1 U3 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U5 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_137 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  NOR2_X1 U1 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  NOR2_X1 U2 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  OAI211_X1 U3 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U5 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_GENERIC_NBIT32_0 ( A, B, C, D, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [31:0] D;
  input [1:0] SEL;
  output [31:0] Y;
  wire   n1, n2, n3, n4, n5, n6;

  MUX41_0 MUXES_0 ( .A(A[0]), .B(B[0]), .C(C[0]), .D(D[0]), .S({n6, n3}), .Y(
        Y[0]) );
  MUX41_167 MUXES_1 ( .A(A[1]), .B(B[1]), .C(C[1]), .D(D[1]), .S({n4, n1}), 
        .Y(Y[1]) );
  MUX41_166 MUXES_2 ( .A(A[2]), .B(B[2]), .C(C[2]), .D(D[2]), .S({n4, n1}), 
        .Y(Y[2]) );
  MUX41_165 MUXES_3 ( .A(A[3]), .B(B[3]), .C(C[3]), .D(D[3]), .S({n4, n1}), 
        .Y(Y[3]) );
  MUX41_164 MUXES_4 ( .A(A[4]), .B(B[4]), .C(C[4]), .D(D[4]), .S({n4, n1}), 
        .Y(Y[4]) );
  MUX41_163 MUXES_5 ( .A(A[5]), .B(B[5]), .C(C[5]), .D(D[5]), .S({n4, n1}), 
        .Y(Y[5]) );
  MUX41_162 MUXES_6 ( .A(A[6]), .B(B[6]), .C(C[6]), .D(D[6]), .S({n4, n1}), 
        .Y(Y[6]) );
  MUX41_161 MUXES_7 ( .A(A[7]), .B(B[7]), .C(C[7]), .D(D[7]), .S({n4, n1}), 
        .Y(Y[7]) );
  MUX41_160 MUXES_8 ( .A(A[8]), .B(B[8]), .C(C[8]), .D(D[8]), .S({n4, n1}), 
        .Y(Y[8]) );
  MUX41_159 MUXES_9 ( .A(A[9]), .B(B[9]), .C(C[9]), .D(D[9]), .S({n4, n1}), 
        .Y(Y[9]) );
  MUX41_158 MUXES_10 ( .A(A[10]), .B(B[10]), .C(C[10]), .D(D[10]), .S({n4, n1}), .Y(Y[10]) );
  MUX41_157 MUXES_11 ( .A(A[11]), .B(B[11]), .C(C[11]), .D(D[11]), .S({n4, n1}), .Y(Y[11]) );
  MUX41_156 MUXES_12 ( .A(A[12]), .B(B[12]), .C(C[12]), .D(D[12]), .S({n4, n2}), .Y(Y[12]) );
  MUX41_155 MUXES_13 ( .A(A[13]), .B(B[13]), .C(C[13]), .D(D[13]), .S({n5, n2}), .Y(Y[13]) );
  MUX41_154 MUXES_14 ( .A(A[14]), .B(B[14]), .C(C[14]), .D(D[14]), .S({n5, n2}), .Y(Y[14]) );
  MUX41_153 MUXES_15 ( .A(A[15]), .B(B[15]), .C(C[15]), .D(D[15]), .S({n5, n2}), .Y(Y[15]) );
  MUX41_152 MUXES_16 ( .A(A[16]), .B(B[16]), .C(C[16]), .D(D[16]), .S({n5, n2}), .Y(Y[16]) );
  MUX41_151 MUXES_17 ( .A(A[17]), .B(B[17]), .C(C[17]), .D(D[17]), .S({n5, n2}), .Y(Y[17]) );
  MUX41_150 MUXES_18 ( .A(A[18]), .B(B[18]), .C(C[18]), .D(D[18]), .S({n5, n2}), .Y(Y[18]) );
  MUX41_149 MUXES_19 ( .A(A[19]), .B(B[19]), .C(C[19]), .D(D[19]), .S({n5, n2}), .Y(Y[19]) );
  MUX41_148 MUXES_20 ( .A(A[20]), .B(B[20]), .C(C[20]), .D(D[20]), .S({n5, n2}), .Y(Y[20]) );
  MUX41_147 MUXES_21 ( .A(A[21]), .B(B[21]), .C(C[21]), .D(D[21]), .S({n5, n2}), .Y(Y[21]) );
  MUX41_146 MUXES_22 ( .A(A[22]), .B(B[22]), .C(C[22]), .D(D[22]), .S({n5, n2}), .Y(Y[22]) );
  MUX41_145 MUXES_23 ( .A(A[23]), .B(B[23]), .C(C[23]), .D(D[23]), .S({n5, n3}), .Y(Y[23]) );
  MUX41_144 MUXES_24 ( .A(A[24]), .B(B[24]), .C(C[24]), .D(D[24]), .S({n5, n3}), .Y(Y[24]) );
  MUX41_143 MUXES_25 ( .A(A[25]), .B(B[25]), .C(C[25]), .D(D[25]), .S({n6, n3}), .Y(Y[25]) );
  MUX41_142 MUXES_26 ( .A(A[26]), .B(B[26]), .C(C[26]), .D(D[26]), .S({n6, n3}), .Y(Y[26]) );
  MUX41_141 MUXES_27 ( .A(A[27]), .B(B[27]), .C(C[27]), .D(D[27]), .S({n6, n3}), .Y(Y[27]) );
  MUX41_140 MUXES_28 ( .A(A[28]), .B(B[28]), .C(C[28]), .D(D[28]), .S({n6, n3}), .Y(Y[28]) );
  MUX41_139 MUXES_29 ( .A(A[29]), .B(B[29]), .C(C[29]), .D(D[29]), .S({n6, n3}), .Y(Y[29]) );
  MUX41_138 MUXES_30 ( .A(A[30]), .B(B[30]), .C(C[30]), .D(D[30]), .S({n6, n3}), .Y(Y[30]) );
  MUX41_137 MUXES_31 ( .A(A[31]), .B(B[31]), .C(C[31]), .D(D[31]), .S({n6, n3}), .Y(Y[31]) );
  BUF_X1 U1 ( .A(SEL[1]), .Z(n4) );
  BUF_X1 U2 ( .A(SEL[1]), .Z(n5) );
  BUF_X1 U3 ( .A(SEL[1]), .Z(n6) );
  BUF_X1 U4 ( .A(SEL[0]), .Z(n1) );
  BUF_X1 U5 ( .A(SEL[0]), .Z(n2) );
  BUF_X1 U6 ( .A(SEL[0]), .Z(n3) );
endmodule


module MUX41_136 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  NOR2_X1 U1 ( .A1(n1), .A2(n8), .ZN(n9) );
  NOR2_X1 U2 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  OAI211_X1 U3 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n13), .ZN(n11) );
  AOI22_X1 U5 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_135 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  OAI211_X2 U1 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  NOR2_X1 U2 ( .A1(n1), .A2(n8), .ZN(n9) );
  NOR2_X1 U3 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  NAND2_X1 U4 ( .A1(B), .A2(n13), .ZN(n11) );
  AOI22_X1 U5 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_134 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  NOR2_X1 U1 ( .A1(n1), .A2(n8), .ZN(n9) );
  NOR2_X1 U2 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  OAI211_X1 U3 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n13), .ZN(n11) );
  AOI22_X1 U5 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_133 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  OAI211_X1 U1 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NOR2_X1 U2 ( .A1(n1), .A2(n8), .ZN(n9) );
  NOR2_X1 U3 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  NAND2_X1 U4 ( .A1(B), .A2(n13), .ZN(n11) );
  AOI22_X1 U5 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_132 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  NOR2_X1 U1 ( .A1(n1), .A2(n8), .ZN(n9) );
  NOR2_X1 U2 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  OAI211_X1 U3 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n13), .ZN(n11) );
  AOI22_X1 U5 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_131 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  NOR2_X1 U1 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  NOR2_X1 U2 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  OAI211_X1 U3 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U5 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_130 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  NOR2_X1 U1 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  NOR2_X1 U2 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  OAI211_X1 U3 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U5 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_129 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  NOR2_X1 U1 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  NOR2_X1 U2 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  OAI211_X1 U3 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U5 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_128 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  NOR2_X1 U1 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  NOR2_X1 U2 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  OAI211_X1 U3 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U5 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_127 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  NOR2_X1 U1 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  NOR2_X1 U2 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  OAI211_X1 U3 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U5 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_126 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  NOR2_X1 U1 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  NOR2_X1 U2 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  OAI211_X1 U3 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U5 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_125 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  NOR2_X1 U1 ( .A1(n1), .A2(n8), .ZN(n9) );
  NOR2_X1 U2 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  OAI211_X1 U3 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n13), .ZN(n11) );
  AOI22_X1 U5 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_124 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  NOR2_X1 U1 ( .A1(n1), .A2(n8), .ZN(n9) );
  NOR2_X1 U2 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  OAI211_X1 U3 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n13), .ZN(n11) );
  AOI22_X1 U5 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_123 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  NOR2_X1 U1 ( .A1(n1), .A2(n8), .ZN(n9) );
  NOR2_X1 U2 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  OAI211_X1 U3 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n13), .ZN(n11) );
  AOI22_X1 U5 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_122 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  NOR2_X1 U1 ( .A1(n1), .A2(n8), .ZN(n9) );
  NOR2_X1 U2 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  OAI211_X1 U3 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n13), .ZN(n11) );
  AOI22_X1 U5 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_121 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  NOR2_X1 U1 ( .A1(n1), .A2(n8), .ZN(n9) );
  NOR2_X1 U2 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  OAI211_X1 U3 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n13), .ZN(n11) );
  AOI22_X1 U5 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_120 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  NOR2_X1 U1 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  NOR2_X1 U2 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  OAI211_X1 U3 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U5 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_119 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  NOR2_X1 U1 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  NOR2_X1 U2 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  OAI211_X1 U3 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U5 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_118 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  NOR2_X1 U1 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  NOR2_X1 U2 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  OAI211_X1 U3 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U5 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_117 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  NOR2_X1 U1 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  NOR2_X1 U2 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  OAI211_X1 U3 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U5 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_116 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  NOR2_X1 U1 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  NOR2_X1 U2 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  OAI211_X1 U3 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U5 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_115 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  NOR2_X1 U1 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  NOR2_X1 U2 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  OAI211_X1 U3 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U5 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_114 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  NOR2_X1 U1 ( .A1(n1), .A2(n8), .ZN(n9) );
  NOR2_X1 U2 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  OAI211_X1 U3 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n13), .ZN(n11) );
  AOI22_X1 U5 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_113 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  NOR2_X1 U1 ( .A1(n1), .A2(n8), .ZN(n9) );
  NOR2_X1 U2 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  OAI211_X1 U3 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n13), .ZN(n11) );
  AOI22_X1 U5 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_112 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  NOR2_X1 U1 ( .A1(n1), .A2(n8), .ZN(n9) );
  NOR2_X1 U2 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  OAI211_X1 U3 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n13), .ZN(n11) );
  AOI22_X1 U5 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_111 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  NOR2_X1 U1 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  NOR2_X1 U2 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  OAI211_X1 U3 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U5 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_110 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  NOR2_X1 U1 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  NOR2_X1 U2 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  OAI211_X1 U3 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U5 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_109 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  NOR2_X1 U1 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  NOR2_X1 U2 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  OAI211_X1 U3 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U5 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_108 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  NOR2_X1 U1 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  NOR2_X1 U2 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  OAI211_X1 U3 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U5 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_107 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  NOR2_X1 U1 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  NOR2_X1 U2 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  OAI211_X1 U3 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U5 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_106 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  NOR2_X1 U1 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  NOR2_X1 U2 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  OAI211_X1 U3 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U5 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_105 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  NOR2_X1 U1 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  NOR2_X1 U2 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  OAI211_X1 U3 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U5 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_GENERIC_NBIT32_2 ( A, B, C, D, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [31:0] D;
  input [1:0] SEL;
  output [31:0] Y;
  wire   n1, n2, n3, n4, n5, n6;

  MUX41_136 MUXES_0 ( .A(A[0]), .B(B[0]), .C(C[0]), .D(D[0]), .S({n4, n1}), 
        .Y(Y[0]) );
  MUX41_135 MUXES_1 ( .A(A[1]), .B(B[1]), .C(C[1]), .D(D[1]), .S({n4, n1}), 
        .Y(Y[1]) );
  MUX41_134 MUXES_2 ( .A(A[2]), .B(B[2]), .C(C[2]), .D(D[2]), .S({n4, n1}), 
        .Y(Y[2]) );
  MUX41_133 MUXES_3 ( .A(A[3]), .B(B[3]), .C(C[3]), .D(D[3]), .S({n4, n1}), 
        .Y(Y[3]) );
  MUX41_132 MUXES_4 ( .A(A[4]), .B(B[4]), .C(C[4]), .D(D[4]), .S({n4, n1}), 
        .Y(Y[4]) );
  MUX41_131 MUXES_5 ( .A(A[5]), .B(B[5]), .C(C[5]), .D(D[5]), .S({n4, n1}), 
        .Y(Y[5]) );
  MUX41_130 MUXES_6 ( .A(A[6]), .B(B[6]), .C(C[6]), .D(D[6]), .S({n4, n1}), 
        .Y(Y[6]) );
  MUX41_129 MUXES_7 ( .A(A[7]), .B(B[7]), .C(C[7]), .D(D[7]), .S({n4, n1}), 
        .Y(Y[7]) );
  MUX41_128 MUXES_8 ( .A(A[8]), .B(B[8]), .C(C[8]), .D(D[8]), .S({n4, n1}), 
        .Y(Y[8]) );
  MUX41_127 MUXES_9 ( .A(A[9]), .B(B[9]), .C(C[9]), .D(D[9]), .S({n4, n1}), 
        .Y(Y[9]) );
  MUX41_126 MUXES_10 ( .A(A[10]), .B(B[10]), .C(C[10]), .D(D[10]), .S({n4, n1}), .Y(Y[10]) );
  MUX41_125 MUXES_11 ( .A(A[11]), .B(B[11]), .C(C[11]), .D(D[11]), .S({n4, n2}), .Y(Y[11]) );
  MUX41_124 MUXES_12 ( .A(A[12]), .B(B[12]), .C(C[12]), .D(D[12]), .S({n5, n2}), .Y(Y[12]) );
  MUX41_123 MUXES_13 ( .A(A[13]), .B(B[13]), .C(C[13]), .D(D[13]), .S({n5, n2}), .Y(Y[13]) );
  MUX41_122 MUXES_14 ( .A(A[14]), .B(B[14]), .C(C[14]), .D(D[14]), .S({n5, n2}), .Y(Y[14]) );
  MUX41_121 MUXES_15 ( .A(A[15]), .B(B[15]), .C(C[15]), .D(D[15]), .S({n5, n2}), .Y(Y[15]) );
  MUX41_120 MUXES_16 ( .A(A[16]), .B(B[16]), .C(C[16]), .D(D[16]), .S({n5, n2}), .Y(Y[16]) );
  MUX41_119 MUXES_17 ( .A(A[17]), .B(B[17]), .C(C[17]), .D(D[17]), .S({n5, n2}), .Y(Y[17]) );
  MUX41_118 MUXES_18 ( .A(A[18]), .B(B[18]), .C(C[18]), .D(D[18]), .S({n5, n2}), .Y(Y[18]) );
  MUX41_117 MUXES_19 ( .A(A[19]), .B(B[19]), .C(C[19]), .D(D[19]), .S({n5, n2}), .Y(Y[19]) );
  MUX41_116 MUXES_20 ( .A(A[20]), .B(B[20]), .C(C[20]), .D(D[20]), .S({n5, n2}), .Y(Y[20]) );
  MUX41_115 MUXES_21 ( .A(A[21]), .B(B[21]), .C(C[21]), .D(D[21]), .S({n5, n2}), .Y(Y[21]) );
  MUX41_114 MUXES_22 ( .A(A[22]), .B(B[22]), .C(C[22]), .D(D[22]), .S({n5, n3}), .Y(Y[22]) );
  MUX41_113 MUXES_23 ( .A(A[23]), .B(B[23]), .C(C[23]), .D(D[23]), .S({n5, n3}), .Y(Y[23]) );
  MUX41_112 MUXES_24 ( .A(A[24]), .B(B[24]), .C(C[24]), .D(D[24]), .S({n6, n3}), .Y(Y[24]) );
  MUX41_111 MUXES_25 ( .A(A[25]), .B(B[25]), .C(C[25]), .D(D[25]), .S({n6, n3}), .Y(Y[25]) );
  MUX41_110 MUXES_26 ( .A(A[26]), .B(B[26]), .C(C[26]), .D(D[26]), .S({n6, n3}), .Y(Y[26]) );
  MUX41_109 MUXES_27 ( .A(A[27]), .B(B[27]), .C(C[27]), .D(D[27]), .S({n6, n3}), .Y(Y[27]) );
  MUX41_108 MUXES_28 ( .A(A[28]), .B(B[28]), .C(C[28]), .D(D[28]), .S({n6, n3}), .Y(Y[28]) );
  MUX41_107 MUXES_29 ( .A(A[29]), .B(B[29]), .C(C[29]), .D(D[29]), .S({n6, n3}), .Y(Y[29]) );
  MUX41_106 MUXES_30 ( .A(A[30]), .B(B[30]), .C(C[30]), .D(D[30]), .S({n6, n3}), .Y(Y[30]) );
  MUX41_105 MUXES_31 ( .A(A[31]), .B(B[31]), .C(C[31]), .D(D[31]), .S({n6, n3}), .Y(Y[31]) );
  BUF_X1 U1 ( .A(SEL[1]), .Z(n5) );
  BUF_X1 U2 ( .A(SEL[1]), .Z(n4) );
  BUF_X1 U3 ( .A(SEL[1]), .Z(n6) );
  BUF_X1 U4 ( .A(SEL[0]), .Z(n2) );
  BUF_X1 U5 ( .A(SEL[0]), .Z(n1) );
  BUF_X1 U6 ( .A(SEL[0]), .Z(n3) );
endmodule


module MUX41_104 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  AOI22_X1 U1 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  NOR2_X1 U2 ( .A1(n1), .A2(n8), .ZN(n9) );
  OAI211_X1 U3 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n13), .ZN(n11) );
  NOR2_X1 U5 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_103 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  AOI22_X1 U1 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  NOR2_X1 U2 ( .A1(n1), .A2(n8), .ZN(n9) );
  OAI211_X1 U3 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n13), .ZN(n11) );
  NOR2_X1 U5 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_102 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  AOI22_X1 U1 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  NOR2_X1 U2 ( .A1(n1), .A2(n8), .ZN(n9) );
  OAI211_X1 U3 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n13), .ZN(n11) );
  NOR2_X1 U5 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_101 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  AOI22_X1 U1 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  NOR2_X1 U2 ( .A1(n1), .A2(n8), .ZN(n9) );
  OAI211_X1 U3 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n13), .ZN(n11) );
  NOR2_X1 U5 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_100 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  AOI22_X1 U1 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  NOR2_X1 U2 ( .A1(n1), .A2(n8), .ZN(n9) );
  OAI211_X1 U3 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n13), .ZN(n11) );
  NOR2_X1 U5 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_99 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  AOI22_X1 U1 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  NOR2_X1 U2 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  OAI211_X1 U3 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  NOR2_X1 U5 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_98 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  AOI22_X1 U1 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  NOR2_X1 U2 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  OAI211_X1 U3 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  NOR2_X1 U5 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_97 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  AOI22_X1 U1 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  NOR2_X1 U2 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  OAI211_X1 U3 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  NOR2_X1 U5 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_96 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  AOI22_X1 U1 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  NOR2_X1 U2 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  OAI211_X1 U3 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  NOR2_X1 U5 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_95 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  AOI22_X1 U1 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  NOR2_X1 U2 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  OAI211_X1 U3 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  NOR2_X1 U5 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_94 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  AOI22_X1 U1 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  NOR2_X1 U2 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  OAI211_X1 U3 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  NOR2_X1 U5 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_93 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  AOI22_X1 U1 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  NOR2_X1 U2 ( .A1(n1), .A2(n8), .ZN(n9) );
  OAI211_X1 U3 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n13), .ZN(n11) );
  NOR2_X1 U5 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_92 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  AOI22_X1 U1 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  NOR2_X1 U2 ( .A1(n1), .A2(n8), .ZN(n9) );
  OAI211_X1 U3 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n13), .ZN(n11) );
  NOR2_X1 U5 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_91 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  AOI22_X1 U1 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  NOR2_X1 U2 ( .A1(n1), .A2(n8), .ZN(n9) );
  OAI211_X1 U3 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n13), .ZN(n11) );
  NOR2_X1 U5 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_90 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  AOI22_X1 U1 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  NOR2_X1 U2 ( .A1(n1), .A2(n8), .ZN(n9) );
  OAI211_X1 U3 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n13), .ZN(n11) );
  NOR2_X1 U5 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_89 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  AOI22_X1 U1 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  NOR2_X1 U2 ( .A1(n1), .A2(n8), .ZN(n9) );
  OAI211_X1 U3 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n13), .ZN(n11) );
  NOR2_X1 U5 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_88 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  AOI22_X1 U1 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  NOR2_X1 U2 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  OAI211_X1 U3 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  NOR2_X1 U5 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_87 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  AOI22_X1 U1 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  NOR2_X1 U2 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  OAI211_X1 U3 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  NOR2_X1 U5 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_86 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  AOI22_X1 U1 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  NOR2_X1 U2 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  OAI211_X1 U3 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  NOR2_X1 U5 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_85 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  AOI22_X1 U1 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  NOR2_X1 U2 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  OAI211_X1 U3 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  NOR2_X1 U5 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_84 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  AOI22_X1 U1 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  NOR2_X1 U2 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  OAI211_X1 U3 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  NOR2_X1 U5 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_83 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  AOI22_X1 U1 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  NOR2_X1 U2 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  OAI211_X1 U3 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  NOR2_X1 U5 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_82 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  AOI22_X1 U1 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  NOR2_X1 U2 ( .A1(n1), .A2(n8), .ZN(n9) );
  OAI211_X1 U3 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n13), .ZN(n11) );
  NOR2_X1 U5 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_81 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  AOI22_X1 U1 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  NOR2_X1 U2 ( .A1(n1), .A2(n8), .ZN(n9) );
  OAI211_X1 U3 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n13), .ZN(n11) );
  NOR2_X1 U5 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_80 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  AOI22_X1 U1 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  NOR2_X1 U2 ( .A1(n1), .A2(n8), .ZN(n9) );
  OAI211_X1 U3 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n13), .ZN(n11) );
  NOR2_X1 U5 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_79 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  AOI22_X1 U1 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  NOR2_X1 U2 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  OAI211_X1 U3 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  NOR2_X1 U5 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_78 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  AOI22_X1 U1 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  NOR2_X1 U2 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  OAI211_X1 U3 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  NOR2_X1 U5 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_77 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  AOI22_X1 U1 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  NOR2_X1 U2 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  OAI211_X1 U3 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  NOR2_X1 U5 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_76 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  AOI22_X1 U1 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  NOR2_X1 U2 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  OAI211_X1 U3 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  NOR2_X1 U5 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_75 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  AOI22_X1 U1 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  NOR2_X1 U2 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  OAI211_X1 U3 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  NOR2_X1 U5 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_74 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  AOI22_X1 U1 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  NOR2_X1 U2 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  OAI211_X1 U3 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  NOR2_X1 U5 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_73 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  AOI22_X1 U1 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  NOR2_X1 U2 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  OAI211_X1 U3 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  NOR2_X1 U5 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_GENERIC_NBIT32_1 ( A, B, C, D, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [31:0] D;
  input [1:0] SEL;
  output [31:0] Y;
  wire   n1, n2, n3, n4, n5, n6;

  MUX41_104 MUXES_0 ( .A(A[0]), .B(B[0]), .C(C[0]), .D(D[0]), .S({n4, n1}), 
        .Y(Y[0]) );
  MUX41_103 MUXES_1 ( .A(A[1]), .B(B[1]), .C(C[1]), .D(D[1]), .S({n4, n1}), 
        .Y(Y[1]) );
  MUX41_102 MUXES_2 ( .A(A[2]), .B(B[2]), .C(C[2]), .D(D[2]), .S({n4, n1}), 
        .Y(Y[2]) );
  MUX41_101 MUXES_3 ( .A(A[3]), .B(B[3]), .C(C[3]), .D(D[3]), .S({n4, n1}), 
        .Y(Y[3]) );
  MUX41_100 MUXES_4 ( .A(A[4]), .B(B[4]), .C(C[4]), .D(D[4]), .S({n4, n1}), 
        .Y(Y[4]) );
  MUX41_99 MUXES_5 ( .A(A[5]), .B(B[5]), .C(C[5]), .D(D[5]), .S({n4, n1}), .Y(
        Y[5]) );
  MUX41_98 MUXES_6 ( .A(A[6]), .B(B[6]), .C(C[6]), .D(D[6]), .S({n4, n1}), .Y(
        Y[6]) );
  MUX41_97 MUXES_7 ( .A(A[7]), .B(B[7]), .C(C[7]), .D(D[7]), .S({n4, n1}), .Y(
        Y[7]) );
  MUX41_96 MUXES_8 ( .A(A[8]), .B(B[8]), .C(C[8]), .D(D[8]), .S({n4, n1}), .Y(
        Y[8]) );
  MUX41_95 MUXES_9 ( .A(A[9]), .B(B[9]), .C(C[9]), .D(D[9]), .S({n4, n1}), .Y(
        Y[9]) );
  MUX41_94 MUXES_10 ( .A(A[10]), .B(B[10]), .C(C[10]), .D(D[10]), .S({n4, n1}), 
        .Y(Y[10]) );
  MUX41_93 MUXES_11 ( .A(A[11]), .B(B[11]), .C(C[11]), .D(D[11]), .S({n4, n2}), 
        .Y(Y[11]) );
  MUX41_92 MUXES_12 ( .A(A[12]), .B(B[12]), .C(C[12]), .D(D[12]), .S({n5, n2}), 
        .Y(Y[12]) );
  MUX41_91 MUXES_13 ( .A(A[13]), .B(B[13]), .C(C[13]), .D(D[13]), .S({n5, n2}), 
        .Y(Y[13]) );
  MUX41_90 MUXES_14 ( .A(A[14]), .B(B[14]), .C(C[14]), .D(D[14]), .S({n5, n2}), 
        .Y(Y[14]) );
  MUX41_89 MUXES_15 ( .A(A[15]), .B(B[15]), .C(C[15]), .D(D[15]), .S({n5, n2}), 
        .Y(Y[15]) );
  MUX41_88 MUXES_16 ( .A(A[16]), .B(B[16]), .C(C[16]), .D(D[16]), .S({n5, n2}), 
        .Y(Y[16]) );
  MUX41_87 MUXES_17 ( .A(A[17]), .B(B[17]), .C(C[17]), .D(D[17]), .S({n5, n2}), 
        .Y(Y[17]) );
  MUX41_86 MUXES_18 ( .A(A[18]), .B(B[18]), .C(C[18]), .D(D[18]), .S({n5, n2}), 
        .Y(Y[18]) );
  MUX41_85 MUXES_19 ( .A(A[19]), .B(B[19]), .C(C[19]), .D(D[19]), .S({n5, n2}), 
        .Y(Y[19]) );
  MUX41_84 MUXES_20 ( .A(A[20]), .B(B[20]), .C(C[20]), .D(D[20]), .S({n5, n2}), 
        .Y(Y[20]) );
  MUX41_83 MUXES_21 ( .A(A[21]), .B(B[21]), .C(C[21]), .D(D[21]), .S({n5, n2}), 
        .Y(Y[21]) );
  MUX41_82 MUXES_22 ( .A(A[22]), .B(B[22]), .C(C[22]), .D(D[22]), .S({n5, n3}), 
        .Y(Y[22]) );
  MUX41_81 MUXES_23 ( .A(A[23]), .B(B[23]), .C(C[23]), .D(D[23]), .S({n5, n3}), 
        .Y(Y[23]) );
  MUX41_80 MUXES_24 ( .A(A[24]), .B(B[24]), .C(C[24]), .D(D[24]), .S({n6, n3}), 
        .Y(Y[24]) );
  MUX41_79 MUXES_25 ( .A(A[25]), .B(B[25]), .C(C[25]), .D(D[25]), .S({n6, n3}), 
        .Y(Y[25]) );
  MUX41_78 MUXES_26 ( .A(A[26]), .B(B[26]), .C(C[26]), .D(D[26]), .S({n6, n3}), 
        .Y(Y[26]) );
  MUX41_77 MUXES_27 ( .A(A[27]), .B(B[27]), .C(C[27]), .D(D[27]), .S({n6, n3}), 
        .Y(Y[27]) );
  MUX41_76 MUXES_28 ( .A(A[28]), .B(B[28]), .C(C[28]), .D(D[28]), .S({n6, n3}), 
        .Y(Y[28]) );
  MUX41_75 MUXES_29 ( .A(A[29]), .B(B[29]), .C(C[29]), .D(D[29]), .S({n6, n3}), 
        .Y(Y[29]) );
  MUX41_74 MUXES_30 ( .A(A[30]), .B(B[30]), .C(C[30]), .D(D[30]), .S({n6, n3}), 
        .Y(Y[30]) );
  MUX41_73 MUXES_31 ( .A(A[31]), .B(B[31]), .C(C[31]), .D(D[31]), .S({n6, n3}), 
        .Y(Y[31]) );
  BUF_X1 U1 ( .A(SEL[1]), .Z(n5) );
  BUF_X1 U2 ( .A(SEL[1]), .Z(n4) );
  BUF_X1 U3 ( .A(SEL[1]), .Z(n6) );
  BUF_X1 U4 ( .A(SEL[0]), .Z(n2) );
  BUF_X1 U5 ( .A(SEL[0]), .Z(n1) );
  BUF_X1 U6 ( .A(SEL[0]), .Z(n3) );
endmodule


module MUX21_466 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_465 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_464 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_463 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_462 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_GENERIC_NBIT5_0 ( A, B, SEL, Y );
  input [4:0] A;
  input [4:0] B;
  output [4:0] Y;
  input SEL;


  MUX21_466 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_465 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_464 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_463 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
  MUX21_462 MUXES_4 ( .A(A[4]), .B(B[4]), .S(SEL), .Y(Y[4]) );
endmodule


module MUX21_360 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_359 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_358 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_357 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_356 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_355 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_354 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_353 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_GENERIC_NBIT8_0 ( A, B, SEL, Y );
  input [7:0] A;
  input [7:0] B;
  output [7:0] Y;
  input SEL;


  MUX21_360 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_359 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_358 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_357 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
  MUX21_356 MUXES_4 ( .A(A[4]), .B(B[4]), .S(SEL), .Y(Y[4]) );
  MUX21_355 MUXES_5 ( .A(A[5]), .B(B[5]), .S(SEL), .Y(Y[5]) );
  MUX21_354 MUXES_6 ( .A(A[6]), .B(B[6]), .S(SEL), .Y(Y[6]) );
  MUX21_353 MUXES_7 ( .A(A[7]), .B(B[7]), .S(SEL), .Y(Y[7]) );
endmodule


module MUX21_352 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_351 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_350 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_349 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_348 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_347 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_346 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_345 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_GENERIC_NBIT8_16 ( A, B, SEL, Y );
  input [7:0] A;
  input [7:0] B;
  output [7:0] Y;
  input SEL;


  MUX21_352 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_351 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_350 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_349 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
  MUX21_348 MUXES_4 ( .A(A[4]), .B(B[4]), .S(SEL), .Y(Y[4]) );
  MUX21_347 MUXES_5 ( .A(A[5]), .B(B[5]), .S(SEL), .Y(Y[5]) );
  MUX21_346 MUXES_6 ( .A(A[6]), .B(B[6]), .S(SEL), .Y(Y[6]) );
  MUX21_345 MUXES_7 ( .A(A[7]), .B(B[7]), .S(SEL), .Y(Y[7]) );
endmodule


module MUX21_344 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_343 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_342 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_341 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_340 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_339 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_338 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_337 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_GENERIC_NBIT8_15 ( A, B, SEL, Y );
  input [7:0] A;
  input [7:0] B;
  output [7:0] Y;
  input SEL;


  MUX21_344 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_343 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_342 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_341 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
  MUX21_340 MUXES_4 ( .A(A[4]), .B(B[4]), .S(SEL), .Y(Y[4]) );
  MUX21_339 MUXES_5 ( .A(A[5]), .B(B[5]), .S(SEL), .Y(Y[5]) );
  MUX21_338 MUXES_6 ( .A(A[6]), .B(B[6]), .S(SEL), .Y(Y[6]) );
  MUX21_337 MUXES_7 ( .A(A[7]), .B(B[7]), .S(SEL), .Y(Y[7]) );
endmodule


module MUX21_336 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_335 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_334 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_333 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_332 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_331 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_330 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_329 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_GENERIC_NBIT8_14 ( A, B, SEL, Y );
  input [7:0] A;
  input [7:0] B;
  output [7:0] Y;
  input SEL;


  MUX21_336 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_335 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_334 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_333 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
  MUX21_332 MUXES_4 ( .A(A[4]), .B(B[4]), .S(SEL), .Y(Y[4]) );
  MUX21_331 MUXES_5 ( .A(A[5]), .B(B[5]), .S(SEL), .Y(Y[5]) );
  MUX21_330 MUXES_6 ( .A(A[6]), .B(B[6]), .S(SEL), .Y(Y[6]) );
  MUX21_329 MUXES_7 ( .A(A[7]), .B(B[7]), .S(SEL), .Y(Y[7]) );
endmodule


module MUX21_328 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_327 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_326 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_325 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_324 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_323 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_322 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_321 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_GENERIC_NBIT8_13 ( A, B, SEL, Y );
  input [7:0] A;
  input [7:0] B;
  output [7:0] Y;
  input SEL;


  MUX21_328 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_327 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_326 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_325 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
  MUX21_324 MUXES_4 ( .A(A[4]), .B(B[4]), .S(SEL), .Y(Y[4]) );
  MUX21_323 MUXES_5 ( .A(A[5]), .B(B[5]), .S(SEL), .Y(Y[5]) );
  MUX21_322 MUXES_6 ( .A(A[6]), .B(B[6]), .S(SEL), .Y(Y[6]) );
  MUX21_321 MUXES_7 ( .A(A[7]), .B(B[7]), .S(SEL), .Y(Y[7]) );
endmodule


module MUX41_32 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  NOR2_X1 U1 ( .A1(n1), .A2(n8), .ZN(n9) );
  OAI211_X1 U2 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND2_X1 U3 ( .A1(B), .A2(n13), .ZN(n11) );
  AOI22_X1 U4 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  NOR2_X1 U5 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_31 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  NOR2_X1 U1 ( .A1(n1), .A2(n8), .ZN(n9) );
  OAI211_X1 U2 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND2_X1 U3 ( .A1(B), .A2(n13), .ZN(n11) );
  AOI22_X1 U4 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  NOR2_X1 U5 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_30 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  NOR2_X1 U1 ( .A1(n1), .A2(n8), .ZN(n9) );
  OAI211_X1 U2 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND2_X1 U3 ( .A1(B), .A2(n13), .ZN(n11) );
  AOI22_X1 U4 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  NOR2_X1 U5 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_29 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  NOR2_X1 U1 ( .A1(n1), .A2(n8), .ZN(n9) );
  OAI211_X1 U2 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND2_X1 U3 ( .A1(B), .A2(n13), .ZN(n11) );
  AOI22_X1 U4 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  NOR2_X1 U5 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_28 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  NOR2_X1 U1 ( .A1(n1), .A2(n8), .ZN(n9) );
  OAI211_X1 U2 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND2_X1 U3 ( .A1(B), .A2(n13), .ZN(n11) );
  AOI22_X1 U4 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  NOR2_X1 U5 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_27 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  NOR2_X1 U1 ( .A1(n1), .A2(n8), .ZN(n9) );
  OAI211_X1 U2 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND2_X1 U3 ( .A1(B), .A2(n13), .ZN(n11) );
  AOI22_X1 U4 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  NOR2_X1 U5 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_26 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  NOR2_X1 U1 ( .A1(n1), .A2(n8), .ZN(n9) );
  OAI211_X1 U2 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  AOI22_X1 U3 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  NAND2_X1 U4 ( .A1(B), .A2(n13), .ZN(n11) );
  NOR2_X1 U5 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_25 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  NOR2_X1 U1 ( .A1(n1), .A2(n8), .ZN(n9) );
  OAI211_X1 U2 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND2_X1 U3 ( .A1(B), .A2(n13), .ZN(n11) );
  AOI22_X1 U4 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  NOR2_X1 U5 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_GENERIC_NBIT8_0 ( A, B, C, D, SEL, Y );
  input [7:0] A;
  input [7:0] B;
  input [7:0] C;
  input [7:0] D;
  input [1:0] SEL;
  output [7:0] Y;


  MUX41_32 MUXES_0 ( .A(A[0]), .B(B[0]), .C(C[0]), .D(D[0]), .S(SEL), .Y(Y[0])
         );
  MUX41_31 MUXES_1 ( .A(A[1]), .B(B[1]), .C(C[1]), .D(D[1]), .S(SEL), .Y(Y[1])
         );
  MUX41_30 MUXES_2 ( .A(A[2]), .B(B[2]), .C(C[2]), .D(D[2]), .S(SEL), .Y(Y[2])
         );
  MUX41_29 MUXES_3 ( .A(A[3]), .B(B[3]), .C(C[3]), .D(D[3]), .S(SEL), .Y(Y[3])
         );
  MUX41_28 MUXES_4 ( .A(A[4]), .B(B[4]), .C(C[4]), .D(D[4]), .S(SEL), .Y(Y[4])
         );
  MUX41_27 MUXES_5 ( .A(A[5]), .B(B[5]), .C(C[5]), .D(D[5]), .S(SEL), .Y(Y[5])
         );
  MUX41_26 MUXES_6 ( .A(A[6]), .B(B[6]), .C(C[6]), .D(D[6]), .S(SEL), .Y(Y[6])
         );
  MUX41_25 MUXES_7 ( .A(A[7]), .B(B[7]), .C(C[7]), .D(D[7]), .S(SEL), .Y(Y[7])
         );
endmodule


module MUX21_320 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_319 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_318 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_317 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_316 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_315 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_314 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_313 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_GENERIC_NBIT8_12 ( A, B, SEL, Y );
  input [7:0] A;
  input [7:0] B;
  output [7:0] Y;
  input SEL;


  MUX21_320 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_319 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_318 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_317 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
  MUX21_316 MUXES_4 ( .A(A[4]), .B(B[4]), .S(SEL), .Y(Y[4]) );
  MUX21_315 MUXES_5 ( .A(A[5]), .B(B[5]), .S(SEL), .Y(Y[5]) );
  MUX21_314 MUXES_6 ( .A(A[6]), .B(B[6]), .S(SEL), .Y(Y[6]) );
  MUX21_313 MUXES_7 ( .A(A[7]), .B(B[7]), .S(SEL), .Y(Y[7]) );
endmodule


module MUX21_312 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_311 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_310 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_309 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_308 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_307 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_306 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_305 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_GENERIC_NBIT8_11 ( A, B, SEL, Y );
  input [7:0] A;
  input [7:0] B;
  output [7:0] Y;
  input SEL;


  MUX21_312 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_311 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_310 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_309 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
  MUX21_308 MUXES_4 ( .A(A[4]), .B(B[4]), .S(SEL), .Y(Y[4]) );
  MUX21_307 MUXES_5 ( .A(A[5]), .B(B[5]), .S(SEL), .Y(Y[5]) );
  MUX21_306 MUXES_6 ( .A(A[6]), .B(B[6]), .S(SEL), .Y(Y[6]) );
  MUX21_305 MUXES_7 ( .A(A[7]), .B(B[7]), .S(SEL), .Y(Y[7]) );
endmodule


module MUX21_304 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_303 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_302 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_301 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_300 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_299 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_298 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_297 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_GENERIC_NBIT8_10 ( A, B, SEL, Y );
  input [7:0] A;
  input [7:0] B;
  output [7:0] Y;
  input SEL;


  MUX21_304 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_303 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_302 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_301 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
  MUX21_300 MUXES_4 ( .A(A[4]), .B(B[4]), .S(SEL), .Y(Y[4]) );
  MUX21_299 MUXES_5 ( .A(A[5]), .B(B[5]), .S(SEL), .Y(Y[5]) );
  MUX21_298 MUXES_6 ( .A(A[6]), .B(B[6]), .S(SEL), .Y(Y[6]) );
  MUX21_297 MUXES_7 ( .A(A[7]), .B(B[7]), .S(SEL), .Y(Y[7]) );
endmodule


module MUX21_296 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_295 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_294 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_293 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_292 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_291 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_290 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_289 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_GENERIC_NBIT8_9 ( A, B, SEL, Y );
  input [7:0] A;
  input [7:0] B;
  output [7:0] Y;
  input SEL;


  MUX21_296 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_295 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_294 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_293 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
  MUX21_292 MUXES_4 ( .A(A[4]), .B(B[4]), .S(SEL), .Y(Y[4]) );
  MUX21_291 MUXES_5 ( .A(A[5]), .B(B[5]), .S(SEL), .Y(Y[5]) );
  MUX21_290 MUXES_6 ( .A(A[6]), .B(B[6]), .S(SEL), .Y(Y[6]) );
  MUX21_289 MUXES_7 ( .A(A[7]), .B(B[7]), .S(SEL), .Y(Y[7]) );
endmodule


module MUX41_24 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  NOR2_X1 U1 ( .A1(n1), .A2(n8), .ZN(n9) );
  OAI211_X1 U2 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND2_X1 U3 ( .A1(B), .A2(n13), .ZN(n11) );
  AOI22_X1 U4 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  NOR2_X1 U5 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_23 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  NOR2_X1 U1 ( .A1(n1), .A2(n8), .ZN(n9) );
  OAI211_X1 U2 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND2_X1 U3 ( .A1(B), .A2(n13), .ZN(n11) );
  AOI22_X1 U4 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  NOR2_X1 U5 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_22 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  NOR2_X1 U1 ( .A1(n1), .A2(n8), .ZN(n9) );
  OAI211_X1 U2 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND2_X1 U3 ( .A1(B), .A2(n13), .ZN(n11) );
  AOI22_X1 U4 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  NOR2_X1 U5 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_21 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  NOR2_X1 U1 ( .A1(n1), .A2(n8), .ZN(n9) );
  OAI211_X1 U2 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND2_X1 U3 ( .A1(B), .A2(n13), .ZN(n11) );
  AOI22_X1 U4 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  NOR2_X1 U5 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_20 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  NOR2_X1 U1 ( .A1(n1), .A2(n8), .ZN(n9) );
  OAI211_X1 U2 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND2_X1 U3 ( .A1(B), .A2(n13), .ZN(n11) );
  AOI22_X1 U4 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  NOR2_X1 U5 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_19 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  NOR2_X1 U1 ( .A1(n1), .A2(n8), .ZN(n9) );
  OAI211_X1 U2 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND2_X1 U3 ( .A1(B), .A2(n13), .ZN(n11) );
  AOI22_X1 U4 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  NOR2_X1 U5 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_18 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  NOR2_X1 U1 ( .A1(n1), .A2(n8), .ZN(n9) );
  OAI211_X1 U2 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND2_X1 U3 ( .A1(B), .A2(n13), .ZN(n11) );
  AOI22_X1 U4 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  NOR2_X1 U5 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_17 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  NOR2_X1 U1 ( .A1(n1), .A2(n8), .ZN(n9) );
  OAI211_X1 U2 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND2_X1 U3 ( .A1(B), .A2(n13), .ZN(n11) );
  AOI22_X1 U4 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  NOR2_X1 U5 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_GENERIC_NBIT8_3 ( A, B, C, D, SEL, Y );
  input [7:0] A;
  input [7:0] B;
  input [7:0] C;
  input [7:0] D;
  input [1:0] SEL;
  output [7:0] Y;


  MUX41_24 MUXES_0 ( .A(A[0]), .B(B[0]), .C(C[0]), .D(D[0]), .S(SEL), .Y(Y[0])
         );
  MUX41_23 MUXES_1 ( .A(A[1]), .B(B[1]), .C(C[1]), .D(D[1]), .S(SEL), .Y(Y[1])
         );
  MUX41_22 MUXES_2 ( .A(A[2]), .B(B[2]), .C(C[2]), .D(D[2]), .S(SEL), .Y(Y[2])
         );
  MUX41_21 MUXES_3 ( .A(A[3]), .B(B[3]), .C(C[3]), .D(D[3]), .S(SEL), .Y(Y[3])
         );
  MUX41_20 MUXES_4 ( .A(A[4]), .B(B[4]), .C(C[4]), .D(D[4]), .S(SEL), .Y(Y[4])
         );
  MUX41_19 MUXES_5 ( .A(A[5]), .B(B[5]), .C(C[5]), .D(D[5]), .S(SEL), .Y(Y[5])
         );
  MUX41_18 MUXES_6 ( .A(A[6]), .B(B[6]), .C(C[6]), .D(D[6]), .S(SEL), .Y(Y[6])
         );
  MUX41_17 MUXES_7 ( .A(A[7]), .B(B[7]), .C(C[7]), .D(D[7]), .S(SEL), .Y(Y[7])
         );
endmodule


module MUX21_288 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_287 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_286 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_285 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_284 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_283 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_282 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_281 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_GENERIC_NBIT8_8 ( A, B, SEL, Y );
  input [7:0] A;
  input [7:0] B;
  output [7:0] Y;
  input SEL;


  MUX21_288 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_287 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_286 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_285 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
  MUX21_284 MUXES_4 ( .A(A[4]), .B(B[4]), .S(SEL), .Y(Y[4]) );
  MUX21_283 MUXES_5 ( .A(A[5]), .B(B[5]), .S(SEL), .Y(Y[5]) );
  MUX21_282 MUXES_6 ( .A(A[6]), .B(B[6]), .S(SEL), .Y(Y[6]) );
  MUX21_281 MUXES_7 ( .A(A[7]), .B(B[7]), .S(SEL), .Y(Y[7]) );
endmodule


module MUX21_280 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_279 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_278 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_277 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_276 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_275 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_274 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_273 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_GENERIC_NBIT8_7 ( A, B, SEL, Y );
  input [7:0] A;
  input [7:0] B;
  output [7:0] Y;
  input SEL;


  MUX21_280 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_279 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_278 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_277 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
  MUX21_276 MUXES_4 ( .A(A[4]), .B(B[4]), .S(SEL), .Y(Y[4]) );
  MUX21_275 MUXES_5 ( .A(A[5]), .B(B[5]), .S(SEL), .Y(Y[5]) );
  MUX21_274 MUXES_6 ( .A(A[6]), .B(B[6]), .S(SEL), .Y(Y[6]) );
  MUX21_273 MUXES_7 ( .A(A[7]), .B(B[7]), .S(SEL), .Y(Y[7]) );
endmodule


module MUX21_272 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_271 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_270 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_269 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_268 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_267 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_266 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_265 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_GENERIC_NBIT8_6 ( A, B, SEL, Y );
  input [7:0] A;
  input [7:0] B;
  output [7:0] Y;
  input SEL;


  MUX21_272 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_271 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_270 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_269 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
  MUX21_268 MUXES_4 ( .A(A[4]), .B(B[4]), .S(SEL), .Y(Y[4]) );
  MUX21_267 MUXES_5 ( .A(A[5]), .B(B[5]), .S(SEL), .Y(Y[5]) );
  MUX21_266 MUXES_6 ( .A(A[6]), .B(B[6]), .S(SEL), .Y(Y[6]) );
  MUX21_265 MUXES_7 ( .A(A[7]), .B(B[7]), .S(SEL), .Y(Y[7]) );
endmodule


module MUX21_264 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_263 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_262 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_261 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_260 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_259 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_258 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_257 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_GENERIC_NBIT8_5 ( A, B, SEL, Y );
  input [7:0] A;
  input [7:0] B;
  output [7:0] Y;
  input SEL;


  MUX21_264 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_263 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_262 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_261 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
  MUX21_260 MUXES_4 ( .A(A[4]), .B(B[4]), .S(SEL), .Y(Y[4]) );
  MUX21_259 MUXES_5 ( .A(A[5]), .B(B[5]), .S(SEL), .Y(Y[5]) );
  MUX21_258 MUXES_6 ( .A(A[6]), .B(B[6]), .S(SEL), .Y(Y[6]) );
  MUX21_257 MUXES_7 ( .A(A[7]), .B(B[7]), .S(SEL), .Y(Y[7]) );
endmodule


module MUX41_16 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  NOR2_X1 U1 ( .A1(n1), .A2(n8), .ZN(n9) );
  OAI211_X1 U2 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND2_X1 U3 ( .A1(B), .A2(n13), .ZN(n11) );
  AOI22_X1 U4 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  NOR2_X1 U5 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_15 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  NOR2_X1 U1 ( .A1(n1), .A2(n8), .ZN(n9) );
  OAI211_X1 U2 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND2_X1 U3 ( .A1(B), .A2(n13), .ZN(n11) );
  AOI22_X1 U4 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  NOR2_X1 U5 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_14 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  NOR2_X1 U1 ( .A1(n1), .A2(n8), .ZN(n9) );
  OAI211_X1 U2 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND2_X1 U3 ( .A1(B), .A2(n13), .ZN(n11) );
  AOI22_X1 U4 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  NOR2_X1 U5 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_13 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  NOR2_X1 U1 ( .A1(n1), .A2(n8), .ZN(n9) );
  OAI211_X1 U2 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND2_X1 U3 ( .A1(B), .A2(n13), .ZN(n11) );
  AOI22_X1 U4 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  NOR2_X1 U5 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_12 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  NOR2_X1 U1 ( .A1(n1), .A2(n8), .ZN(n9) );
  OAI211_X1 U2 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND2_X1 U3 ( .A1(B), .A2(n13), .ZN(n11) );
  AOI22_X1 U4 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  NOR2_X1 U5 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_11 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  NOR2_X1 U1 ( .A1(n1), .A2(n8), .ZN(n9) );
  OAI211_X1 U2 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND2_X1 U3 ( .A1(B), .A2(n13), .ZN(n11) );
  AOI22_X1 U4 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  NOR2_X1 U5 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_10 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  NOR2_X1 U1 ( .A1(n1), .A2(n8), .ZN(n9) );
  OAI211_X1 U2 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND2_X1 U3 ( .A1(B), .A2(n13), .ZN(n11) );
  AOI22_X1 U4 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  NOR2_X1 U5 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_9 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  NOR2_X1 U1 ( .A1(n1), .A2(n8), .ZN(n9) );
  OAI211_X1 U2 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND2_X1 U3 ( .A1(B), .A2(n13), .ZN(n11) );
  AOI22_X1 U4 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  NOR2_X1 U5 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_GENERIC_NBIT8_2 ( A, B, C, D, SEL, Y );
  input [7:0] A;
  input [7:0] B;
  input [7:0] C;
  input [7:0] D;
  input [1:0] SEL;
  output [7:0] Y;


  MUX41_16 MUXES_0 ( .A(A[0]), .B(B[0]), .C(C[0]), .D(D[0]), .S(SEL), .Y(Y[0])
         );
  MUX41_15 MUXES_1 ( .A(A[1]), .B(B[1]), .C(C[1]), .D(D[1]), .S(SEL), .Y(Y[1])
         );
  MUX41_14 MUXES_2 ( .A(A[2]), .B(B[2]), .C(C[2]), .D(D[2]), .S(SEL), .Y(Y[2])
         );
  MUX41_13 MUXES_3 ( .A(A[3]), .B(B[3]), .C(C[3]), .D(D[3]), .S(SEL), .Y(Y[3])
         );
  MUX41_12 MUXES_4 ( .A(A[4]), .B(B[4]), .C(C[4]), .D(D[4]), .S(SEL), .Y(Y[4])
         );
  MUX41_11 MUXES_5 ( .A(A[5]), .B(B[5]), .C(C[5]), .D(D[5]), .S(SEL), .Y(Y[5])
         );
  MUX41_10 MUXES_6 ( .A(A[6]), .B(B[6]), .C(C[6]), .D(D[6]), .S(SEL), .Y(Y[6])
         );
  MUX41_9 MUXES_7 ( .A(A[7]), .B(B[7]), .C(C[7]), .D(D[7]), .S(SEL), .Y(Y[7])
         );
endmodule


module MUX21_256 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_255 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_254 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_253 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_252 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_251 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_250 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_249 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_GENERIC_NBIT8_4 ( A, B, SEL, Y );
  input [7:0] A;
  input [7:0] B;
  output [7:0] Y;
  input SEL;


  MUX21_256 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_255 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_254 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_253 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
  MUX21_252 MUXES_4 ( .A(A[4]), .B(B[4]), .S(SEL), .Y(Y[4]) );
  MUX21_251 MUXES_5 ( .A(A[5]), .B(B[5]), .S(SEL), .Y(Y[5]) );
  MUX21_250 MUXES_6 ( .A(A[6]), .B(B[6]), .S(SEL), .Y(Y[6]) );
  MUX21_249 MUXES_7 ( .A(A[7]), .B(B[7]), .S(SEL), .Y(Y[7]) );
endmodule


module MUX21_248 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_247 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_246 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_245 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_244 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_243 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_242 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_241 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_GENERIC_NBIT8_3 ( A, B, SEL, Y );
  input [7:0] A;
  input [7:0] B;
  output [7:0] Y;
  input SEL;


  MUX21_248 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_247 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_246 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_245 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
  MUX21_244 MUXES_4 ( .A(A[4]), .B(B[4]), .S(SEL), .Y(Y[4]) );
  MUX21_243 MUXES_5 ( .A(A[5]), .B(B[5]), .S(SEL), .Y(Y[5]) );
  MUX21_242 MUXES_6 ( .A(A[6]), .B(B[6]), .S(SEL), .Y(Y[6]) );
  MUX21_241 MUXES_7 ( .A(A[7]), .B(B[7]), .S(SEL), .Y(Y[7]) );
endmodule


module MUX21_240 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_239 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_238 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_237 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_236 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_235 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_234 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_233 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_GENERIC_NBIT8_2 ( A, B, SEL, Y );
  input [7:0] A;
  input [7:0] B;
  output [7:0] Y;
  input SEL;


  MUX21_240 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_239 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_238 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_237 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
  MUX21_236 MUXES_4 ( .A(A[4]), .B(B[4]), .S(SEL), .Y(Y[4]) );
  MUX21_235 MUXES_5 ( .A(A[5]), .B(B[5]), .S(SEL), .Y(Y[5]) );
  MUX21_234 MUXES_6 ( .A(A[6]), .B(B[6]), .S(SEL), .Y(Y[6]) );
  MUX21_233 MUXES_7 ( .A(A[7]), .B(B[7]), .S(SEL), .Y(Y[7]) );
endmodule


module MUX21_232 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_231 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_230 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_229 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_228 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_227 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_226 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_225 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_GENERIC_NBIT8_1 ( A, B, SEL, Y );
  input [7:0] A;
  input [7:0] B;
  output [7:0] Y;
  input SEL;


  MUX21_232 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_231 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_230 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_229 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
  MUX21_228 MUXES_4 ( .A(A[4]), .B(B[4]), .S(SEL), .Y(Y[4]) );
  MUX21_227 MUXES_5 ( .A(A[5]), .B(B[5]), .S(SEL), .Y(Y[5]) );
  MUX21_226 MUXES_6 ( .A(A[6]), .B(B[6]), .S(SEL), .Y(Y[6]) );
  MUX21_225 MUXES_7 ( .A(A[7]), .B(B[7]), .S(SEL), .Y(Y[7]) );
endmodule


module MUX41_8 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  NOR2_X1 U1 ( .A1(n1), .A2(n8), .ZN(n9) );
  OAI211_X1 U2 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND2_X1 U3 ( .A1(B), .A2(n13), .ZN(n11) );
  AOI22_X1 U4 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  NOR2_X1 U5 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_7 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  NOR2_X1 U1 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  OAI211_X1 U2 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U3 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U4 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  NOR2_X1 U5 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_6 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  NOR2_X1 U1 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  OAI211_X1 U2 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U3 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U4 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  NOR2_X1 U5 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_5 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  NOR2_X1 U1 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  OAI211_X1 U2 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U3 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U4 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  NOR2_X1 U5 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_4 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  NOR2_X1 U1 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  OAI211_X1 U2 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U3 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U4 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  NOR2_X1 U5 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_3 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  NOR2_X1 U1 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  OAI211_X1 U2 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U3 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U4 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  NOR2_X1 U5 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_2 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  OAI211_X1 U1 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  AOI22_X1 U2 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  NOR2_X1 U3 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  NOR2_X1 U5 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_1 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  AOI22_X1 U1 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  NOR2_X1 U2 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  OAI211_X1 U3 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  NOR2_X1 U5 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_GENERIC_NBIT8_1 ( A, B, C, D, SEL, Y );
  input [7:0] A;
  input [7:0] B;
  input [7:0] C;
  input [7:0] D;
  input [1:0] SEL;
  output [7:0] Y;


  MUX41_8 MUXES_0 ( .A(A[0]), .B(B[0]), .C(C[0]), .D(D[0]), .S(SEL), .Y(Y[0])
         );
  MUX41_7 MUXES_1 ( .A(A[1]), .B(B[1]), .C(C[1]), .D(D[1]), .S(SEL), .Y(Y[1])
         );
  MUX41_6 MUXES_2 ( .A(A[2]), .B(B[2]), .C(C[2]), .D(D[2]), .S(SEL), .Y(Y[2])
         );
  MUX41_5 MUXES_3 ( .A(A[3]), .B(B[3]), .C(C[3]), .D(D[3]), .S(SEL), .Y(Y[3])
         );
  MUX41_4 MUXES_4 ( .A(A[4]), .B(B[4]), .C(C[4]), .D(D[4]), .S(SEL), .Y(Y[4])
         );
  MUX41_3 MUXES_5 ( .A(A[5]), .B(B[5]), .C(C[5]), .D(D[5]), .S(SEL), .Y(Y[5])
         );
  MUX41_2 MUXES_6 ( .A(A[6]), .B(B[6]), .C(C[6]), .D(D[6]), .S(SEL), .Y(Y[6])
         );
  MUX41_1 MUXES_7 ( .A(A[7]), .B(B[7]), .C(C[7]), .D(D[7]), .S(SEL), .Y(Y[7])
         );
endmodule


module mask_generator_NBITS32 ( R1, R2, LnR, AnL, RnS, mask0, mask8, mask16, 
        mask24 );
  input [31:0] R1;
  input [31:0] R2;
  output [39:0] mask0;
  output [39:0] mask8;
  output [39:0] mask16;
  output [39:0] mask24;
  input LnR, AnL, RnS;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9;
  wire   [7:0] shr_new_block;

  MUX21_GENERIC_NBIT8_0 MUX_shift_type ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .B({n9, n9, n9, n9, n9, n9, n9, n9}), .SEL(AnL), 
        .Y(shr_new_block) );
  MUX21_GENERIC_NBIT8_16 MUX_mask0_LSB_0_0 ( .A(R1[7:0]), .B({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .SEL(n3), .Y(mask0[7:0]) );
  MUX21_GENERIC_NBIT8_15 MUX_mask0_0_1 ( .A(R1[15:8]), .B(R1[7:0]), .SEL(n8), 
        .Y(mask0[15:8]) );
  MUX21_GENERIC_NBIT8_14 MUX_mask0_0_2 ( .A(R1[23:16]), .B(R1[15:8]), .SEL(n8), 
        .Y(mask0[23:16]) );
  MUX21_GENERIC_NBIT8_13 MUX_mask0_0_3 ( .A({n9, R1[30:24]}), .B(R1[23:16]), 
        .SEL(n7), .Y(mask0[31:24]) );
  MUX41_GENERIC_NBIT8_0 MUX_mask_MSB_0_4 ( .A(shr_new_block), .B(R1[7:0]), .C(
        {n9, R1[30:24]}), .D({n9, R1[30:24]}), .SEL({n3, n1}), .Y(mask0[39:32]) );
  MUX21_GENERIC_NBIT8_12 MUX_mask_LSB_1_0 ( .A(mask0[15:8]), .B({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .SEL(n7), .Y(mask8[7:0]) );
  MUX21_GENERIC_NBIT8_11 MUX_mask_1_1 ( .A(mask0[23:16]), .B(mask0[7:0]), 
        .SEL(n7), .Y(mask8[15:8]) );
  MUX21_GENERIC_NBIT8_10 MUX_mask_1_2 ( .A(mask0[31:24]), .B(mask0[15:8]), 
        .SEL(n6), .Y(mask8[23:16]) );
  MUX21_GENERIC_NBIT8_9 MUX_mask_1_3 ( .A(mask0[39:32]), .B(mask0[23:16]), 
        .SEL(n6), .Y(mask8[31:24]) );
  MUX41_GENERIC_NBIT8_3 MUX_mask_MSB_1_4 ( .A(shr_new_block), .B(mask0[15:8]), 
        .C(mask0[31:24]), .D(mask0[31:24]), .SEL({n2, n1}), .Y(mask8[39:32])
         );
  MUX21_GENERIC_NBIT8_8 MUX_mask_LSB_2_0 ( .A(mask8[15:8]), .B({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .SEL(n6), .Y(mask16[7:0]) );
  MUX21_GENERIC_NBIT8_7 MUX_mask_2_1 ( .A(mask8[23:16]), .B(mask8[7:0]), .SEL(
        n5), .Y(mask16[15:8]) );
  MUX21_GENERIC_NBIT8_6 MUX_mask_2_2 ( .A(mask8[31:24]), .B(mask8[15:8]), 
        .SEL(n5), .Y(mask16[23:16]) );
  MUX21_GENERIC_NBIT8_5 MUX_mask_2_3 ( .A(mask8[39:32]), .B(mask8[23:16]), 
        .SEL(n4), .Y(mask16[31:24]) );
  MUX41_GENERIC_NBIT8_2 MUX_mask_MSB_2_4 ( .A(shr_new_block), .B(mask8[15:8]), 
        .C(mask8[31:24]), .D(mask8[31:24]), .SEL({n2, n1}), .Y(mask16[39:32])
         );
  MUX21_GENERIC_NBIT8_4 MUX_mask_LSB_3_0 ( .A(mask16[15:8]), .B({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .SEL(n5), .Y(mask24[7:0]) );
  MUX21_GENERIC_NBIT8_3 MUX_mask_3_1 ( .A(mask16[23:16]), .B(mask16[7:0]), 
        .SEL(n4), .Y(mask24[15:8]) );
  MUX21_GENERIC_NBIT8_2 MUX_mask_3_2 ( .A(mask16[31:24]), .B(mask16[15:8]), 
        .SEL(n4), .Y(mask24[23:16]) );
  MUX21_GENERIC_NBIT8_1 MUX_mask_3_3 ( .A(mask16[39:32]), .B(mask16[23:16]), 
        .SEL(n3), .Y(mask24[31:24]) );
  MUX41_GENERIC_NBIT8_1 MUX_mask_MSB_3_4 ( .A(shr_new_block), .B(mask16[15:8]), 
        .C(mask16[31:24]), .D(mask16[31:24]), .SEL({n2, n1}), .Y(mask24[39:32]) );
  BUF_X2 U2 ( .A(LnR), .Z(n2) );
  BUF_X2 U3 ( .A(LnR), .Z(n4) );
  BUF_X2 U4 ( .A(LnR), .Z(n6) );
  BUF_X2 U5 ( .A(LnR), .Z(n5) );
  BUF_X2 U6 ( .A(LnR), .Z(n7) );
  BUF_X2 U7 ( .A(LnR), .Z(n3) );
  BUF_X1 U8 ( .A(R1[31]), .Z(n9) );
  BUF_X2 U9 ( .A(LnR), .Z(n8) );
  BUF_X2 U10 ( .A(RnS), .Z(n1) );
endmodule


module MUX41_72 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  NOR2_X1 U1 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  AOI22_X1 U2 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  NOR2_X1 U3 ( .A1(n1), .A2(n8), .ZN(n9) );
  OAI211_X1 U4 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND2_X1 U5 ( .A1(B), .A2(n13), .ZN(n11) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_71 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  NOR2_X1 U1 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  AOI22_X1 U2 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  NOR2_X1 U3 ( .A1(n1), .A2(n8), .ZN(n9) );
  OAI211_X1 U4 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND2_X1 U5 ( .A1(B), .A2(n13), .ZN(n11) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_70 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  NOR2_X1 U1 ( .A1(n1), .A2(n8), .ZN(n9) );
  NOR2_X1 U2 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  OAI211_X1 U3 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n13), .ZN(n11) );
  AOI22_X1 U5 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_69 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  NOR2_X1 U1 ( .A1(n1), .A2(n8), .ZN(n9) );
  NOR2_X1 U2 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  OAI211_X1 U3 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n13), .ZN(n11) );
  AOI22_X1 U5 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_68 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  NOR2_X1 U1 ( .A1(n1), .A2(n8), .ZN(n9) );
  NOR2_X1 U2 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  OAI211_X1 U3 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n13), .ZN(n11) );
  AOI22_X1 U5 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_67 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  NOR2_X1 U1 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  NOR2_X1 U2 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  OAI211_X1 U3 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U5 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_66 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  NOR2_X1 U1 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  NOR2_X1 U2 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  OAI211_X1 U3 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U5 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_65 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  NOR2_X1 U1 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  NOR2_X1 U2 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  OAI211_X1 U3 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U5 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_64 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  NOR2_X1 U1 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  NOR2_X1 U2 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  OAI211_X1 U3 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U5 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_63 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  NOR2_X1 U1 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  NOR2_X1 U2 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  OAI211_X1 U3 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U5 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_62 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  NOR2_X1 U1 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  NOR2_X1 U2 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  OAI211_X1 U3 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U5 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_61 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  NOR2_X1 U1 ( .A1(n1), .A2(n8), .ZN(n9) );
  NOR2_X1 U2 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  OAI211_X1 U3 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n13), .ZN(n11) );
  AOI22_X1 U5 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_60 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  NOR2_X1 U1 ( .A1(n1), .A2(n8), .ZN(n9) );
  NOR2_X1 U2 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  OAI211_X1 U3 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n13), .ZN(n11) );
  AOI22_X1 U5 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_59 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  NOR2_X1 U1 ( .A1(n1), .A2(n8), .ZN(n9) );
  NOR2_X1 U2 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  OAI211_X1 U3 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n13), .ZN(n11) );
  AOI22_X1 U5 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_58 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  NOR2_X1 U1 ( .A1(n1), .A2(n8), .ZN(n9) );
  NOR2_X1 U2 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  OAI211_X1 U3 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n13), .ZN(n11) );
  AOI22_X1 U5 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_57 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  NOR2_X1 U1 ( .A1(n1), .A2(n8), .ZN(n9) );
  NOR2_X1 U2 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  OAI211_X1 U3 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n13), .ZN(n11) );
  AOI22_X1 U5 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_56 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  NOR2_X1 U1 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  NOR2_X1 U2 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  OAI211_X1 U3 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U5 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_55 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  NOR2_X1 U1 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  NOR2_X1 U2 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  OAI211_X1 U3 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U5 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_54 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  NOR2_X1 U1 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  NOR2_X1 U2 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  OAI211_X1 U3 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U5 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_53 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  NOR2_X1 U1 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  NOR2_X1 U2 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  OAI211_X1 U3 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U5 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_52 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  NOR2_X1 U1 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  NOR2_X1 U2 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  OAI211_X1 U3 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U5 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_51 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  NOR2_X1 U1 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  NOR2_X1 U2 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  OAI211_X1 U3 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U5 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_50 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  NOR2_X1 U1 ( .A1(n1), .A2(n8), .ZN(n9) );
  NOR2_X1 U2 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  OAI211_X1 U3 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n13), .ZN(n11) );
  AOI22_X1 U5 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_49 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  NOR2_X1 U1 ( .A1(n1), .A2(n8), .ZN(n9) );
  NOR2_X1 U2 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  OAI211_X1 U3 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n13), .ZN(n11) );
  AOI22_X1 U5 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_48 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  NOR2_X1 U1 ( .A1(n1), .A2(n8), .ZN(n9) );
  NOR2_X1 U2 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  OAI211_X1 U3 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n13), .ZN(n11) );
  AOI22_X1 U5 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_47 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  NOR2_X1 U1 ( .A1(n1), .A2(n8), .ZN(n9) );
  NOR2_X1 U2 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  OAI211_X1 U3 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n13), .ZN(n11) );
  AOI22_X1 U5 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_46 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12, n13;

  NAND3_X1 U8 ( .A1(n2), .A2(n8), .A3(A), .ZN(n10) );
  NOR2_X1 U1 ( .A1(n1), .A2(n8), .ZN(n9) );
  NOR2_X1 U2 ( .A1(n2), .A2(S[1]), .ZN(n13) );
  OAI211_X1 U3 ( .C1(n13), .C2(n12), .A(n11), .B(n10), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n13), .ZN(n11) );
  AOI22_X1 U5 ( .A1(D), .A2(n1), .B1(n9), .B2(C), .ZN(n12) );
  INV_X1 U6 ( .A(n2), .ZN(n1) );
  INV_X1 U7 ( .A(S[0]), .ZN(n2) );
  INV_X1 U9 ( .A(S[1]), .ZN(n8) );
endmodule


module MUX41_45 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  NOR2_X1 U1 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  NOR2_X1 U2 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  OAI211_X1 U3 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U5 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_44 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  NOR2_X1 U1 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  NOR2_X1 U2 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  OAI211_X1 U3 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U5 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_43 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  NOR2_X1 U1 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  NOR2_X1 U2 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  OAI211_X1 U3 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U5 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_42 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  NOR2_X1 U1 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  NOR2_X1 U2 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  OAI211_X1 U3 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U5 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_41 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  NOR2_X1 U1 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  NOR2_X1 U2 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  OAI211_X1 U3 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U5 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_40 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  NOR2_X1 U1 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  NOR2_X1 U2 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  OAI211_X1 U3 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U5 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_39 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  NOR2_X1 U1 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  NOR2_X1 U2 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  OAI211_X1 U3 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U5 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_38 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  NOR2_X1 U1 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  NOR2_X1 U2 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  OAI211_X1 U3 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U5 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_37 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  NOR2_X1 U1 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  NOR2_X1 U2 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  OAI211_X1 U3 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U5 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_36 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  NOR2_X1 U1 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  NOR2_X1 U2 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  OAI211_X1 U3 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U5 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_35 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  NOR2_X1 U1 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  NOR2_X1 U2 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  OAI211_X1 U3 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U4 ( .A1(B), .A2(n12), .ZN(n10) );
  AOI22_X1 U5 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_34 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  NOR2_X1 U1 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  AOI22_X1 U2 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  NOR2_X1 U3 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  OAI211_X1 U4 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  NAND2_X1 U5 ( .A1(B), .A2(n12), .ZN(n10) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_33 ( A, B, C, D, S, Y );
  input [1:0] S;
  input A, B, C, D;
  output Y;
  wire   n1, n2, n8, n9, n10, n11, n12;

  NAND3_X1 U8 ( .A1(n1), .A2(n2), .A3(A), .ZN(n9) );
  NOR2_X1 U1 ( .A1(n1), .A2(S[1]), .ZN(n12) );
  OAI211_X1 U2 ( .C1(n12), .C2(n11), .A(n10), .B(n9), .ZN(Y) );
  AOI22_X1 U3 ( .A1(D), .A2(S[0]), .B1(n8), .B2(C), .ZN(n11) );
  NOR2_X1 U4 ( .A1(S[0]), .A2(n2), .ZN(n8) );
  NAND2_X1 U5 ( .A1(B), .A2(n12), .ZN(n10) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
endmodule


module MUX41_GENERIC_NBIT40 ( A, B, C, D, SEL, Y );
  input [39:0] A;
  input [39:0] B;
  input [39:0] C;
  input [39:0] D;
  input [1:0] SEL;
  output [39:0] Y;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12;

  MUX41_72 MUXES_0 ( .A(A[0]), .B(B[0]), .C(C[0]), .D(D[0]), .S({n9, n3}), .Y(
        Y[0]) );
  MUX41_71 MUXES_1 ( .A(A[1]), .B(B[1]), .C(C[1]), .D(D[1]), .S({n9, n3}), .Y(
        Y[1]) );
  MUX41_70 MUXES_2 ( .A(A[2]), .B(B[2]), .C(C[2]), .D(D[2]), .S({n9, n3}), .Y(
        Y[2]) );
  MUX41_69 MUXES_3 ( .A(A[3]), .B(B[3]), .C(C[3]), .D(D[3]), .S({n9, n3}), .Y(
        Y[3]) );
  MUX41_68 MUXES_4 ( .A(A[4]), .B(B[4]), .C(C[4]), .D(D[4]), .S({n9, n3}), .Y(
        Y[4]) );
  MUX41_67 MUXES_5 ( .A(A[5]), .B(B[5]), .C(C[5]), .D(D[5]), .S({n9, n3}), .Y(
        Y[5]) );
  MUX41_66 MUXES_6 ( .A(A[6]), .B(B[6]), .C(C[6]), .D(D[6]), .S({n9, n3}), .Y(
        Y[6]) );
  MUX41_65 MUXES_7 ( .A(A[7]), .B(B[7]), .C(C[7]), .D(D[7]), .S({n9, n3}), .Y(
        Y[7]) );
  MUX41_64 MUXES_8 ( .A(A[8]), .B(B[8]), .C(C[8]), .D(D[8]), .S({n9, n3}), .Y(
        Y[8]) );
  MUX41_63 MUXES_9 ( .A(A[9]), .B(B[9]), .C(C[9]), .D(D[9]), .S({n9, n3}), .Y(
        Y[9]) );
  MUX41_62 MUXES_10 ( .A(A[10]), .B(B[10]), .C(C[10]), .D(D[10]), .S({n9, n3}), 
        .Y(Y[10]) );
  MUX41_61 MUXES_11 ( .A(A[11]), .B(B[11]), .C(C[11]), .D(D[11]), .S({n9, n4}), 
        .Y(Y[11]) );
  MUX41_60 MUXES_12 ( .A(A[12]), .B(B[12]), .C(C[12]), .D(D[12]), .S({n10, n4}), .Y(Y[12]) );
  MUX41_59 MUXES_13 ( .A(A[13]), .B(B[13]), .C(C[13]), .D(D[13]), .S({n10, n4}), .Y(Y[13]) );
  MUX41_58 MUXES_14 ( .A(A[14]), .B(B[14]), .C(C[14]), .D(D[14]), .S({n10, n4}), .Y(Y[14]) );
  MUX41_57 MUXES_15 ( .A(A[15]), .B(B[15]), .C(C[15]), .D(D[15]), .S({n10, n4}), .Y(Y[15]) );
  MUX41_56 MUXES_16 ( .A(A[16]), .B(B[16]), .C(C[16]), .D(D[16]), .S({n10, n4}), .Y(Y[16]) );
  MUX41_55 MUXES_17 ( .A(A[17]), .B(B[17]), .C(C[17]), .D(D[17]), .S({n10, n4}), .Y(Y[17]) );
  MUX41_54 MUXES_18 ( .A(A[18]), .B(B[18]), .C(C[18]), .D(D[18]), .S({n10, n4}), .Y(Y[18]) );
  MUX41_53 MUXES_19 ( .A(A[19]), .B(B[19]), .C(C[19]), .D(D[19]), .S({n10, n4}), .Y(Y[19]) );
  MUX41_52 MUXES_20 ( .A(A[20]), .B(B[20]), .C(C[20]), .D(D[20]), .S({n10, n4}), .Y(Y[20]) );
  MUX41_51 MUXES_21 ( .A(A[21]), .B(B[21]), .C(C[21]), .D(D[21]), .S({n10, n4}), .Y(Y[21]) );
  MUX41_50 MUXES_22 ( .A(A[22]), .B(B[22]), .C(C[22]), .D(D[22]), .S({n10, n5}), .Y(Y[22]) );
  MUX41_49 MUXES_23 ( .A(A[23]), .B(B[23]), .C(C[23]), .D(D[23]), .S({n10, n5}), .Y(Y[23]) );
  MUX41_48 MUXES_24 ( .A(A[24]), .B(B[24]), .C(C[24]), .D(D[24]), .S({n11, n5}), .Y(Y[24]) );
  MUX41_47 MUXES_25 ( .A(A[25]), .B(B[25]), .C(C[25]), .D(D[25]), .S({n11, n5}), .Y(Y[25]) );
  MUX41_46 MUXES_26 ( .A(A[26]), .B(B[26]), .C(C[26]), .D(D[26]), .S({n11, n5}), .Y(Y[26]) );
  MUX41_45 MUXES_27 ( .A(A[27]), .B(B[27]), .C(C[27]), .D(D[27]), .S({n11, n5}), .Y(Y[27]) );
  MUX41_44 MUXES_28 ( .A(A[28]), .B(B[28]), .C(C[28]), .D(D[28]), .S({n11, n5}), .Y(Y[28]) );
  MUX41_43 MUXES_29 ( .A(A[29]), .B(B[29]), .C(C[29]), .D(D[29]), .S({n11, n5}), .Y(Y[29]) );
  MUX41_42 MUXES_30 ( .A(A[30]), .B(B[30]), .C(C[30]), .D(D[30]), .S({n11, n5}), .Y(Y[30]) );
  MUX41_41 MUXES_31 ( .A(A[31]), .B(B[31]), .C(C[31]), .D(D[31]), .S({n11, n5}), .Y(Y[31]) );
  MUX41_40 MUXES_32 ( .A(A[32]), .B(B[32]), .C(C[32]), .D(D[32]), .S({n11, n5}), .Y(Y[32]) );
  MUX41_39 MUXES_33 ( .A(A[33]), .B(B[33]), .C(C[33]), .D(D[33]), .S({n11, n6}), .Y(Y[33]) );
  MUX41_38 MUXES_34 ( .A(A[34]), .B(B[34]), .C(C[34]), .D(D[34]), .S({n11, n6}), .Y(Y[34]) );
  MUX41_37 MUXES_35 ( .A(A[35]), .B(B[35]), .C(C[35]), .D(D[35]), .S({n11, n6}), .Y(Y[35]) );
  MUX41_36 MUXES_36 ( .A(A[36]), .B(B[36]), .C(C[36]), .D(D[36]), .S({n12, n6}), .Y(Y[36]) );
  MUX41_35 MUXES_37 ( .A(A[37]), .B(B[37]), .C(C[37]), .D(D[37]), .S({n12, n6}), .Y(Y[37]) );
  MUX41_34 MUXES_38 ( .A(A[38]), .B(B[38]), .C(C[38]), .D(D[38]), .S({n12, n6}), .Y(Y[38]) );
  MUX41_33 MUXES_39 ( .A(A[39]), .B(B[39]), .C(C[39]), .D(D[39]), .S({n12, n6}), .Y(Y[39]) );
  BUF_X1 U1 ( .A(n7), .Z(n10) );
  BUF_X1 U2 ( .A(n7), .Z(n9) );
  BUF_X1 U3 ( .A(n8), .Z(n11) );
  BUF_X1 U4 ( .A(n8), .Z(n12) );
  BUF_X1 U5 ( .A(n1), .Z(n4) );
  BUF_X1 U6 ( .A(n1), .Z(n3) );
  BUF_X1 U7 ( .A(n2), .Z(n5) );
  BUF_X1 U8 ( .A(n2), .Z(n6) );
  BUF_X1 U9 ( .A(SEL[0]), .Z(n1) );
  BUF_X1 U10 ( .A(SEL[1]), .Z(n7) );
  BUF_X1 U11 ( .A(SEL[0]), .Z(n2) );
  BUF_X1 U12 ( .A(SEL[1]), .Z(n8) );
endmodule


module mask_shifter_NBITS40 ( R1, LnR, mask_sh0, mask_sh1, mask_sh2, mask_sh3, 
        mask_sh4, mask_sh5, mask_sh6, mask_sh7 );
  input [39:0] R1;
  output [31:0] mask_sh0;
  output [31:0] mask_sh1;
  output [31:0] mask_sh2;
  output [31:0] mask_sh3;
  output [31:0] mask_sh4;
  output [31:0] mask_sh5;
  output [31:0] mask_sh6;
  output [31:0] mask_sh7;
  input LnR;
  wire   R1_3, R1_2, R1_1, R1_0, \R1[35] , \R1[34] , \R1[33] , \R1[32] ,
         \R1[31] , \R1[30] , \R1[29] , \R1[28] , \R1[27] , \R1[26] , \R1[25] ,
         \R1[24] , \R1[23] , \R1[22] , \R1[21] , \R1[20] , \R1[19] , \R1[18] ,
         \R1[17] , \R1[16] , \R1[15] , \R1[14] , \R1[13] , \R1[12] , \R1[11] ,
         \R1[10] , \R1[9] , \R1[8] , \R1[7] , \R1[6] , \R1[5] , \R1[4] , n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n1,
         n2, n3, n4, n5, n6, n7, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95;
  assign R1_3 = R1[3];
  assign R1_2 = R1[2];
  assign R1_1 = R1[1];
  assign R1_0 = R1[0];
  assign mask_sh4[31] = \R1[35] ;
  assign \R1[35]  = R1[35];
  assign mask_sh4[30] = \R1[34] ;
  assign \R1[34]  = R1[34];
  assign mask_sh4[29] = \R1[33] ;
  assign \R1[33]  = R1[33];
  assign mask_sh4[28] = \R1[32] ;
  assign \R1[32]  = R1[32];
  assign mask_sh4[27] = \R1[31] ;
  assign \R1[31]  = R1[31];
  assign mask_sh4[26] = \R1[30] ;
  assign \R1[30]  = R1[30];
  assign mask_sh4[25] = \R1[29] ;
  assign \R1[29]  = R1[29];
  assign mask_sh4[24] = \R1[28] ;
  assign \R1[28]  = R1[28];
  assign mask_sh4[23] = \R1[27] ;
  assign \R1[27]  = R1[27];
  assign mask_sh4[22] = \R1[26] ;
  assign \R1[26]  = R1[26];
  assign mask_sh4[21] = \R1[25] ;
  assign \R1[25]  = R1[25];
  assign mask_sh4[20] = \R1[24] ;
  assign \R1[24]  = R1[24];
  assign mask_sh4[19] = \R1[23] ;
  assign \R1[23]  = R1[23];
  assign mask_sh4[18] = \R1[22] ;
  assign \R1[22]  = R1[22];
  assign mask_sh4[17] = \R1[21] ;
  assign \R1[21]  = R1[21];
  assign mask_sh4[16] = \R1[20] ;
  assign \R1[20]  = R1[20];
  assign mask_sh4[15] = \R1[19] ;
  assign \R1[19]  = R1[19];
  assign mask_sh4[14] = \R1[18] ;
  assign \R1[18]  = R1[18];
  assign mask_sh4[13] = \R1[17] ;
  assign \R1[17]  = R1[17];
  assign mask_sh4[12] = \R1[16] ;
  assign \R1[16]  = R1[16];
  assign mask_sh4[11] = \R1[15] ;
  assign \R1[15]  = R1[15];
  assign mask_sh4[10] = \R1[14] ;
  assign \R1[14]  = R1[14];
  assign mask_sh4[9] = \R1[13] ;
  assign \R1[13]  = R1[13];
  assign mask_sh4[8] = \R1[12] ;
  assign \R1[12]  = R1[12];
  assign mask_sh4[7] = \R1[11] ;
  assign \R1[11]  = R1[11];
  assign mask_sh4[6] = \R1[10] ;
  assign \R1[10]  = R1[10];
  assign mask_sh4[5] = \R1[9] ;
  assign \R1[9]  = R1[9];
  assign mask_sh4[4] = \R1[8] ;
  assign \R1[8]  = R1[8];
  assign mask_sh4[3] = \R1[7] ;
  assign \R1[7]  = R1[7];
  assign mask_sh4[2] = \R1[6] ;
  assign \R1[6]  = R1[6];
  assign mask_sh4[1] = \R1[5] ;
  assign \R1[5]  = R1[5];
  assign mask_sh4[0] = \R1[4] ;
  assign \R1[4]  = R1[4];

  NAND2_X1 U1 ( .A1(n58), .A2(n62), .ZN(mask_sh6[13]) );
  NAND2_X1 U2 ( .A1(n60), .A2(n64), .ZN(mask_sh6[12]) );
  NAND2_X1 U3 ( .A1(n61), .A2(n66), .ZN(mask_sh6[11]) );
  NAND2_X1 U4 ( .A1(n50), .A2(n53), .ZN(mask_sh6[17]) );
  NAND2_X1 U5 ( .A1(n30), .A2(n51), .ZN(mask_sh2[22]) );
  NAND2_X1 U6 ( .A1(n32), .A2(n53), .ZN(mask_sh2[21]) );
  NAND2_X1 U7 ( .A1(n52), .A2(n55), .ZN(mask_sh6[16]) );
  NAND2_X1 U8 ( .A1(n54), .A2(n57), .ZN(mask_sh6[15]) );
  NAND2_X1 U9 ( .A1(n56), .A2(n59), .ZN(mask_sh6[14]) );
  NAND2_X1 U10 ( .A1(n34), .A2(n55), .ZN(mask_sh2[20]) );
  NAND2_X1 U11 ( .A1(n37), .A2(n57), .ZN(mask_sh2[19]) );
  NAND2_X1 U12 ( .A1(n39), .A2(n59), .ZN(mask_sh2[18]) );
  NAND2_X1 U13 ( .A1(n34), .A2(n51), .ZN(mask_sh3[21]) );
  NAND2_X1 U14 ( .A1(n37), .A2(n53), .ZN(mask_sh3[20]) );
  NAND2_X1 U15 ( .A1(n39), .A2(n55), .ZN(mask_sh3[19]) );
  NAND2_X1 U16 ( .A1(n26), .A2(n47), .ZN(mask_sh2[24]) );
  NAND2_X1 U17 ( .A1(n28), .A2(n49), .ZN(mask_sh2[23]) );
  NAND2_X1 U18 ( .A1(n30), .A2(n47), .ZN(mask_sh3[23]) );
  NAND2_X1 U19 ( .A1(n32), .A2(n49), .ZN(mask_sh3[22]) );
  NAND2_X1 U20 ( .A1(n22), .A2(n42), .ZN(mask_sh2[26]) );
  NAND2_X1 U21 ( .A1(n23), .A2(n44), .ZN(mask_sh2[25]) );
  NAND2_X1 U22 ( .A1(n34), .A2(n38), .ZN(mask_sh6[24]) );
  NAND2_X1 U23 ( .A1(n26), .A2(n42), .ZN(mask_sh3[25]) );
  NAND2_X1 U24 ( .A1(n28), .A2(n44), .ZN(mask_sh3[24]) );
  NAND2_X1 U25 ( .A1(n37), .A2(n40), .ZN(mask_sh6[23]) );
  NAND2_X1 U26 ( .A1(n22), .A2(n38), .ZN(mask_sh3[27]) );
  NAND2_X1 U27 ( .A1(n23), .A2(n40), .ZN(mask_sh3[26]) );
  NAND2_X1 U28 ( .A1(n8), .A2(n13), .ZN(mask_sh6[8]) );
  NAND2_X1 U29 ( .A1(n10), .A2(n14), .ZN(mask_sh6[7]) );
  NAND2_X1 U30 ( .A1(n8), .A2(n46), .ZN(mask_sh3[5]) );
  NAND2_X1 U31 ( .A1(n11), .A2(n54), .ZN(mask_sh3[12]) );
  NAND2_X1 U32 ( .A1(n16), .A2(n60), .ZN(mask_sh3[9]) );
  NAND2_X1 U33 ( .A1(n14), .A2(n58), .ZN(mask_sh3[10]) );
  NAND2_X1 U34 ( .A1(n20), .A2(n63), .ZN(mask_sh3[7]) );
  NAND2_X1 U35 ( .A1(n18), .A2(n61), .ZN(mask_sh3[8]) );
  NAND2_X1 U36 ( .A1(n24), .A2(n65), .ZN(mask_sh3[6]) );
  NAND2_X1 U37 ( .A1(n13), .A2(n56), .ZN(mask_sh3[11]) );
  NAND2_X1 U38 ( .A1(n38), .A2(n70), .ZN(mask_sh2[28]) );
  NAND2_X1 U39 ( .A1(n40), .A2(n68), .ZN(mask_sh2[27]) );
  NAND2_X1 U40 ( .A1(n36), .A2(n73), .ZN(mask_sh2[29]) );
  NAND2_X1 U41 ( .A1(n36), .A2(n68), .ZN(mask_sh3[28]) );
  NAND2_X1 U42 ( .A1(n30), .A2(n35), .ZN(mask_sh6[26]) );
  NAND2_X1 U43 ( .A1(n22), .A2(n27), .ZN(mask_sh6[30]) );
  NAND2_X1 U44 ( .A1(n23), .A2(n29), .ZN(mask_sh6[29]) );
  NAND2_X1 U45 ( .A1(n26), .A2(n31), .ZN(mask_sh6[28]) );
  NAND2_X1 U46 ( .A1(n28), .A2(n33), .ZN(mask_sh6[27]) );
  NAND2_X1 U47 ( .A1(n54), .A2(n62), .ZN(mask_sh5[14]) );
  NAND2_X1 U48 ( .A1(n56), .A2(n64), .ZN(mask_sh5[13]) );
  NAND2_X1 U49 ( .A1(n58), .A2(n66), .ZN(mask_sh5[12]) );
  NAND2_X1 U50 ( .A1(n65), .A2(n66), .ZN(mask_sh7[10]) );
  NAND2_X1 U51 ( .A1(n43), .A2(n51), .ZN(mask_sh5[19]) );
  NAND2_X1 U52 ( .A1(n45), .A2(n53), .ZN(mask_sh5[18]) );
  NAND2_X1 U53 ( .A1(n48), .A2(n55), .ZN(mask_sh5[17]) );
  NAND2_X1 U54 ( .A1(n50), .A2(n57), .ZN(mask_sh5[16]) );
  NAND2_X1 U55 ( .A1(n52), .A2(n59), .ZN(mask_sh5[15]) );
  NAND2_X1 U56 ( .A1(n39), .A2(n47), .ZN(mask_sh5[21]) );
  NAND2_X1 U57 ( .A1(n41), .A2(n49), .ZN(mask_sh5[20]) );
  NAND2_X1 U58 ( .A1(n34), .A2(n42), .ZN(mask_sh5[23]) );
  NAND2_X1 U59 ( .A1(n37), .A2(n44), .ZN(mask_sh5[22]) );
  NAND2_X1 U60 ( .A1(n30), .A2(n38), .ZN(mask_sh5[25]) );
  NAND2_X1 U61 ( .A1(n32), .A2(n40), .ZN(mask_sh5[24]) );
  NAND2_X1 U62 ( .A1(n8), .A2(n16), .ZN(mask_sh5[7]) );
  NAND2_X1 U63 ( .A1(n12), .A2(n20), .ZN(mask_sh5[5]) );
  NAND2_X1 U64 ( .A1(n8), .A2(n9), .ZN(mask_sh7[9]) );
  NAND2_X1 U65 ( .A1(n10), .A2(n18), .ZN(mask_sh5[6]) );
  NAND2_X1 U66 ( .A1(n9), .A2(n60), .ZN(mask_sh5[11]) );
  NAND2_X1 U67 ( .A1(n47), .A2(n48), .ZN(mask_sh7[19]) );
  NAND2_X1 U68 ( .A1(n49), .A2(n50), .ZN(mask_sh7[18]) );
  NAND2_X1 U69 ( .A1(n13), .A2(n63), .ZN(mask_sh5[9]) );
  NAND2_X1 U70 ( .A1(n42), .A2(n43), .ZN(mask_sh7[21]) );
  NAND2_X1 U71 ( .A1(n44), .A2(n45), .ZN(mask_sh7[20]) );
  NAND2_X1 U72 ( .A1(n11), .A2(n61), .ZN(mask_sh5[10]) );
  NAND2_X1 U73 ( .A1(n14), .A2(n65), .ZN(mask_sh5[8]) );
  NAND2_X1 U74 ( .A1(n40), .A2(n41), .ZN(mask_sh7[22]) );
  NAND2_X1 U75 ( .A1(n26), .A2(n35), .ZN(mask_sh5[27]) );
  NAND2_X1 U76 ( .A1(n34), .A2(n35), .ZN(mask_sh7[25]) );
  NAND2_X1 U77 ( .A1(n22), .A2(n31), .ZN(mask_sh5[29]) );
  NAND2_X1 U78 ( .A1(n23), .A2(n33), .ZN(mask_sh5[28]) );
  NAND2_X1 U79 ( .A1(n32), .A2(n33), .ZN(mask_sh7[26]) );
  NAND2_X1 U80 ( .A1(n68), .A2(n29), .ZN(mask_sh5[30]) );
  NAND2_X1 U81 ( .A1(n70), .A2(n27), .ZN(mask_sh5[31]) );
  NAND2_X1 U82 ( .A1(n41), .A2(n62), .ZN(mask_sh2[17]) );
  NAND2_X1 U83 ( .A1(n43), .A2(n64), .ZN(mask_sh2[16]) );
  NAND2_X1 U84 ( .A1(n45), .A2(n66), .ZN(mask_sh2[15]) );
  NAND2_X1 U85 ( .A1(n45), .A2(n62), .ZN(mask_sh3[16]) );
  NAND2_X1 U86 ( .A1(n48), .A2(n64), .ZN(mask_sh3[15]) );
  NAND2_X1 U87 ( .A1(n50), .A2(n66), .ZN(mask_sh3[14]) );
  NAND2_X1 U88 ( .A1(n41), .A2(n57), .ZN(mask_sh3[18]) );
  NAND2_X1 U89 ( .A1(n43), .A2(n59), .ZN(mask_sh3[17]) );
  NAND2_X1 U90 ( .A1(n13), .A2(n52), .ZN(mask_sh2[12]) );
  NAND2_X1 U91 ( .A1(n14), .A2(n54), .ZN(mask_sh2[11]) );
  NAND2_X1 U92 ( .A1(n20), .A2(n60), .ZN(mask_sh2[8]) );
  NAND2_X1 U93 ( .A1(n9), .A2(n48), .ZN(mask_sh2[14]) );
  NAND2_X1 U94 ( .A1(n11), .A2(n50), .ZN(mask_sh2[13]) );
  NAND2_X1 U95 ( .A1(n18), .A2(n58), .ZN(mask_sh2[9]) );
  NAND2_X1 U96 ( .A1(n46), .A2(n63), .ZN(mask_sh2[6]) );
  NAND2_X1 U97 ( .A1(n9), .A2(n52), .ZN(mask_sh3[13]) );
  NAND2_X1 U98 ( .A1(n24), .A2(n61), .ZN(mask_sh2[7]) );
  NAND2_X1 U99 ( .A1(n16), .A2(n56), .ZN(mask_sh2[10]) );
  NAND2_X1 U100 ( .A1(n35), .A2(n72), .ZN(mask_sh2[30]) );
  NAND2_X1 U101 ( .A1(n35), .A2(n70), .ZN(mask_sh3[29]) );
  NAND2_X1 U102 ( .A1(n33), .A2(n76), .ZN(mask_sh2[31]) );
  NAND2_X1 U103 ( .A1(n33), .A2(n73), .ZN(mask_sh3[30]) );
  NAND2_X1 U104 ( .A1(n31), .A2(n72), .ZN(mask_sh3[31]) );
  NAND2_X1 U105 ( .A1(\R1[19] ), .A2(n78), .ZN(n62) );
  NAND2_X1 U106 ( .A1(\R1[18] ), .A2(n78), .ZN(n64) );
  NAND2_X1 U107 ( .A1(\R1[17] ), .A2(n78), .ZN(n66) );
  NAND2_X1 U108 ( .A1(\R1[24] ), .A2(n7), .ZN(n51) );
  NAND2_X1 U109 ( .A1(\R1[23] ), .A2(n78), .ZN(n53) );
  NAND2_X1 U110 ( .A1(\R1[22] ), .A2(n78), .ZN(n55) );
  NAND2_X1 U111 ( .A1(\R1[21] ), .A2(n78), .ZN(n57) );
  NAND2_X1 U112 ( .A1(\R1[20] ), .A2(n78), .ZN(n59) );
  NAND2_X1 U113 ( .A1(\R1[26] ), .A2(n7), .ZN(n47) );
  NAND2_X1 U114 ( .A1(\R1[25] ), .A2(n78), .ZN(n49) );
  NAND2_X1 U115 ( .A1(n89), .A2(\R1[16] ), .ZN(n56) );
  NAND2_X1 U116 ( .A1(\R1[18] ), .A2(n79), .ZN(n52) );
  NAND2_X1 U117 ( .A1(\R1[17] ), .A2(n87), .ZN(n54) );
  NAND2_X1 U118 ( .A1(\R1[14] ), .A2(n87), .ZN(n60) );
  NAND2_X1 U119 ( .A1(\R1[28] ), .A2(n7), .ZN(n42) );
  NAND2_X1 U120 ( .A1(\R1[27] ), .A2(n78), .ZN(n44) );
  NAND2_X1 U121 ( .A1(\R1[30] ), .A2(n7), .ZN(n38) );
  NAND2_X1 U122 ( .A1(\R1[20] ), .A2(n79), .ZN(n48) );
  NAND2_X1 U123 ( .A1(\R1[19] ), .A2(n80), .ZN(n50) );
  NAND2_X1 U124 ( .A1(\R1[15] ), .A2(n86), .ZN(n58) );
  NAND2_X1 U125 ( .A1(\R1[12] ), .A2(n85), .ZN(n63) );
  NAND2_X1 U126 ( .A1(\R1[29] ), .A2(n78), .ZN(n40) );
  NAND2_X1 U127 ( .A1(\R1[31] ), .A2(n7), .ZN(n36) );
  NAND2_X1 U128 ( .A1(\R1[22] ), .A2(n81), .ZN(n43) );
  NAND2_X1 U129 ( .A1(\R1[21] ), .A2(n80), .ZN(n45) );
  NAND2_X1 U130 ( .A1(\R1[13] ), .A2(n86), .ZN(n61) );
  NAND2_X1 U131 ( .A1(\R1[11] ), .A2(n84), .ZN(n65) );
  NAND2_X1 U132 ( .A1(\R1[14] ), .A2(n78), .ZN(n13) );
  NAND2_X1 U133 ( .A1(\R1[12] ), .A2(n78), .ZN(n16) );
  NAND2_X1 U134 ( .A1(\R1[8] ), .A2(n78), .ZN(n46) );
  NAND2_X1 U135 ( .A1(\R1[24] ), .A2(n81), .ZN(n39) );
  NAND2_X1 U136 ( .A1(\R1[23] ), .A2(n81), .ZN(n41) );
  NAND2_X1 U137 ( .A1(\R1[10] ), .A2(n7), .ZN(n20) );
  NAND2_X1 U138 ( .A1(\R1[16] ), .A2(n78), .ZN(n9) );
  NAND2_X1 U139 ( .A1(\R1[15] ), .A2(n78), .ZN(n11) );
  NAND2_X1 U140 ( .A1(\R1[13] ), .A2(n78), .ZN(n14) );
  NAND2_X1 U141 ( .A1(\R1[11] ), .A2(n78), .ZN(n18) );
  NAND2_X1 U142 ( .A1(\R1[9] ), .A2(n7), .ZN(n24) );
  NAND2_X1 U143 ( .A1(\R1[25] ), .A2(n82), .ZN(n37) );
  NAND2_X1 U144 ( .A1(\R1[32] ), .A2(n82), .ZN(n22) );
  NAND2_X1 U145 ( .A1(\R1[31] ), .A2(n83), .ZN(n23) );
  NAND2_X1 U146 ( .A1(\R1[9] ), .A2(n83), .ZN(n10) );
  NAND2_X1 U147 ( .A1(\R1[8] ), .A2(n80), .ZN(n12) );
  NAND2_X1 U148 ( .A1(\R1[30] ), .A2(n84), .ZN(n26) );
  NAND2_X1 U149 ( .A1(\R1[29] ), .A2(n83), .ZN(n28) );
  NAND2_X1 U150 ( .A1(\R1[28] ), .A2(n82), .ZN(n30) );
  NAND2_X1 U151 ( .A1(\R1[27] ), .A2(n81), .ZN(n32) );
  NAND2_X1 U152 ( .A1(\R1[26] ), .A2(n82), .ZN(n34) );
  NAND2_X1 U153 ( .A1(\R1[10] ), .A2(n86), .ZN(n8) );
  NAND2_X1 U154 ( .A1(\R1[32] ), .A2(n7), .ZN(n35) );
  NAND2_X1 U155 ( .A1(\R1[33] ), .A2(n84), .ZN(n68) );
  NAND2_X1 U156 ( .A1(\R1[33] ), .A2(n7), .ZN(n33) );
  NAND2_X1 U157 ( .A1(\R1[34] ), .A2(n84), .ZN(n70) );
  NAND2_X1 U158 ( .A1(\R1[34] ), .A2(n7), .ZN(n31) );
  NAND2_X1 U159 ( .A1(R1[36]), .A2(n7), .ZN(n27) );
  NAND2_X1 U160 ( .A1(\R1[35] ), .A2(n7), .ZN(n29) );
  OAI21_X1 U161 ( .B1(n88), .B2(n93), .A(n68), .ZN(mask_sh6[31]) );
  NAND2_X1 U162 ( .A1(n43), .A2(n47), .ZN(mask_sh6[20]) );
  NAND2_X1 U163 ( .A1(n45), .A2(n49), .ZN(mask_sh6[19]) );
  NAND2_X1 U164 ( .A1(n10), .A2(n67), .ZN(mask_sh3[4]) );
  NAND2_X1 U165 ( .A1(n12), .A2(n16), .ZN(mask_sh6[6]) );
  NAND2_X1 U166 ( .A1(n9), .A2(n63), .ZN(mask_sh6[10]) );
  NAND2_X1 U167 ( .A1(n11), .A2(n65), .ZN(mask_sh6[9]) );
  NAND2_X1 U168 ( .A1(n46), .A2(n21), .ZN(mask_sh6[2]) );
  NAND2_X1 U169 ( .A1(n20), .A2(n17), .ZN(mask_sh6[4]) );
  NAND2_X1 U170 ( .A1(n18), .A2(n15), .ZN(mask_sh6[5]) );
  NAND2_X1 U171 ( .A1(n12), .A2(n69), .ZN(mask_sh3[3]) );
  NAND2_X1 U172 ( .A1(n24), .A2(n19), .ZN(mask_sh6[3]) );
  INV_X1 U173 ( .A(R1[37]), .ZN(n93) );
  NAND2_X1 U174 ( .A1(n39), .A2(n42), .ZN(mask_sh6[22]) );
  NAND2_X1 U175 ( .A1(n41), .A2(n44), .ZN(mask_sh6[21]) );
  NAND2_X1 U176 ( .A1(n48), .A2(n51), .ZN(mask_sh6[18]) );
  NAND2_X1 U177 ( .A1(n32), .A2(n36), .ZN(mask_sh6[25]) );
  NAND2_X1 U178 ( .A1(n46), .A2(n17), .ZN(mask_sh5[3]) );
  NAND2_X1 U179 ( .A1(n14), .A2(n15), .ZN(mask_sh7[6]) );
  NAND2_X1 U180 ( .A1(n24), .A2(n15), .ZN(mask_sh5[4]) );
  NAND2_X1 U181 ( .A1(R1[36]), .A2(n85), .ZN(n72) );
  NAND2_X1 U182 ( .A1(\R1[35] ), .A2(n85), .ZN(n73) );
  OAI21_X1 U183 ( .B1(n95), .B2(n78), .A(n36), .ZN(mask_sh0[31]) );
  INV_X1 U184 ( .A(R1[39]), .ZN(n95) );
  OAI21_X1 U185 ( .B1(n78), .B2(n94), .A(n38), .ZN(mask_sh0[30]) );
  NAND2_X1 U186 ( .A1(n40), .A2(n76), .ZN(mask_sh0[29]) );
  NAND2_X1 U187 ( .A1(n42), .A2(n72), .ZN(mask_sh0[28]) );
  NAND2_X1 U188 ( .A1(n44), .A2(n73), .ZN(mask_sh0[27]) );
  NAND2_X1 U189 ( .A1(n47), .A2(n70), .ZN(mask_sh0[26]) );
  NAND2_X1 U190 ( .A1(n49), .A2(n68), .ZN(mask_sh0[25]) );
  NAND2_X1 U191 ( .A1(n22), .A2(n51), .ZN(mask_sh0[24]) );
  NAND2_X1 U192 ( .A1(n23), .A2(n53), .ZN(mask_sh0[23]) );
  NAND2_X1 U193 ( .A1(n26), .A2(n55), .ZN(mask_sh0[22]) );
  NAND2_X1 U194 ( .A1(n28), .A2(n57), .ZN(mask_sh0[21]) );
  NAND2_X1 U195 ( .A1(n30), .A2(n59), .ZN(mask_sh0[20]) );
  NAND2_X1 U196 ( .A1(n32), .A2(n62), .ZN(mask_sh0[19]) );
  NAND2_X1 U197 ( .A1(n34), .A2(n64), .ZN(mask_sh0[18]) );
  NAND2_X1 U198 ( .A1(n9), .A2(n39), .ZN(mask_sh0[16]) );
  NAND2_X1 U199 ( .A1(n11), .A2(n41), .ZN(mask_sh0[15]) );
  NAND2_X1 U200 ( .A1(n13), .A2(n43), .ZN(mask_sh0[14]) );
  NAND2_X1 U201 ( .A1(n14), .A2(n45), .ZN(mask_sh0[13]) );
  NAND2_X1 U202 ( .A1(n16), .A2(n48), .ZN(mask_sh0[12]) );
  NAND2_X1 U203 ( .A1(n18), .A2(n50), .ZN(mask_sh0[11]) );
  NAND2_X1 U204 ( .A1(n20), .A2(n52), .ZN(mask_sh0[10]) );
  NAND2_X1 U205 ( .A1(n24), .A2(n54), .ZN(mask_sh0[9]) );
  NAND2_X1 U206 ( .A1(n46), .A2(n56), .ZN(mask_sh0[8]) );
  NAND2_X1 U207 ( .A1(n58), .A2(n67), .ZN(mask_sh0[7]) );
  NAND2_X1 U208 ( .A1(n60), .A2(n69), .ZN(mask_sh0[6]) );
  NAND2_X1 U209 ( .A1(n61), .A2(n71), .ZN(mask_sh0[5]) );
  NAND2_X1 U210 ( .A1(n63), .A2(n74), .ZN(mask_sh0[4]) );
  NAND2_X1 U211 ( .A1(n65), .A2(n75), .ZN(mask_sh0[3]) );
  NAND2_X1 U212 ( .A1(n8), .A2(n77), .ZN(mask_sh0[2]) );
  OAI21_X1 U213 ( .B1(n7), .B2(n92), .A(n69), .ZN(mask_sh6[0]) );
  NAND2_X1 U214 ( .A1(R1[37]), .A2(n85), .ZN(n76) );
  NAND2_X1 U215 ( .A1(n37), .A2(n66), .ZN(mask_sh0[17]) );
  NAND2_X1 U216 ( .A1(n65), .A2(n67), .ZN(mask_sh2[5]) );
  NAND2_X1 U217 ( .A1(n67), .A2(n25), .ZN(mask_sh6[1]) );
  NAND2_X1 U218 ( .A1(n8), .A2(n69), .ZN(mask_sh2[4]) );
  NAND2_X1 U219 ( .A1(n10), .A2(n71), .ZN(mask_sh2[3]) );
  NAND2_X1 U220 ( .A1(n12), .A2(n74), .ZN(mask_sh2[2]) );
  NAND2_X1 U221 ( .A1(n15), .A2(n71), .ZN(mask_sh3[2]) );
  NAND2_X1 U222 ( .A1(n15), .A2(n75), .ZN(mask_sh2[1]) );
  NAND2_X1 U223 ( .A1(n67), .A2(n19), .ZN(mask_sh5[2]) );
  NAND2_X1 U224 ( .A1(n17), .A2(n74), .ZN(mask_sh3[1]) );
  NAND2_X1 U225 ( .A1(n19), .A2(n75), .ZN(mask_sh3[0]) );
  NAND2_X1 U226 ( .A1(n17), .A2(n77), .ZN(mask_sh2[0]) );
  NAND2_X1 U227 ( .A1(n69), .A2(n21), .ZN(mask_sh5[1]) );
  NAND2_X1 U228 ( .A1(n71), .A2(n25), .ZN(mask_sh5[0]) );
  INV_X1 U229 ( .A(n88), .ZN(n7) );
  INV_X1 U230 ( .A(n89), .ZN(n78) );
  NAND2_X1 U231 ( .A1(\R1[7] ), .A2(n7), .ZN(n67) );
  NAND2_X1 U232 ( .A1(n28), .A2(n36), .ZN(mask_sh5[26]) );
  NAND2_X1 U233 ( .A1(n36), .A2(n37), .ZN(mask_sh7[24]) );
  NAND2_X1 U234 ( .A1(n38), .A2(n39), .ZN(mask_sh7[23]) );
  NAND2_X1 U235 ( .A1(n51), .A2(n52), .ZN(mask_sh7[17]) );
  NAND2_X1 U236 ( .A1(n53), .A2(n54), .ZN(mask_sh7[16]) );
  NAND2_X1 U237 ( .A1(n55), .A2(n56), .ZN(mask_sh7[15]) );
  NAND2_X1 U238 ( .A1(n57), .A2(n58), .ZN(mask_sh7[14]) );
  NAND2_X1 U239 ( .A1(n59), .A2(n60), .ZN(mask_sh7[13]) );
  NAND2_X1 U240 ( .A1(n61), .A2(n62), .ZN(mask_sh7[12]) );
  NAND2_X1 U241 ( .A1(n63), .A2(n64), .ZN(mask_sh7[11]) );
  NAND2_X1 U242 ( .A1(n10), .A2(n11), .ZN(mask_sh7[8]) );
  NAND2_X1 U243 ( .A1(n12), .A2(n13), .ZN(mask_sh7[7]) );
  NAND2_X1 U244 ( .A1(n16), .A2(n17), .ZN(mask_sh7[5]) );
  NAND2_X1 U245 ( .A1(n18), .A2(n19), .ZN(mask_sh7[4]) );
  NAND2_X1 U246 ( .A1(n20), .A2(n21), .ZN(mask_sh7[3]) );
  NAND2_X1 U247 ( .A1(n24), .A2(n25), .ZN(mask_sh7[2]) );
  OAI21_X1 U248 ( .B1(n78), .B2(n92), .A(n46), .ZN(mask_sh7[1]) );
  OAI21_X1 U249 ( .B1(n88), .B2(n94), .A(n22), .ZN(mask_sh7[31]) );
  OAI21_X1 U250 ( .B1(n87), .B2(n93), .A(n23), .ZN(mask_sh7[30]) );
  NAND2_X1 U251 ( .A1(n26), .A2(n27), .ZN(mask_sh7[29]) );
  NAND2_X1 U252 ( .A1(n28), .A2(n29), .ZN(mask_sh7[28]) );
  NAND2_X1 U253 ( .A1(n30), .A2(n31), .ZN(mask_sh7[27]) );
  OAI21_X1 U254 ( .B1(n78), .B2(n91), .A(n67), .ZN(mask_sh7[0]) );
  NAND2_X1 U255 ( .A1(n23), .A2(n49), .ZN(mask_sh1[24]) );
  NAND2_X1 U256 ( .A1(n26), .A2(n51), .ZN(mask_sh1[23]) );
  NAND2_X1 U257 ( .A1(n28), .A2(n53), .ZN(mask_sh1[22]) );
  NAND2_X1 U258 ( .A1(n30), .A2(n55), .ZN(mask_sh1[21]) );
  NAND2_X1 U259 ( .A1(n32), .A2(n57), .ZN(mask_sh1[20]) );
  NAND2_X1 U260 ( .A1(n34), .A2(n59), .ZN(mask_sh1[19]) );
  NAND2_X1 U261 ( .A1(n37), .A2(n62), .ZN(mask_sh1[18]) );
  NAND2_X1 U262 ( .A1(n39), .A2(n64), .ZN(mask_sh1[17]) );
  NAND2_X1 U263 ( .A1(n41), .A2(n66), .ZN(mask_sh1[16]) );
  NAND2_X1 U264 ( .A1(n9), .A2(n43), .ZN(mask_sh1[15]) );
  NAND2_X1 U265 ( .A1(n11), .A2(n45), .ZN(mask_sh1[14]) );
  NAND2_X1 U266 ( .A1(n13), .A2(n48), .ZN(mask_sh1[13]) );
  NAND2_X1 U267 ( .A1(n14), .A2(n50), .ZN(mask_sh1[12]) );
  NAND2_X1 U268 ( .A1(n16), .A2(n52), .ZN(mask_sh1[11]) );
  NAND2_X1 U269 ( .A1(n18), .A2(n54), .ZN(mask_sh1[10]) );
  NAND2_X1 U270 ( .A1(n20), .A2(n56), .ZN(mask_sh1[9]) );
  NAND2_X1 U271 ( .A1(n24), .A2(n58), .ZN(mask_sh1[8]) );
  NAND2_X1 U272 ( .A1(n46), .A2(n60), .ZN(mask_sh1[7]) );
  NAND2_X1 U273 ( .A1(n61), .A2(n67), .ZN(mask_sh1[6]) );
  NAND2_X1 U274 ( .A1(n63), .A2(n69), .ZN(mask_sh1[5]) );
  NAND2_X1 U275 ( .A1(n65), .A2(n71), .ZN(mask_sh1[4]) );
  NAND2_X1 U276 ( .A1(n8), .A2(n74), .ZN(mask_sh1[3]) );
  NAND2_X1 U277 ( .A1(n10), .A2(n75), .ZN(mask_sh1[2]) );
  NAND2_X1 U278 ( .A1(n12), .A2(n77), .ZN(mask_sh1[1]) );
  OAI21_X1 U279 ( .B1(n7), .B2(n94), .A(n35), .ZN(mask_sh1[31]) );
  NAND2_X1 U280 ( .A1(n36), .A2(n76), .ZN(mask_sh1[30]) );
  NAND2_X1 U281 ( .A1(n38), .A2(n72), .ZN(mask_sh1[29]) );
  NAND2_X1 U282 ( .A1(n40), .A2(n73), .ZN(mask_sh1[28]) );
  NAND2_X1 U283 ( .A1(n42), .A2(n70), .ZN(mask_sh1[27]) );
  NAND2_X1 U284 ( .A1(n44), .A2(n68), .ZN(mask_sh1[26]) );
  NAND2_X1 U285 ( .A1(n22), .A2(n47), .ZN(mask_sh1[25]) );
  OAI21_X1 U286 ( .B1(n88), .B2(n90), .A(n12), .ZN(mask_sh0[0]) );
  INV_X1 U287 ( .A(R1[38]), .ZN(n94) );
  NAND2_X1 U288 ( .A1(\R1[6] ), .A2(n7), .ZN(n69) );
  NAND2_X1 U289 ( .A1(\R1[7] ), .A2(n86), .ZN(n15) );
  NAND2_X1 U290 ( .A1(\R1[5] ), .A2(n7), .ZN(n71) );
  NAND2_X1 U291 ( .A1(\R1[6] ), .A2(n83), .ZN(n17) );
  NAND2_X1 U292 ( .A1(\R1[4] ), .A2(n7), .ZN(n74) );
  NAND2_X1 U293 ( .A1(R1_3), .A2(n7), .ZN(n75) );
  NAND2_X1 U294 ( .A1(\R1[5] ), .A2(n80), .ZN(n19) );
  NAND2_X1 U295 ( .A1(R1_2), .A2(n7), .ZN(n77) );
  OAI21_X1 U296 ( .B1(n88), .B2(n91), .A(n10), .ZN(mask_sh0[1]) );
  NAND2_X1 U297 ( .A1(\R1[4] ), .A2(n79), .ZN(n21) );
  NAND2_X1 U298 ( .A1(R1_3), .A2(n79), .ZN(n25) );
  OAI21_X1 U299 ( .B1(n87), .B2(n91), .A(n15), .ZN(mask_sh1[0]) );
  INV_X1 U300 ( .A(R1_2), .ZN(n92) );
  BUF_X1 U301 ( .A(n4), .Z(n88) );
  BUF_X1 U302 ( .A(n2), .Z(n82) );
  BUF_X1 U303 ( .A(n1), .Z(n81) );
  BUF_X1 U304 ( .A(n1), .Z(n79) );
  BUF_X1 U305 ( .A(n3), .Z(n85) );
  BUF_X1 U306 ( .A(n2), .Z(n84) );
  BUF_X1 U307 ( .A(n3), .Z(n86) );
  BUF_X1 U308 ( .A(n2), .Z(n83) );
  BUF_X1 U309 ( .A(n1), .Z(n80) );
  BUF_X1 U310 ( .A(n3), .Z(n87) );
  BUF_X1 U311 ( .A(n4), .Z(n89) );
  INV_X1 U312 ( .A(R1_1), .ZN(n91) );
  INV_X1 U313 ( .A(R1_0), .ZN(n90) );
  BUF_X1 U314 ( .A(n5), .Z(n3) );
  BUF_X1 U315 ( .A(n6), .Z(n2) );
  BUF_X1 U316 ( .A(n6), .Z(n1) );
  BUF_X1 U317 ( .A(n5), .Z(n4) );
  BUF_X1 U318 ( .A(LnR), .Z(n5) );
  BUF_X1 U319 ( .A(LnR), .Z(n6) );
endmodule


module MUX81_0 ( A, B, C, D, E, F, G, H, S, Y );
  input [2:0] S;
  input A, B, C, D, E, F, G, H;
  output Y;
  wire   n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n1,
         n2, n3, n4, n5, n6;

  NAND3_X1 U20 ( .A1(S[1]), .A2(n6), .A3(H), .ZN(n19) );
  NAND3_X1 U21 ( .A1(S[0]), .A2(n2), .A3(F), .ZN(n17) );
  INV_X1 U1 ( .A(n15), .ZN(n5) );
  NOR2_X1 U2 ( .A1(n1), .A2(S[2]), .ZN(n15) );
  INV_X1 U3 ( .A(n10), .ZN(n4) );
  INV_X1 U4 ( .A(n20), .ZN(n6) );
  NAND2_X1 U5 ( .A1(n7), .A2(n8), .ZN(Y) );
  NAND4_X1 U6 ( .A1(A), .A2(n1), .A3(n2), .A4(n3), .ZN(n8) );
  AOI22_X1 U7 ( .A1(n9), .A2(n4), .B1(B), .B2(n10), .ZN(n7) );
  OAI21_X1 U8 ( .B1(n11), .B2(n12), .A(n13), .ZN(n9) );
  NAND2_X1 U9 ( .A1(C), .A2(n12), .ZN(n13) );
  AOI22_X1 U10 ( .A1(n14), .A2(n5), .B1(D), .B2(n15), .ZN(n11) );
  NOR3_X1 U11 ( .A1(S[0]), .A2(S[2]), .A3(n2), .ZN(n12) );
  NAND4_X1 U12 ( .A1(n16), .A2(n17), .A3(n18), .A4(n19), .ZN(n14) );
  NAND4_X1 U13 ( .A1(E), .A2(S[2]), .A3(n1), .A4(n2), .ZN(n16) );
  NAND2_X1 U14 ( .A1(G), .A2(n20), .ZN(n18) );
  NOR3_X1 U15 ( .A1(S[1]), .A2(S[2]), .A3(n1), .ZN(n10) );
  NOR2_X1 U16 ( .A1(n2), .A2(S[0]), .ZN(n20) );
  INV_X1 U17 ( .A(S[0]), .ZN(n1) );
  INV_X1 U18 ( .A(S[1]), .ZN(n2) );
  INV_X1 U19 ( .A(S[2]), .ZN(n3) );
endmodule


module MUX81_31 ( A, B, C, D, E, F, G, H, S, Y );
  input [2:0] S;
  input A, B, C, D, E, F, G, H;
  output Y;
  wire   n1, n2, n3, n4, n5, n6, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35;

  NAND3_X1 U20 ( .A1(S[1]), .A2(n21), .A3(H), .ZN(n23) );
  NAND3_X1 U21 ( .A1(S[0]), .A2(n2), .A3(F), .ZN(n25) );
  INV_X1 U1 ( .A(n27), .ZN(n6) );
  NOR2_X1 U2 ( .A1(n1), .A2(n3), .ZN(n27) );
  INV_X1 U3 ( .A(n22), .ZN(n21) );
  AOI22_X1 U4 ( .A1(n33), .A2(n5), .B1(B), .B2(n32), .ZN(n35) );
  INV_X1 U5 ( .A(n32), .ZN(n5) );
  NOR3_X1 U6 ( .A1(S[1]), .A2(n3), .A3(n1), .ZN(n32) );
  OAI21_X1 U7 ( .B1(n31), .B2(n30), .A(n29), .ZN(n33) );
  NAND2_X1 U8 ( .A1(C), .A2(n30), .ZN(n29) );
  AOI22_X1 U9 ( .A1(n28), .A2(n6), .B1(D), .B2(n27), .ZN(n31) );
  NOR3_X1 U10 ( .A1(S[0]), .A2(n3), .A3(n2), .ZN(n30) );
  NAND4_X1 U11 ( .A1(n26), .A2(n25), .A3(n24), .A4(n23), .ZN(n28) );
  NAND4_X1 U12 ( .A1(E), .A2(n3), .A3(n1), .A4(n2), .ZN(n26) );
  NAND2_X1 U13 ( .A1(G), .A2(n22), .ZN(n24) );
  NAND2_X1 U14 ( .A1(n35), .A2(n34), .ZN(Y) );
  NOR2_X1 U15 ( .A1(n2), .A2(S[0]), .ZN(n22) );
  NAND4_X1 U16 ( .A1(A), .A2(n1), .A3(n2), .A4(n4), .ZN(n34) );
  INV_X1 U17 ( .A(S[0]), .ZN(n1) );
  INV_X1 U18 ( .A(S[1]), .ZN(n2) );
  INV_X1 U19 ( .A(n4), .ZN(n3) );
  INV_X1 U22 ( .A(S[2]), .ZN(n4) );
endmodule


module MUX81_30 ( A, B, C, D, E, F, G, H, S, Y );
  input [2:0] S;
  input A, B, C, D, E, F, G, H;
  output Y;
  wire   n1, n2, n3, n4, n5, n6, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35;

  NAND3_X1 U20 ( .A1(S[1]), .A2(n21), .A3(H), .ZN(n23) );
  NAND3_X1 U21 ( .A1(S[0]), .A2(n2), .A3(F), .ZN(n25) );
  INV_X1 U1 ( .A(n27), .ZN(n6) );
  NOR2_X1 U2 ( .A1(n1), .A2(n3), .ZN(n27) );
  NAND4_X1 U3 ( .A1(A), .A2(n1), .A3(n2), .A4(n4), .ZN(n34) );
  INV_X1 U4 ( .A(n22), .ZN(n21) );
  AOI22_X1 U5 ( .A1(n33), .A2(n5), .B1(B), .B2(n32), .ZN(n35) );
  INV_X1 U6 ( .A(n32), .ZN(n5) );
  NOR3_X1 U7 ( .A1(S[1]), .A2(n3), .A3(n1), .ZN(n32) );
  OAI21_X1 U8 ( .B1(n31), .B2(n30), .A(n29), .ZN(n33) );
  NAND2_X1 U9 ( .A1(C), .A2(n30), .ZN(n29) );
  AOI22_X1 U10 ( .A1(n28), .A2(n6), .B1(D), .B2(n27), .ZN(n31) );
  NOR3_X1 U11 ( .A1(S[0]), .A2(n3), .A3(n2), .ZN(n30) );
  NAND4_X1 U12 ( .A1(n26), .A2(n25), .A3(n24), .A4(n23), .ZN(n28) );
  NAND4_X1 U13 ( .A1(E), .A2(n3), .A3(n1), .A4(n2), .ZN(n26) );
  NAND2_X1 U14 ( .A1(G), .A2(n22), .ZN(n24) );
  NAND2_X1 U15 ( .A1(n35), .A2(n34), .ZN(Y) );
  NOR2_X1 U16 ( .A1(n2), .A2(S[0]), .ZN(n22) );
  INV_X1 U17 ( .A(S[0]), .ZN(n1) );
  INV_X1 U18 ( .A(S[1]), .ZN(n2) );
  INV_X1 U19 ( .A(n4), .ZN(n3) );
  INV_X1 U22 ( .A(S[2]), .ZN(n4) );
endmodule


module MUX81_29 ( A, B, C, D, E, F, G, H, S, Y );
  input [2:0] S;
  input A, B, C, D, E, F, G, H;
  output Y;
  wire   n1, n2, n3, n4, n5, n6, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35;

  NAND3_X1 U20 ( .A1(S[1]), .A2(n21), .A3(H), .ZN(n23) );
  NAND3_X1 U21 ( .A1(S[0]), .A2(n2), .A3(F), .ZN(n25) );
  INV_X1 U1 ( .A(n27), .ZN(n6) );
  NOR2_X1 U2 ( .A1(n1), .A2(n3), .ZN(n27) );
  NAND4_X1 U3 ( .A1(A), .A2(n1), .A3(n2), .A4(n4), .ZN(n34) );
  INV_X1 U4 ( .A(n22), .ZN(n21) );
  AOI22_X1 U5 ( .A1(n33), .A2(n5), .B1(B), .B2(n32), .ZN(n35) );
  INV_X1 U6 ( .A(n32), .ZN(n5) );
  NOR3_X1 U7 ( .A1(S[1]), .A2(n3), .A3(n1), .ZN(n32) );
  OAI21_X1 U8 ( .B1(n31), .B2(n30), .A(n29), .ZN(n33) );
  NAND2_X1 U9 ( .A1(C), .A2(n30), .ZN(n29) );
  AOI22_X1 U10 ( .A1(n28), .A2(n6), .B1(D), .B2(n27), .ZN(n31) );
  NOR3_X1 U11 ( .A1(S[0]), .A2(n3), .A3(n2), .ZN(n30) );
  NAND4_X1 U12 ( .A1(n26), .A2(n25), .A3(n24), .A4(n23), .ZN(n28) );
  NAND4_X1 U13 ( .A1(E), .A2(n3), .A3(n1), .A4(n2), .ZN(n26) );
  NAND2_X1 U14 ( .A1(G), .A2(n22), .ZN(n24) );
  NAND2_X1 U15 ( .A1(n35), .A2(n34), .ZN(Y) );
  NOR2_X1 U16 ( .A1(n2), .A2(S[0]), .ZN(n22) );
  INV_X1 U17 ( .A(S[0]), .ZN(n1) );
  INV_X1 U18 ( .A(S[1]), .ZN(n2) );
  INV_X1 U19 ( .A(n4), .ZN(n3) );
  INV_X1 U22 ( .A(S[2]), .ZN(n4) );
endmodule


module MUX81_28 ( A, B, C, D, E, F, G, H, S, Y );
  input [2:0] S;
  input A, B, C, D, E, F, G, H;
  output Y;
  wire   n1, n2, n3, n4, n5, n6, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35;

  NAND3_X1 U20 ( .A1(S[1]), .A2(n21), .A3(H), .ZN(n23) );
  NAND3_X1 U21 ( .A1(S[0]), .A2(n2), .A3(F), .ZN(n25) );
  INV_X1 U1 ( .A(n27), .ZN(n6) );
  NOR2_X1 U2 ( .A1(n1), .A2(n3), .ZN(n27) );
  NAND4_X1 U3 ( .A1(A), .A2(n1), .A3(n2), .A4(n4), .ZN(n34) );
  INV_X1 U4 ( .A(n22), .ZN(n21) );
  AOI22_X1 U5 ( .A1(n33), .A2(n5), .B1(B), .B2(n32), .ZN(n35) );
  INV_X1 U6 ( .A(n32), .ZN(n5) );
  NOR3_X1 U7 ( .A1(S[1]), .A2(n3), .A3(n1), .ZN(n32) );
  OAI21_X1 U8 ( .B1(n31), .B2(n30), .A(n29), .ZN(n33) );
  NAND2_X1 U9 ( .A1(C), .A2(n30), .ZN(n29) );
  AOI22_X1 U10 ( .A1(n28), .A2(n6), .B1(D), .B2(n27), .ZN(n31) );
  NOR3_X1 U11 ( .A1(S[0]), .A2(n3), .A3(n2), .ZN(n30) );
  NAND4_X1 U12 ( .A1(n26), .A2(n25), .A3(n24), .A4(n23), .ZN(n28) );
  NAND4_X1 U13 ( .A1(E), .A2(n3), .A3(n1), .A4(n2), .ZN(n26) );
  NAND2_X1 U14 ( .A1(G), .A2(n22), .ZN(n24) );
  NOR2_X1 U15 ( .A1(n2), .A2(S[0]), .ZN(n22) );
  NAND2_X1 U16 ( .A1(n35), .A2(n34), .ZN(Y) );
  INV_X1 U17 ( .A(S[0]), .ZN(n1) );
  INV_X1 U18 ( .A(S[1]), .ZN(n2) );
  INV_X1 U19 ( .A(n4), .ZN(n3) );
  INV_X1 U22 ( .A(S[2]), .ZN(n4) );
endmodule


module MUX81_27 ( A, B, C, D, E, F, G, H, S, Y );
  input [2:0] S;
  input A, B, C, D, E, F, G, H;
  output Y;
  wire   n1, n2, n3, n4, n5, n6, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35;

  NAND3_X1 U20 ( .A1(S[1]), .A2(n21), .A3(H), .ZN(n23) );
  NAND3_X1 U21 ( .A1(S[0]), .A2(n2), .A3(F), .ZN(n25) );
  INV_X1 U1 ( .A(n27), .ZN(n6) );
  NOR2_X1 U2 ( .A1(n1), .A2(n3), .ZN(n27) );
  NAND4_X1 U3 ( .A1(A), .A2(n1), .A3(n2), .A4(n4), .ZN(n34) );
  INV_X1 U4 ( .A(n22), .ZN(n21) );
  AOI22_X1 U5 ( .A1(n33), .A2(n5), .B1(B), .B2(n32), .ZN(n35) );
  INV_X1 U6 ( .A(n32), .ZN(n5) );
  NOR3_X1 U7 ( .A1(S[1]), .A2(n3), .A3(n1), .ZN(n32) );
  OAI21_X1 U8 ( .B1(n31), .B2(n30), .A(n29), .ZN(n33) );
  NAND2_X1 U9 ( .A1(C), .A2(n30), .ZN(n29) );
  AOI22_X1 U10 ( .A1(n28), .A2(n6), .B1(D), .B2(n27), .ZN(n31) );
  NOR3_X1 U11 ( .A1(S[0]), .A2(n3), .A3(n2), .ZN(n30) );
  NAND4_X1 U12 ( .A1(n26), .A2(n25), .A3(n24), .A4(n23), .ZN(n28) );
  NAND4_X1 U13 ( .A1(E), .A2(n3), .A3(n1), .A4(n2), .ZN(n26) );
  NAND2_X1 U14 ( .A1(G), .A2(n22), .ZN(n24) );
  NAND2_X1 U15 ( .A1(n35), .A2(n34), .ZN(Y) );
  NOR2_X1 U16 ( .A1(n2), .A2(S[0]), .ZN(n22) );
  INV_X1 U17 ( .A(S[0]), .ZN(n1) );
  INV_X1 U18 ( .A(S[1]), .ZN(n2) );
  INV_X1 U19 ( .A(n4), .ZN(n3) );
  INV_X1 U22 ( .A(S[2]), .ZN(n4) );
endmodule


module MUX81_26 ( A, B, C, D, E, F, G, H, S, Y );
  input [2:0] S;
  input A, B, C, D, E, F, G, H;
  output Y;
  wire   n1, n2, n3, n4, n5, n6, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35;

  NAND3_X1 U20 ( .A1(S[1]), .A2(n21), .A3(H), .ZN(n23) );
  NAND3_X1 U21 ( .A1(S[0]), .A2(n2), .A3(F), .ZN(n25) );
  INV_X1 U1 ( .A(n27), .ZN(n6) );
  NAND2_X1 U2 ( .A1(G), .A2(n22), .ZN(n24) );
  NOR2_X1 U3 ( .A1(n1), .A2(n3), .ZN(n27) );
  NAND4_X1 U4 ( .A1(A), .A2(n1), .A3(n2), .A4(n4), .ZN(n34) );
  INV_X1 U5 ( .A(n22), .ZN(n21) );
  AOI22_X1 U6 ( .A1(n33), .A2(n5), .B1(B), .B2(n32), .ZN(n35) );
  INV_X1 U7 ( .A(n32), .ZN(n5) );
  NOR3_X1 U8 ( .A1(S[1]), .A2(n3), .A3(n1), .ZN(n32) );
  OAI21_X1 U9 ( .B1(n31), .B2(n30), .A(n29), .ZN(n33) );
  NAND2_X1 U10 ( .A1(C), .A2(n30), .ZN(n29) );
  AOI22_X1 U11 ( .A1(n28), .A2(n6), .B1(D), .B2(n27), .ZN(n31) );
  NOR3_X1 U12 ( .A1(S[0]), .A2(n3), .A3(n2), .ZN(n30) );
  NAND4_X1 U13 ( .A1(n26), .A2(n25), .A3(n24), .A4(n23), .ZN(n28) );
  NAND4_X1 U14 ( .A1(E), .A2(n3), .A3(n1), .A4(n2), .ZN(n26) );
  NAND2_X1 U15 ( .A1(n35), .A2(n34), .ZN(Y) );
  NOR2_X1 U16 ( .A1(n2), .A2(S[0]), .ZN(n22) );
  INV_X1 U17 ( .A(S[0]), .ZN(n1) );
  INV_X1 U18 ( .A(S[1]), .ZN(n2) );
  INV_X1 U19 ( .A(n4), .ZN(n3) );
  INV_X1 U22 ( .A(S[2]), .ZN(n4) );
endmodule


module MUX81_25 ( A, B, C, D, E, F, G, H, S, Y );
  input [2:0] S;
  input A, B, C, D, E, F, G, H;
  output Y;
  wire   n1, n2, n3, n4, n5, n6, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35;

  NAND3_X1 U20 ( .A1(S[1]), .A2(n21), .A3(H), .ZN(n23) );
  NAND3_X1 U21 ( .A1(S[0]), .A2(n2), .A3(F), .ZN(n25) );
  INV_X1 U1 ( .A(n27), .ZN(n6) );
  NOR2_X1 U2 ( .A1(n1), .A2(n3), .ZN(n27) );
  NAND4_X1 U3 ( .A1(A), .A2(n1), .A3(n2), .A4(n4), .ZN(n34) );
  INV_X1 U4 ( .A(n22), .ZN(n21) );
  AOI22_X1 U5 ( .A1(n33), .A2(n5), .B1(B), .B2(n32), .ZN(n35) );
  INV_X1 U6 ( .A(n32), .ZN(n5) );
  NOR3_X1 U7 ( .A1(S[1]), .A2(n3), .A3(n1), .ZN(n32) );
  OAI21_X1 U8 ( .B1(n31), .B2(n30), .A(n29), .ZN(n33) );
  NAND2_X1 U9 ( .A1(C), .A2(n30), .ZN(n29) );
  AOI22_X1 U10 ( .A1(n28), .A2(n6), .B1(D), .B2(n27), .ZN(n31) );
  NOR3_X1 U11 ( .A1(S[0]), .A2(n3), .A3(n2), .ZN(n30) );
  NAND4_X1 U12 ( .A1(n26), .A2(n25), .A3(n24), .A4(n23), .ZN(n28) );
  NAND4_X1 U13 ( .A1(E), .A2(n3), .A3(n1), .A4(n2), .ZN(n26) );
  NAND2_X1 U14 ( .A1(G), .A2(n22), .ZN(n24) );
  NAND2_X1 U15 ( .A1(n35), .A2(n34), .ZN(Y) );
  NOR2_X1 U16 ( .A1(n2), .A2(S[0]), .ZN(n22) );
  INV_X1 U17 ( .A(S[0]), .ZN(n1) );
  INV_X1 U18 ( .A(S[1]), .ZN(n2) );
  INV_X1 U19 ( .A(n4), .ZN(n3) );
  INV_X1 U22 ( .A(S[2]), .ZN(n4) );
endmodule


module MUX81_24 ( A, B, C, D, E, F, G, H, S, Y );
  input [2:0] S;
  input A, B, C, D, E, F, G, H;
  output Y;
  wire   n1, n2, n3, n4, n5, n6, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35;

  NAND3_X1 U20 ( .A1(S[1]), .A2(n21), .A3(H), .ZN(n23) );
  NAND3_X1 U21 ( .A1(S[0]), .A2(n2), .A3(F), .ZN(n25) );
  INV_X1 U1 ( .A(n27), .ZN(n6) );
  NOR2_X1 U2 ( .A1(n1), .A2(n3), .ZN(n27) );
  NAND4_X1 U3 ( .A1(A), .A2(n1), .A3(n2), .A4(n4), .ZN(n34) );
  INV_X1 U4 ( .A(n22), .ZN(n21) );
  AOI22_X1 U5 ( .A1(n33), .A2(n5), .B1(B), .B2(n32), .ZN(n35) );
  INV_X1 U6 ( .A(n32), .ZN(n5) );
  NOR3_X1 U7 ( .A1(S[1]), .A2(n3), .A3(n1), .ZN(n32) );
  OAI21_X1 U8 ( .B1(n31), .B2(n30), .A(n29), .ZN(n33) );
  NAND2_X1 U9 ( .A1(C), .A2(n30), .ZN(n29) );
  AOI22_X1 U10 ( .A1(n28), .A2(n6), .B1(D), .B2(n27), .ZN(n31) );
  NOR3_X1 U11 ( .A1(S[0]), .A2(n3), .A3(n2), .ZN(n30) );
  NAND4_X1 U12 ( .A1(n26), .A2(n25), .A3(n24), .A4(n23), .ZN(n28) );
  NAND4_X1 U13 ( .A1(E), .A2(n3), .A3(n1), .A4(n2), .ZN(n26) );
  NAND2_X1 U14 ( .A1(G), .A2(n22), .ZN(n24) );
  NOR2_X1 U15 ( .A1(n2), .A2(S[0]), .ZN(n22) );
  NAND2_X1 U16 ( .A1(n35), .A2(n34), .ZN(Y) );
  INV_X1 U17 ( .A(S[0]), .ZN(n1) );
  INV_X1 U18 ( .A(S[1]), .ZN(n2) );
  INV_X1 U19 ( .A(n4), .ZN(n3) );
  INV_X1 U22 ( .A(S[2]), .ZN(n4) );
endmodule


module MUX81_23 ( A, B, C, D, E, F, G, H, S, Y );
  input [2:0] S;
  input A, B, C, D, E, F, G, H;
  output Y;
  wire   n1, n2, n3, n4, n5, n6, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34;

  NAND3_X1 U20 ( .A1(S[1]), .A2(n6), .A3(H), .ZN(n22) );
  NAND3_X1 U21 ( .A1(S[0]), .A2(n2), .A3(F), .ZN(n24) );
  INV_X1 U1 ( .A(n26), .ZN(n5) );
  NAND2_X1 U2 ( .A1(G), .A2(n21), .ZN(n23) );
  NOR2_X1 U3 ( .A1(n1), .A2(S[2]), .ZN(n26) );
  NAND4_X1 U4 ( .A1(A), .A2(n1), .A3(n2), .A4(n3), .ZN(n33) );
  INV_X1 U5 ( .A(n21), .ZN(n6) );
  AOI22_X1 U6 ( .A1(n32), .A2(n4), .B1(B), .B2(n31), .ZN(n34) );
  INV_X1 U7 ( .A(n31), .ZN(n4) );
  NOR3_X1 U8 ( .A1(S[1]), .A2(S[2]), .A3(n1), .ZN(n31) );
  OAI21_X1 U9 ( .B1(n30), .B2(n29), .A(n28), .ZN(n32) );
  NAND2_X1 U10 ( .A1(C), .A2(n29), .ZN(n28) );
  AOI22_X1 U11 ( .A1(n27), .A2(n5), .B1(D), .B2(n26), .ZN(n30) );
  NOR3_X1 U12 ( .A1(S[0]), .A2(S[2]), .A3(n2), .ZN(n29) );
  NAND4_X1 U13 ( .A1(n25), .A2(n24), .A3(n23), .A4(n22), .ZN(n27) );
  NAND4_X1 U14 ( .A1(E), .A2(S[2]), .A3(n1), .A4(n2), .ZN(n25) );
  NAND2_X1 U15 ( .A1(n34), .A2(n33), .ZN(Y) );
  NOR2_X1 U16 ( .A1(n2), .A2(S[0]), .ZN(n21) );
  INV_X1 U17 ( .A(S[0]), .ZN(n1) );
  INV_X1 U18 ( .A(S[1]), .ZN(n2) );
  INV_X1 U19 ( .A(S[2]), .ZN(n3) );
endmodule


module MUX81_22 ( A, B, C, D, E, F, G, H, S, Y );
  input [2:0] S;
  input A, B, C, D, E, F, G, H;
  output Y;
  wire   n1, n2, n3, n4, n5, n6, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34;

  NAND3_X1 U20 ( .A1(S[1]), .A2(n6), .A3(H), .ZN(n22) );
  NAND3_X1 U21 ( .A1(S[0]), .A2(n2), .A3(F), .ZN(n24) );
  INV_X1 U1 ( .A(n26), .ZN(n5) );
  NAND2_X1 U2 ( .A1(G), .A2(n21), .ZN(n23) );
  NOR2_X1 U3 ( .A1(n1), .A2(S[2]), .ZN(n26) );
  NAND4_X1 U4 ( .A1(A), .A2(n1), .A3(n2), .A4(n3), .ZN(n33) );
  INV_X1 U5 ( .A(n21), .ZN(n6) );
  NAND2_X1 U6 ( .A1(n34), .A2(n33), .ZN(Y) );
  AOI22_X1 U7 ( .A1(n32), .A2(n4), .B1(B), .B2(n31), .ZN(n34) );
  INV_X1 U8 ( .A(n31), .ZN(n4) );
  NOR3_X1 U9 ( .A1(S[1]), .A2(S[2]), .A3(n1), .ZN(n31) );
  OAI21_X1 U10 ( .B1(n30), .B2(n29), .A(n28), .ZN(n32) );
  NAND2_X1 U11 ( .A1(C), .A2(n29), .ZN(n28) );
  AOI22_X1 U12 ( .A1(n27), .A2(n5), .B1(D), .B2(n26), .ZN(n30) );
  NOR3_X1 U13 ( .A1(S[0]), .A2(S[2]), .A3(n2), .ZN(n29) );
  NAND4_X1 U14 ( .A1(n25), .A2(n24), .A3(n23), .A4(n22), .ZN(n27) );
  NAND4_X1 U15 ( .A1(E), .A2(S[2]), .A3(n1), .A4(n2), .ZN(n25) );
  NOR2_X1 U16 ( .A1(n2), .A2(S[0]), .ZN(n21) );
  INV_X1 U17 ( .A(S[0]), .ZN(n1) );
  INV_X1 U18 ( .A(S[1]), .ZN(n2) );
  INV_X1 U19 ( .A(S[2]), .ZN(n3) );
endmodule


module MUX81_21 ( A, B, C, D, E, F, G, H, S, Y );
  input [2:0] S;
  input A, B, C, D, E, F, G, H;
  output Y;
  wire   n1, n2, n3, n4, n5, n6, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34;

  NAND3_X1 U20 ( .A1(S[1]), .A2(n6), .A3(H), .ZN(n22) );
  NAND3_X1 U21 ( .A1(S[0]), .A2(n2), .A3(F), .ZN(n24) );
  INV_X1 U1 ( .A(n26), .ZN(n5) );
  NOR2_X1 U2 ( .A1(n1), .A2(S[2]), .ZN(n26) );
  NAND4_X1 U3 ( .A1(A), .A2(n1), .A3(n2), .A4(n3), .ZN(n33) );
  NAND2_X1 U4 ( .A1(n34), .A2(n33), .ZN(Y) );
  INV_X1 U5 ( .A(n21), .ZN(n6) );
  AOI22_X1 U6 ( .A1(n32), .A2(n4), .B1(B), .B2(n31), .ZN(n34) );
  INV_X1 U7 ( .A(n31), .ZN(n4) );
  NOR3_X1 U8 ( .A1(S[1]), .A2(S[2]), .A3(n1), .ZN(n31) );
  OAI21_X1 U9 ( .B1(n30), .B2(n29), .A(n28), .ZN(n32) );
  NAND2_X1 U10 ( .A1(C), .A2(n29), .ZN(n28) );
  AOI22_X1 U11 ( .A1(n27), .A2(n5), .B1(D), .B2(n26), .ZN(n30) );
  NOR3_X1 U12 ( .A1(S[0]), .A2(S[2]), .A3(n2), .ZN(n29) );
  NAND4_X1 U13 ( .A1(n25), .A2(n24), .A3(n23), .A4(n22), .ZN(n27) );
  NAND4_X1 U14 ( .A1(E), .A2(S[2]), .A3(n1), .A4(n2), .ZN(n25) );
  NAND2_X1 U15 ( .A1(G), .A2(n21), .ZN(n23) );
  NOR2_X1 U16 ( .A1(n2), .A2(S[0]), .ZN(n21) );
  INV_X1 U17 ( .A(S[0]), .ZN(n1) );
  INV_X1 U18 ( .A(S[1]), .ZN(n2) );
  INV_X1 U19 ( .A(S[2]), .ZN(n3) );
endmodule


module MUX81_20 ( A, B, C, D, E, F, G, H, S, Y );
  input [2:0] S;
  input A, B, C, D, E, F, G, H;
  output Y;
  wire   n1, n2, n3, n4, n5, n6, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35;

  NAND3_X1 U20 ( .A1(S[1]), .A2(n21), .A3(H), .ZN(n23) );
  NAND3_X1 U21 ( .A1(S[0]), .A2(n2), .A3(F), .ZN(n25) );
  INV_X1 U1 ( .A(n27), .ZN(n6) );
  NOR2_X1 U2 ( .A1(n1), .A2(n3), .ZN(n27) );
  NAND4_X1 U3 ( .A1(A), .A2(n1), .A3(n2), .A4(n4), .ZN(n34) );
  INV_X1 U4 ( .A(n22), .ZN(n21) );
  AOI22_X1 U5 ( .A1(n33), .A2(n5), .B1(B), .B2(n32), .ZN(n35) );
  INV_X1 U6 ( .A(n32), .ZN(n5) );
  NOR3_X1 U7 ( .A1(S[1]), .A2(n3), .A3(n1), .ZN(n32) );
  OAI21_X1 U8 ( .B1(n31), .B2(n30), .A(n29), .ZN(n33) );
  NAND2_X1 U9 ( .A1(C), .A2(n30), .ZN(n29) );
  AOI22_X1 U10 ( .A1(n28), .A2(n6), .B1(D), .B2(n27), .ZN(n31) );
  NOR3_X1 U11 ( .A1(S[0]), .A2(n3), .A3(n2), .ZN(n30) );
  NAND4_X1 U12 ( .A1(n26), .A2(n25), .A3(n24), .A4(n23), .ZN(n28) );
  NAND4_X1 U13 ( .A1(E), .A2(n3), .A3(n1), .A4(n2), .ZN(n26) );
  NAND2_X1 U14 ( .A1(G), .A2(n22), .ZN(n24) );
  NOR2_X1 U15 ( .A1(n2), .A2(S[0]), .ZN(n22) );
  NAND2_X1 U16 ( .A1(n35), .A2(n34), .ZN(Y) );
  INV_X1 U17 ( .A(S[0]), .ZN(n1) );
  INV_X1 U18 ( .A(S[1]), .ZN(n2) );
  INV_X1 U19 ( .A(n4), .ZN(n3) );
  INV_X1 U22 ( .A(S[2]), .ZN(n4) );
endmodule


module MUX81_19 ( A, B, C, D, E, F, G, H, S, Y );
  input [2:0] S;
  input A, B, C, D, E, F, G, H;
  output Y;
  wire   n1, n2, n3, n4, n5, n6, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35;

  NAND3_X1 U20 ( .A1(S[1]), .A2(n21), .A3(H), .ZN(n23) );
  NAND3_X1 U21 ( .A1(S[0]), .A2(n2), .A3(F), .ZN(n25) );
  INV_X1 U1 ( .A(n27), .ZN(n6) );
  NOR2_X1 U2 ( .A1(n1), .A2(n3), .ZN(n27) );
  NAND4_X1 U3 ( .A1(A), .A2(n1), .A3(n2), .A4(n4), .ZN(n34) );
  NAND2_X1 U4 ( .A1(n35), .A2(n34), .ZN(Y) );
  INV_X1 U5 ( .A(n22), .ZN(n21) );
  AOI22_X1 U6 ( .A1(n33), .A2(n5), .B1(B), .B2(n32), .ZN(n35) );
  INV_X1 U7 ( .A(n32), .ZN(n5) );
  NOR3_X1 U8 ( .A1(S[1]), .A2(n3), .A3(n1), .ZN(n32) );
  OAI21_X1 U9 ( .B1(n31), .B2(n30), .A(n29), .ZN(n33) );
  NAND2_X1 U10 ( .A1(C), .A2(n30), .ZN(n29) );
  AOI22_X1 U11 ( .A1(n28), .A2(n6), .B1(D), .B2(n27), .ZN(n31) );
  NOR3_X1 U12 ( .A1(S[0]), .A2(n3), .A3(n2), .ZN(n30) );
  NAND4_X1 U13 ( .A1(n26), .A2(n25), .A3(n24), .A4(n23), .ZN(n28) );
  NAND4_X1 U14 ( .A1(E), .A2(n3), .A3(n1), .A4(n2), .ZN(n26) );
  NAND2_X1 U15 ( .A1(G), .A2(n22), .ZN(n24) );
  NOR2_X1 U16 ( .A1(n2), .A2(S[0]), .ZN(n22) );
  INV_X1 U17 ( .A(S[0]), .ZN(n1) );
  INV_X1 U18 ( .A(S[1]), .ZN(n2) );
  INV_X1 U19 ( .A(n4), .ZN(n3) );
  INV_X1 U22 ( .A(S[2]), .ZN(n4) );
endmodule


module MUX81_18 ( A, B, C, D, E, F, G, H, S, Y );
  input [2:0] S;
  input A, B, C, D, E, F, G, H;
  output Y;
  wire   n1, n2, n3, n4, n5, n6, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35;

  NAND3_X1 U20 ( .A1(S[1]), .A2(n21), .A3(H), .ZN(n23) );
  NAND3_X1 U21 ( .A1(S[0]), .A2(n2), .A3(F), .ZN(n25) );
  INV_X1 U1 ( .A(n27), .ZN(n6) );
  NOR2_X1 U2 ( .A1(n1), .A2(n3), .ZN(n27) );
  NAND4_X1 U3 ( .A1(A), .A2(n1), .A3(n2), .A4(n4), .ZN(n34) );
  NAND2_X1 U4 ( .A1(n35), .A2(n34), .ZN(Y) );
  INV_X1 U5 ( .A(n22), .ZN(n21) );
  AOI22_X1 U6 ( .A1(n33), .A2(n5), .B1(B), .B2(n32), .ZN(n35) );
  INV_X1 U7 ( .A(n32), .ZN(n5) );
  NOR3_X1 U8 ( .A1(S[1]), .A2(n3), .A3(n1), .ZN(n32) );
  OAI21_X1 U9 ( .B1(n31), .B2(n30), .A(n29), .ZN(n33) );
  NAND2_X1 U10 ( .A1(C), .A2(n30), .ZN(n29) );
  AOI22_X1 U11 ( .A1(n28), .A2(n6), .B1(D), .B2(n27), .ZN(n31) );
  NOR3_X1 U12 ( .A1(S[0]), .A2(n3), .A3(n2), .ZN(n30) );
  NAND4_X1 U13 ( .A1(n26), .A2(n25), .A3(n24), .A4(n23), .ZN(n28) );
  NAND4_X1 U14 ( .A1(E), .A2(n3), .A3(n1), .A4(n2), .ZN(n26) );
  NAND2_X1 U15 ( .A1(G), .A2(n22), .ZN(n24) );
  NOR2_X1 U16 ( .A1(n2), .A2(S[0]), .ZN(n22) );
  INV_X1 U17 ( .A(S[0]), .ZN(n1) );
  INV_X1 U18 ( .A(S[1]), .ZN(n2) );
  INV_X1 U19 ( .A(n4), .ZN(n3) );
  INV_X1 U22 ( .A(S[2]), .ZN(n4) );
endmodule


module MUX81_17 ( A, B, C, D, E, F, G, H, S, Y );
  input [2:0] S;
  input A, B, C, D, E, F, G, H;
  output Y;
  wire   n1, n2, n3, n4, n5, n6, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35;

  NAND3_X1 U20 ( .A1(S[1]), .A2(n21), .A3(H), .ZN(n23) );
  NAND3_X1 U21 ( .A1(S[0]), .A2(n2), .A3(F), .ZN(n25) );
  INV_X1 U1 ( .A(n27), .ZN(n6) );
  NOR2_X1 U2 ( .A1(n1), .A2(n3), .ZN(n27) );
  NAND4_X1 U3 ( .A1(A), .A2(n1), .A3(n2), .A4(n4), .ZN(n34) );
  NAND2_X1 U4 ( .A1(n35), .A2(n34), .ZN(Y) );
  INV_X1 U5 ( .A(n22), .ZN(n21) );
  AOI22_X1 U6 ( .A1(n33), .A2(n5), .B1(B), .B2(n32), .ZN(n35) );
  INV_X1 U7 ( .A(n32), .ZN(n5) );
  NOR3_X1 U8 ( .A1(S[1]), .A2(n3), .A3(n1), .ZN(n32) );
  OAI21_X1 U9 ( .B1(n31), .B2(n30), .A(n29), .ZN(n33) );
  NAND2_X1 U10 ( .A1(C), .A2(n30), .ZN(n29) );
  AOI22_X1 U11 ( .A1(n28), .A2(n6), .B1(D), .B2(n27), .ZN(n31) );
  NOR3_X1 U12 ( .A1(S[0]), .A2(n3), .A3(n2), .ZN(n30) );
  NAND4_X1 U13 ( .A1(n26), .A2(n25), .A3(n24), .A4(n23), .ZN(n28) );
  NAND4_X1 U14 ( .A1(E), .A2(n3), .A3(n1), .A4(n2), .ZN(n26) );
  NAND2_X1 U15 ( .A1(G), .A2(n22), .ZN(n24) );
  NOR2_X1 U16 ( .A1(n2), .A2(S[0]), .ZN(n22) );
  INV_X1 U17 ( .A(S[0]), .ZN(n1) );
  INV_X1 U18 ( .A(S[1]), .ZN(n2) );
  INV_X1 U19 ( .A(n4), .ZN(n3) );
  INV_X1 U22 ( .A(S[2]), .ZN(n4) );
endmodule


module MUX81_16 ( A, B, C, D, E, F, G, H, S, Y );
  input [2:0] S;
  input A, B, C, D, E, F, G, H;
  output Y;
  wire   n1, n2, n3, n4, n5, n6, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35;

  NAND3_X1 U20 ( .A1(S[1]), .A2(n21), .A3(H), .ZN(n23) );
  NAND3_X1 U21 ( .A1(S[0]), .A2(n2), .A3(F), .ZN(n25) );
  INV_X1 U1 ( .A(n27), .ZN(n6) );
  NOR2_X1 U2 ( .A1(n1), .A2(n3), .ZN(n27) );
  NAND4_X1 U3 ( .A1(A), .A2(n1), .A3(n2), .A4(n4), .ZN(n34) );
  INV_X1 U4 ( .A(n22), .ZN(n21) );
  AOI22_X1 U5 ( .A1(n33), .A2(n5), .B1(B), .B2(n32), .ZN(n35) );
  INV_X1 U6 ( .A(n32), .ZN(n5) );
  NOR3_X1 U7 ( .A1(S[1]), .A2(n3), .A3(n1), .ZN(n32) );
  OAI21_X1 U8 ( .B1(n31), .B2(n30), .A(n29), .ZN(n33) );
  NAND2_X1 U9 ( .A1(C), .A2(n30), .ZN(n29) );
  AOI22_X1 U10 ( .A1(n28), .A2(n6), .B1(D), .B2(n27), .ZN(n31) );
  NOR3_X1 U11 ( .A1(S[0]), .A2(n3), .A3(n2), .ZN(n30) );
  NAND4_X1 U12 ( .A1(n26), .A2(n25), .A3(n24), .A4(n23), .ZN(n28) );
  NAND4_X1 U13 ( .A1(E), .A2(n3), .A3(n1), .A4(n2), .ZN(n26) );
  NAND2_X1 U14 ( .A1(G), .A2(n22), .ZN(n24) );
  NOR2_X1 U15 ( .A1(n2), .A2(S[0]), .ZN(n22) );
  NAND2_X1 U16 ( .A1(n35), .A2(n34), .ZN(Y) );
  INV_X1 U17 ( .A(S[0]), .ZN(n1) );
  INV_X1 U18 ( .A(S[1]), .ZN(n2) );
  INV_X1 U19 ( .A(n4), .ZN(n3) );
  INV_X1 U22 ( .A(S[2]), .ZN(n4) );
endmodule


module MUX81_15 ( A, B, C, D, E, F, G, H, S, Y );
  input [2:0] S;
  input A, B, C, D, E, F, G, H;
  output Y;
  wire   n1, n2, n3, n4, n5, n6, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35;

  NAND3_X1 U20 ( .A1(S[1]), .A2(n21), .A3(H), .ZN(n23) );
  NAND3_X1 U21 ( .A1(S[0]), .A2(n2), .A3(F), .ZN(n25) );
  INV_X1 U1 ( .A(n27), .ZN(n6) );
  NOR2_X1 U2 ( .A1(n1), .A2(n3), .ZN(n27) );
  NAND4_X1 U3 ( .A1(A), .A2(n1), .A3(n2), .A4(n4), .ZN(n34) );
  INV_X1 U4 ( .A(n22), .ZN(n21) );
  AOI22_X1 U5 ( .A1(n33), .A2(n5), .B1(B), .B2(n32), .ZN(n35) );
  INV_X1 U6 ( .A(n32), .ZN(n5) );
  NOR3_X1 U7 ( .A1(S[1]), .A2(n3), .A3(n1), .ZN(n32) );
  OAI21_X1 U8 ( .B1(n31), .B2(n30), .A(n29), .ZN(n33) );
  NAND2_X1 U9 ( .A1(C), .A2(n30), .ZN(n29) );
  AOI22_X1 U10 ( .A1(n28), .A2(n6), .B1(D), .B2(n27), .ZN(n31) );
  NOR3_X1 U11 ( .A1(S[0]), .A2(n3), .A3(n2), .ZN(n30) );
  NAND4_X1 U12 ( .A1(n26), .A2(n25), .A3(n24), .A4(n23), .ZN(n28) );
  NAND4_X1 U13 ( .A1(E), .A2(n3), .A3(n1), .A4(n2), .ZN(n26) );
  NAND2_X1 U14 ( .A1(G), .A2(n22), .ZN(n24) );
  NAND2_X1 U15 ( .A1(n35), .A2(n34), .ZN(Y) );
  NOR2_X1 U16 ( .A1(n2), .A2(S[0]), .ZN(n22) );
  INV_X1 U17 ( .A(S[0]), .ZN(n1) );
  INV_X1 U18 ( .A(S[1]), .ZN(n2) );
  INV_X1 U19 ( .A(n4), .ZN(n3) );
  INV_X1 U22 ( .A(S[2]), .ZN(n4) );
endmodule


module MUX81_14 ( A, B, C, D, E, F, G, H, S, Y );
  input [2:0] S;
  input A, B, C, D, E, F, G, H;
  output Y;
  wire   n1, n2, n3, n4, n5, n6, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35;

  NAND3_X1 U20 ( .A1(S[1]), .A2(n21), .A3(H), .ZN(n23) );
  NAND3_X1 U21 ( .A1(S[0]), .A2(n2), .A3(F), .ZN(n25) );
  INV_X1 U1 ( .A(n27), .ZN(n6) );
  NAND2_X1 U2 ( .A1(G), .A2(n22), .ZN(n24) );
  NOR2_X1 U3 ( .A1(n1), .A2(n3), .ZN(n27) );
  NAND4_X1 U4 ( .A1(A), .A2(n1), .A3(n2), .A4(n4), .ZN(n34) );
  INV_X1 U5 ( .A(n22), .ZN(n21) );
  AOI22_X1 U6 ( .A1(n33), .A2(n5), .B1(B), .B2(n32), .ZN(n35) );
  INV_X1 U7 ( .A(n32), .ZN(n5) );
  NOR3_X1 U8 ( .A1(S[1]), .A2(n3), .A3(n1), .ZN(n32) );
  OAI21_X1 U9 ( .B1(n31), .B2(n30), .A(n29), .ZN(n33) );
  NAND2_X1 U10 ( .A1(C), .A2(n30), .ZN(n29) );
  AOI22_X1 U11 ( .A1(n28), .A2(n6), .B1(D), .B2(n27), .ZN(n31) );
  NOR3_X1 U12 ( .A1(S[0]), .A2(n3), .A3(n2), .ZN(n30) );
  NAND4_X1 U13 ( .A1(n26), .A2(n25), .A3(n24), .A4(n23), .ZN(n28) );
  NAND4_X1 U14 ( .A1(E), .A2(n3), .A3(n1), .A4(n2), .ZN(n26) );
  NAND2_X1 U15 ( .A1(n35), .A2(n34), .ZN(Y) );
  NOR2_X1 U16 ( .A1(n2), .A2(S[0]), .ZN(n22) );
  INV_X1 U17 ( .A(S[0]), .ZN(n1) );
  INV_X1 U18 ( .A(S[1]), .ZN(n2) );
  INV_X1 U19 ( .A(n4), .ZN(n3) );
  INV_X1 U22 ( .A(S[2]), .ZN(n4) );
endmodule


module MUX81_13 ( A, B, C, D, E, F, G, H, S, Y );
  input [2:0] S;
  input A, B, C, D, E, F, G, H;
  output Y;
  wire   n1, n2, n3, n4, n5, n6, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35;

  NAND3_X1 U20 ( .A1(S[1]), .A2(n21), .A3(H), .ZN(n23) );
  NAND3_X1 U21 ( .A1(S[0]), .A2(n2), .A3(F), .ZN(n25) );
  INV_X1 U1 ( .A(n27), .ZN(n6) );
  NAND2_X1 U2 ( .A1(G), .A2(n22), .ZN(n24) );
  NOR2_X1 U3 ( .A1(n1), .A2(n3), .ZN(n27) );
  NAND4_X1 U4 ( .A1(A), .A2(n1), .A3(n2), .A4(n4), .ZN(n34) );
  INV_X1 U5 ( .A(n22), .ZN(n21) );
  NAND2_X1 U6 ( .A1(n35), .A2(n34), .ZN(Y) );
  AOI22_X1 U7 ( .A1(n33), .A2(n5), .B1(B), .B2(n32), .ZN(n35) );
  INV_X1 U8 ( .A(n32), .ZN(n5) );
  NOR3_X1 U9 ( .A1(S[1]), .A2(n3), .A3(n1), .ZN(n32) );
  OAI21_X1 U10 ( .B1(n31), .B2(n30), .A(n29), .ZN(n33) );
  NAND2_X1 U11 ( .A1(C), .A2(n30), .ZN(n29) );
  AOI22_X1 U12 ( .A1(n28), .A2(n6), .B1(D), .B2(n27), .ZN(n31) );
  NOR3_X1 U13 ( .A1(S[0]), .A2(n3), .A3(n2), .ZN(n30) );
  NAND4_X1 U14 ( .A1(n26), .A2(n25), .A3(n24), .A4(n23), .ZN(n28) );
  NAND4_X1 U15 ( .A1(E), .A2(n3), .A3(n1), .A4(n2), .ZN(n26) );
  NOR2_X1 U16 ( .A1(n2), .A2(S[0]), .ZN(n22) );
  INV_X1 U17 ( .A(S[0]), .ZN(n1) );
  INV_X1 U18 ( .A(S[1]), .ZN(n2) );
  INV_X1 U19 ( .A(n4), .ZN(n3) );
  INV_X1 U22 ( .A(S[2]), .ZN(n4) );
endmodule


module MUX81_12 ( A, B, C, D, E, F, G, H, S, Y );
  input [2:0] S;
  input A, B, C, D, E, F, G, H;
  output Y;
  wire   n1, n2, n3, n4, n5, n6, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34;

  NAND3_X1 U20 ( .A1(S[1]), .A2(n6), .A3(H), .ZN(n22) );
  NAND3_X1 U21 ( .A1(S[0]), .A2(n2), .A3(F), .ZN(n24) );
  INV_X1 U1 ( .A(n26), .ZN(n5) );
  NAND2_X1 U2 ( .A1(G), .A2(n21), .ZN(n23) );
  NOR2_X1 U3 ( .A1(n1), .A2(S[2]), .ZN(n26) );
  NAND4_X1 U4 ( .A1(A), .A2(n1), .A3(n2), .A4(n3), .ZN(n33) );
  INV_X1 U5 ( .A(n21), .ZN(n6) );
  AOI22_X1 U6 ( .A1(n32), .A2(n4), .B1(B), .B2(n31), .ZN(n34) );
  INV_X1 U7 ( .A(n31), .ZN(n4) );
  NOR3_X1 U8 ( .A1(S[1]), .A2(S[2]), .A3(n1), .ZN(n31) );
  OAI21_X1 U9 ( .B1(n30), .B2(n29), .A(n28), .ZN(n32) );
  NAND2_X1 U10 ( .A1(C), .A2(n29), .ZN(n28) );
  AOI22_X1 U11 ( .A1(n27), .A2(n5), .B1(D), .B2(n26), .ZN(n30) );
  NOR3_X1 U12 ( .A1(S[0]), .A2(S[2]), .A3(n2), .ZN(n29) );
  NAND4_X1 U13 ( .A1(n25), .A2(n24), .A3(n23), .A4(n22), .ZN(n27) );
  NAND4_X1 U14 ( .A1(E), .A2(S[2]), .A3(n1), .A4(n2), .ZN(n25) );
  NOR2_X1 U15 ( .A1(n2), .A2(S[0]), .ZN(n21) );
  NAND2_X1 U16 ( .A1(n34), .A2(n33), .ZN(Y) );
  INV_X1 U17 ( .A(S[0]), .ZN(n1) );
  INV_X1 U18 ( .A(S[1]), .ZN(n2) );
  INV_X1 U19 ( .A(S[2]), .ZN(n3) );
endmodule


module MUX81_11 ( A, B, C, D, E, F, G, H, S, Y );
  input [2:0] S;
  input A, B, C, D, E, F, G, H;
  output Y;
  wire   n1, n2, n3, n4, n5, n6, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34;

  NAND3_X1 U20 ( .A1(S[1]), .A2(n6), .A3(H), .ZN(n22) );
  NAND3_X1 U21 ( .A1(S[0]), .A2(n2), .A3(F), .ZN(n24) );
  INV_X1 U1 ( .A(n26), .ZN(n5) );
  NAND2_X1 U2 ( .A1(G), .A2(n21), .ZN(n23) );
  NOR2_X1 U3 ( .A1(n1), .A2(S[2]), .ZN(n26) );
  NAND4_X1 U4 ( .A1(A), .A2(n1), .A3(n2), .A4(n3), .ZN(n33) );
  INV_X1 U5 ( .A(n21), .ZN(n6) );
  NAND2_X1 U6 ( .A1(n34), .A2(n33), .ZN(Y) );
  AOI22_X1 U7 ( .A1(n32), .A2(n4), .B1(B), .B2(n31), .ZN(n34) );
  INV_X1 U8 ( .A(n31), .ZN(n4) );
  NOR3_X1 U9 ( .A1(S[1]), .A2(S[2]), .A3(n1), .ZN(n31) );
  OAI21_X1 U10 ( .B1(n30), .B2(n29), .A(n28), .ZN(n32) );
  NAND2_X1 U11 ( .A1(C), .A2(n29), .ZN(n28) );
  AOI22_X1 U12 ( .A1(n27), .A2(n5), .B1(D), .B2(n26), .ZN(n30) );
  NOR3_X1 U13 ( .A1(S[0]), .A2(S[2]), .A3(n2), .ZN(n29) );
  NAND4_X1 U14 ( .A1(n25), .A2(n24), .A3(n23), .A4(n22), .ZN(n27) );
  NAND4_X1 U15 ( .A1(E), .A2(S[2]), .A3(n1), .A4(n2), .ZN(n25) );
  NOR2_X1 U16 ( .A1(n2), .A2(S[0]), .ZN(n21) );
  INV_X1 U17 ( .A(S[0]), .ZN(n1) );
  INV_X1 U18 ( .A(S[1]), .ZN(n2) );
  INV_X1 U19 ( .A(S[2]), .ZN(n3) );
endmodule


module MUX81_10 ( A, B, C, D, E, F, G, H, S, Y );
  input [2:0] S;
  input A, B, C, D, E, F, G, H;
  output Y;
  wire   n1, n2, n3, n4, n5, n6, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34;

  NAND3_X1 U20 ( .A1(S[1]), .A2(n6), .A3(H), .ZN(n22) );
  NAND3_X1 U21 ( .A1(S[0]), .A2(n2), .A3(F), .ZN(n24) );
  INV_X1 U1 ( .A(n26), .ZN(n5) );
  NAND2_X1 U2 ( .A1(G), .A2(n21), .ZN(n23) );
  NOR2_X1 U3 ( .A1(n1), .A2(S[2]), .ZN(n26) );
  NAND4_X1 U4 ( .A1(A), .A2(n1), .A3(n2), .A4(n3), .ZN(n33) );
  INV_X1 U5 ( .A(n21), .ZN(n6) );
  NAND2_X1 U6 ( .A1(n34), .A2(n33), .ZN(Y) );
  AOI22_X1 U7 ( .A1(n32), .A2(n4), .B1(B), .B2(n31), .ZN(n34) );
  INV_X1 U8 ( .A(n31), .ZN(n4) );
  NOR3_X1 U9 ( .A1(S[1]), .A2(S[2]), .A3(n1), .ZN(n31) );
  OAI21_X1 U10 ( .B1(n30), .B2(n29), .A(n28), .ZN(n32) );
  NAND2_X1 U11 ( .A1(C), .A2(n29), .ZN(n28) );
  AOI22_X1 U12 ( .A1(n27), .A2(n5), .B1(D), .B2(n26), .ZN(n30) );
  NOR3_X1 U13 ( .A1(S[0]), .A2(S[2]), .A3(n2), .ZN(n29) );
  NAND4_X1 U14 ( .A1(n25), .A2(n24), .A3(n23), .A4(n22), .ZN(n27) );
  NAND4_X1 U15 ( .A1(E), .A2(S[2]), .A3(n1), .A4(n2), .ZN(n25) );
  NOR2_X1 U16 ( .A1(n2), .A2(S[0]), .ZN(n21) );
  INV_X1 U17 ( .A(S[0]), .ZN(n1) );
  INV_X1 U18 ( .A(S[1]), .ZN(n2) );
  INV_X1 U19 ( .A(S[2]), .ZN(n3) );
endmodule


module MUX81_9 ( A, B, C, D, E, F, G, H, S, Y );
  input [2:0] S;
  input A, B, C, D, E, F, G, H;
  output Y;
  wire   n1, n2, n3, n4, n5, n6, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35;

  NAND3_X1 U20 ( .A1(S[1]), .A2(n21), .A3(H), .ZN(n23) );
  NAND3_X1 U21 ( .A1(S[0]), .A2(n2), .A3(F), .ZN(n25) );
  INV_X1 U1 ( .A(n27), .ZN(n6) );
  NOR2_X1 U2 ( .A1(n1), .A2(n3), .ZN(n27) );
  NAND4_X1 U3 ( .A1(A), .A2(n1), .A3(n2), .A4(n4), .ZN(n34) );
  INV_X1 U4 ( .A(n22), .ZN(n21) );
  AOI22_X1 U5 ( .A1(n33), .A2(n5), .B1(B), .B2(n32), .ZN(n35) );
  INV_X1 U6 ( .A(n32), .ZN(n5) );
  NOR3_X1 U7 ( .A1(S[1]), .A2(n3), .A3(n1), .ZN(n32) );
  OAI21_X1 U8 ( .B1(n31), .B2(n30), .A(n29), .ZN(n33) );
  NAND2_X1 U9 ( .A1(C), .A2(n30), .ZN(n29) );
  AOI22_X1 U10 ( .A1(n28), .A2(n6), .B1(D), .B2(n27), .ZN(n31) );
  NOR3_X1 U11 ( .A1(S[0]), .A2(n3), .A3(n2), .ZN(n30) );
  NAND4_X1 U12 ( .A1(n26), .A2(n25), .A3(n24), .A4(n23), .ZN(n28) );
  NAND4_X1 U13 ( .A1(E), .A2(n3), .A3(n1), .A4(n2), .ZN(n26) );
  NAND2_X1 U14 ( .A1(G), .A2(n22), .ZN(n24) );
  NAND2_X1 U15 ( .A1(n35), .A2(n34), .ZN(Y) );
  NOR2_X1 U16 ( .A1(n2), .A2(S[0]), .ZN(n22) );
  INV_X1 U17 ( .A(S[0]), .ZN(n1) );
  INV_X1 U18 ( .A(S[1]), .ZN(n2) );
  INV_X1 U19 ( .A(n4), .ZN(n3) );
  INV_X1 U22 ( .A(S[2]), .ZN(n4) );
endmodule


module MUX81_8 ( A, B, C, D, E, F, G, H, S, Y );
  input [2:0] S;
  input A, B, C, D, E, F, G, H;
  output Y;
  wire   n1, n2, n3, n4, n5, n6, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35;

  NAND3_X1 U20 ( .A1(S[1]), .A2(n21), .A3(H), .ZN(n23) );
  NAND3_X1 U21 ( .A1(S[0]), .A2(n2), .A3(F), .ZN(n25) );
  INV_X1 U1 ( .A(n27), .ZN(n6) );
  NOR2_X1 U2 ( .A1(n1), .A2(n3), .ZN(n27) );
  NAND4_X1 U3 ( .A1(A), .A2(n1), .A3(n2), .A4(n4), .ZN(n34) );
  INV_X1 U4 ( .A(n22), .ZN(n21) );
  AOI22_X1 U5 ( .A1(n33), .A2(n5), .B1(B), .B2(n32), .ZN(n35) );
  INV_X1 U6 ( .A(n32), .ZN(n5) );
  NOR3_X1 U7 ( .A1(S[1]), .A2(n3), .A3(n1), .ZN(n32) );
  OAI21_X1 U8 ( .B1(n31), .B2(n30), .A(n29), .ZN(n33) );
  NAND2_X1 U9 ( .A1(C), .A2(n30), .ZN(n29) );
  AOI22_X1 U10 ( .A1(n28), .A2(n6), .B1(D), .B2(n27), .ZN(n31) );
  NOR3_X1 U11 ( .A1(S[0]), .A2(n3), .A3(n2), .ZN(n30) );
  NAND4_X1 U12 ( .A1(n26), .A2(n25), .A3(n24), .A4(n23), .ZN(n28) );
  NAND4_X1 U13 ( .A1(E), .A2(n3), .A3(n1), .A4(n2), .ZN(n26) );
  NAND2_X1 U14 ( .A1(G), .A2(n22), .ZN(n24) );
  NOR2_X1 U15 ( .A1(n2), .A2(S[0]), .ZN(n22) );
  NAND2_X1 U16 ( .A1(n35), .A2(n34), .ZN(Y) );
  INV_X1 U17 ( .A(S[0]), .ZN(n1) );
  INV_X1 U18 ( .A(S[1]), .ZN(n2) );
  INV_X1 U19 ( .A(n4), .ZN(n3) );
  INV_X1 U22 ( .A(S[2]), .ZN(n4) );
endmodule


module MUX81_7 ( A, B, C, D, E, F, G, H, S, Y );
  input [2:0] S;
  input A, B, C, D, E, F, G, H;
  output Y;
  wire   n1, n2, n3, n4, n5, n6, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35;

  NAND3_X1 U20 ( .A1(S[1]), .A2(n21), .A3(H), .ZN(n23) );
  NAND3_X1 U21 ( .A1(S[0]), .A2(n2), .A3(F), .ZN(n25) );
  INV_X1 U1 ( .A(n27), .ZN(n6) );
  NAND2_X1 U2 ( .A1(G), .A2(n22), .ZN(n24) );
  NOR2_X1 U3 ( .A1(n1), .A2(n3), .ZN(n27) );
  NAND4_X1 U4 ( .A1(A), .A2(n1), .A3(n2), .A4(n4), .ZN(n34) );
  INV_X1 U5 ( .A(n22), .ZN(n21) );
  AOI22_X1 U6 ( .A1(n33), .A2(n5), .B1(B), .B2(n32), .ZN(n35) );
  INV_X1 U7 ( .A(n32), .ZN(n5) );
  NOR3_X1 U8 ( .A1(S[1]), .A2(n3), .A3(n1), .ZN(n32) );
  OAI21_X1 U9 ( .B1(n31), .B2(n30), .A(n29), .ZN(n33) );
  NAND2_X1 U10 ( .A1(C), .A2(n30), .ZN(n29) );
  AOI22_X1 U11 ( .A1(n28), .A2(n6), .B1(D), .B2(n27), .ZN(n31) );
  NOR3_X1 U12 ( .A1(S[0]), .A2(n3), .A3(n2), .ZN(n30) );
  NAND4_X1 U13 ( .A1(n26), .A2(n25), .A3(n24), .A4(n23), .ZN(n28) );
  NAND4_X1 U14 ( .A1(E), .A2(n3), .A3(n1), .A4(n2), .ZN(n26) );
  NAND2_X1 U15 ( .A1(n35), .A2(n34), .ZN(Y) );
  NOR2_X1 U16 ( .A1(n2), .A2(S[0]), .ZN(n22) );
  INV_X1 U17 ( .A(S[0]), .ZN(n1) );
  INV_X1 U18 ( .A(S[1]), .ZN(n2) );
  INV_X1 U19 ( .A(n4), .ZN(n3) );
  INV_X1 U22 ( .A(S[2]), .ZN(n4) );
endmodule


module MUX81_6 ( A, B, C, D, E, F, G, H, S, Y );
  input [2:0] S;
  input A, B, C, D, E, F, G, H;
  output Y;
  wire   n1, n2, n3, n4, n5, n6, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35;

  NAND3_X1 U20 ( .A1(S[1]), .A2(n21), .A3(H), .ZN(n23) );
  NAND3_X1 U21 ( .A1(S[0]), .A2(n2), .A3(F), .ZN(n25) );
  INV_X1 U1 ( .A(n27), .ZN(n6) );
  NOR2_X1 U2 ( .A1(n1), .A2(n3), .ZN(n27) );
  NAND4_X1 U3 ( .A1(A), .A2(n1), .A3(n2), .A4(n4), .ZN(n34) );
  INV_X1 U4 ( .A(n22), .ZN(n21) );
  AOI22_X1 U5 ( .A1(n33), .A2(n5), .B1(B), .B2(n32), .ZN(n35) );
  INV_X1 U6 ( .A(n32), .ZN(n5) );
  NOR3_X1 U7 ( .A1(S[1]), .A2(n3), .A3(n1), .ZN(n32) );
  OAI21_X1 U8 ( .B1(n31), .B2(n30), .A(n29), .ZN(n33) );
  NAND2_X1 U9 ( .A1(C), .A2(n30), .ZN(n29) );
  AOI22_X1 U10 ( .A1(n28), .A2(n6), .B1(D), .B2(n27), .ZN(n31) );
  NOR3_X1 U11 ( .A1(S[0]), .A2(n3), .A3(n2), .ZN(n30) );
  NAND4_X1 U12 ( .A1(n26), .A2(n25), .A3(n24), .A4(n23), .ZN(n28) );
  NAND4_X1 U13 ( .A1(E), .A2(n3), .A3(n1), .A4(n2), .ZN(n26) );
  NAND2_X1 U14 ( .A1(G), .A2(n22), .ZN(n24) );
  NAND2_X1 U15 ( .A1(n35), .A2(n34), .ZN(Y) );
  NOR2_X1 U16 ( .A1(n2), .A2(S[0]), .ZN(n22) );
  INV_X1 U17 ( .A(S[0]), .ZN(n1) );
  INV_X1 U18 ( .A(S[1]), .ZN(n2) );
  INV_X1 U19 ( .A(n4), .ZN(n3) );
  INV_X1 U22 ( .A(S[2]), .ZN(n4) );
endmodule


module MUX81_5 ( A, B, C, D, E, F, G, H, S, Y );
  input [2:0] S;
  input A, B, C, D, E, F, G, H;
  output Y;
  wire   n1, n2, n3, n4, n5, n6, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35;

  NAND3_X1 U20 ( .A1(S[1]), .A2(n21), .A3(H), .ZN(n23) );
  NAND3_X1 U21 ( .A1(S[0]), .A2(n2), .A3(F), .ZN(n25) );
  INV_X1 U1 ( .A(n27), .ZN(n6) );
  NOR2_X1 U2 ( .A1(n1), .A2(n3), .ZN(n27) );
  NAND4_X1 U3 ( .A1(A), .A2(n1), .A3(n2), .A4(n4), .ZN(n34) );
  INV_X1 U4 ( .A(n22), .ZN(n21) );
  AOI22_X1 U5 ( .A1(n33), .A2(n5), .B1(B), .B2(n32), .ZN(n35) );
  INV_X1 U6 ( .A(n32), .ZN(n5) );
  NOR3_X1 U7 ( .A1(S[1]), .A2(n3), .A3(n1), .ZN(n32) );
  OAI21_X1 U8 ( .B1(n31), .B2(n30), .A(n29), .ZN(n33) );
  NAND2_X1 U9 ( .A1(C), .A2(n30), .ZN(n29) );
  AOI22_X1 U10 ( .A1(n28), .A2(n6), .B1(D), .B2(n27), .ZN(n31) );
  NOR3_X1 U11 ( .A1(S[0]), .A2(n3), .A3(n2), .ZN(n30) );
  NAND4_X1 U12 ( .A1(n26), .A2(n25), .A3(n24), .A4(n23), .ZN(n28) );
  NAND4_X1 U13 ( .A1(E), .A2(n3), .A3(n1), .A4(n2), .ZN(n26) );
  NAND2_X1 U14 ( .A1(G), .A2(n22), .ZN(n24) );
  NAND2_X1 U15 ( .A1(n35), .A2(n34), .ZN(Y) );
  NOR2_X1 U16 ( .A1(n2), .A2(S[0]), .ZN(n22) );
  INV_X1 U17 ( .A(S[0]), .ZN(n1) );
  INV_X1 U18 ( .A(S[1]), .ZN(n2) );
  INV_X1 U19 ( .A(n4), .ZN(n3) );
  INV_X1 U22 ( .A(S[2]), .ZN(n4) );
endmodule


module MUX81_4 ( A, B, C, D, E, F, G, H, S, Y );
  input [2:0] S;
  input A, B, C, D, E, F, G, H;
  output Y;
  wire   n1, n2, n3, n4, n5, n6, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35;

  NAND3_X1 U20 ( .A1(S[1]), .A2(n21), .A3(H), .ZN(n23) );
  NAND3_X1 U21 ( .A1(S[0]), .A2(n2), .A3(F), .ZN(n25) );
  INV_X1 U1 ( .A(n27), .ZN(n6) );
  NOR2_X1 U2 ( .A1(n1), .A2(n3), .ZN(n27) );
  NAND4_X1 U3 ( .A1(A), .A2(n1), .A3(n2), .A4(n4), .ZN(n34) );
  INV_X1 U4 ( .A(n22), .ZN(n21) );
  AOI22_X1 U5 ( .A1(n33), .A2(n5), .B1(B), .B2(n32), .ZN(n35) );
  INV_X1 U6 ( .A(n32), .ZN(n5) );
  NOR3_X1 U7 ( .A1(S[1]), .A2(n3), .A3(n1), .ZN(n32) );
  OAI21_X1 U8 ( .B1(n31), .B2(n30), .A(n29), .ZN(n33) );
  NAND2_X1 U9 ( .A1(C), .A2(n30), .ZN(n29) );
  AOI22_X1 U10 ( .A1(n28), .A2(n6), .B1(D), .B2(n27), .ZN(n31) );
  NOR3_X1 U11 ( .A1(S[0]), .A2(n3), .A3(n2), .ZN(n30) );
  NAND4_X1 U12 ( .A1(n26), .A2(n25), .A3(n24), .A4(n23), .ZN(n28) );
  NAND4_X1 U13 ( .A1(E), .A2(n3), .A3(n1), .A4(n2), .ZN(n26) );
  NAND2_X1 U14 ( .A1(G), .A2(n22), .ZN(n24) );
  NOR2_X1 U15 ( .A1(n2), .A2(S[0]), .ZN(n22) );
  NAND2_X1 U16 ( .A1(n35), .A2(n34), .ZN(Y) );
  INV_X1 U17 ( .A(S[0]), .ZN(n1) );
  INV_X1 U18 ( .A(S[1]), .ZN(n2) );
  INV_X1 U19 ( .A(n4), .ZN(n3) );
  INV_X1 U22 ( .A(S[2]), .ZN(n4) );
endmodule


module MUX81_3 ( A, B, C, D, E, F, G, H, S, Y );
  input [2:0] S;
  input A, B, C, D, E, F, G, H;
  output Y;
  wire   n1, n2, n3, n4, n5, n6, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35;

  NAND3_X1 U20 ( .A1(S[1]), .A2(n21), .A3(H), .ZN(n23) );
  NAND3_X1 U21 ( .A1(S[0]), .A2(n2), .A3(F), .ZN(n25) );
  INV_X1 U1 ( .A(n27), .ZN(n6) );
  NOR2_X1 U2 ( .A1(n1), .A2(n3), .ZN(n27) );
  NAND4_X1 U3 ( .A1(A), .A2(n1), .A3(n2), .A4(n4), .ZN(n34) );
  INV_X1 U4 ( .A(n22), .ZN(n21) );
  AOI22_X1 U5 ( .A1(n33), .A2(n5), .B1(B), .B2(n32), .ZN(n35) );
  INV_X1 U6 ( .A(n32), .ZN(n5) );
  NOR3_X1 U7 ( .A1(S[1]), .A2(n3), .A3(n1), .ZN(n32) );
  OAI21_X1 U8 ( .B1(n31), .B2(n30), .A(n29), .ZN(n33) );
  NAND2_X1 U9 ( .A1(C), .A2(n30), .ZN(n29) );
  AOI22_X1 U10 ( .A1(n28), .A2(n6), .B1(D), .B2(n27), .ZN(n31) );
  NOR3_X1 U11 ( .A1(S[0]), .A2(n3), .A3(n2), .ZN(n30) );
  NAND4_X1 U12 ( .A1(n26), .A2(n25), .A3(n24), .A4(n23), .ZN(n28) );
  NAND4_X1 U13 ( .A1(E), .A2(n3), .A3(n1), .A4(n2), .ZN(n26) );
  NAND2_X1 U14 ( .A1(G), .A2(n22), .ZN(n24) );
  NAND2_X1 U15 ( .A1(n35), .A2(n34), .ZN(Y) );
  NOR2_X1 U16 ( .A1(n2), .A2(S[0]), .ZN(n22) );
  INV_X1 U17 ( .A(S[0]), .ZN(n1) );
  INV_X1 U18 ( .A(S[1]), .ZN(n2) );
  INV_X1 U19 ( .A(n4), .ZN(n3) );
  INV_X1 U22 ( .A(S[2]), .ZN(n4) );
endmodule


module MUX81_2 ( A, B, C, D, E, F, G, H, S, Y );
  input [2:0] S;
  input A, B, C, D, E, F, G, H;
  output Y;
  wire   n1, n2, n3, n4, n5, n6, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34;

  NAND3_X1 U20 ( .A1(S[1]), .A2(n6), .A3(H), .ZN(n22) );
  NAND3_X1 U21 ( .A1(S[0]), .A2(n2), .A3(F), .ZN(n24) );
  INV_X1 U1 ( .A(n26), .ZN(n5) );
  NOR2_X1 U2 ( .A1(n1), .A2(S[2]), .ZN(n26) );
  NAND4_X1 U3 ( .A1(A), .A2(n1), .A3(n2), .A4(n3), .ZN(n33) );
  INV_X1 U4 ( .A(n21), .ZN(n6) );
  AOI22_X1 U5 ( .A1(n32), .A2(n4), .B1(B), .B2(n31), .ZN(n34) );
  INV_X1 U6 ( .A(n31), .ZN(n4) );
  NOR3_X1 U7 ( .A1(S[1]), .A2(S[2]), .A3(n1), .ZN(n31) );
  OAI21_X1 U8 ( .B1(n30), .B2(n29), .A(n28), .ZN(n32) );
  NAND2_X1 U9 ( .A1(C), .A2(n29), .ZN(n28) );
  AOI22_X1 U10 ( .A1(n27), .A2(n5), .B1(D), .B2(n26), .ZN(n30) );
  NOR3_X1 U11 ( .A1(S[0]), .A2(S[2]), .A3(n2), .ZN(n29) );
  NAND4_X1 U12 ( .A1(n25), .A2(n24), .A3(n23), .A4(n22), .ZN(n27) );
  NAND4_X1 U13 ( .A1(E), .A2(S[2]), .A3(n1), .A4(n2), .ZN(n25) );
  NAND2_X1 U14 ( .A1(G), .A2(n21), .ZN(n23) );
  NAND2_X1 U15 ( .A1(n34), .A2(n33), .ZN(Y) );
  NOR2_X1 U16 ( .A1(n2), .A2(S[0]), .ZN(n21) );
  INV_X1 U17 ( .A(S[0]), .ZN(n1) );
  INV_X1 U18 ( .A(S[1]), .ZN(n2) );
  INV_X1 U19 ( .A(S[2]), .ZN(n3) );
endmodule


module MUX81_1 ( A, B, C, D, E, F, G, H, S, Y );
  input [2:0] S;
  input A, B, C, D, E, F, G, H;
  output Y;
  wire   n1, n2, n3, n4, n5, n6, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34;

  NAND3_X1 U20 ( .A1(S[1]), .A2(n6), .A3(H), .ZN(n22) );
  NAND3_X1 U21 ( .A1(S[0]), .A2(n2), .A3(F), .ZN(n24) );
  INV_X1 U1 ( .A(n26), .ZN(n5) );
  NOR2_X1 U2 ( .A1(n1), .A2(S[2]), .ZN(n26) );
  NAND4_X1 U3 ( .A1(A), .A2(n1), .A3(n2), .A4(n3), .ZN(n33) );
  INV_X1 U4 ( .A(n21), .ZN(n6) );
  AOI22_X1 U5 ( .A1(n32), .A2(n4), .B1(B), .B2(n31), .ZN(n34) );
  INV_X1 U6 ( .A(n31), .ZN(n4) );
  NOR3_X1 U7 ( .A1(S[1]), .A2(S[2]), .A3(n1), .ZN(n31) );
  OAI21_X1 U8 ( .B1(n30), .B2(n29), .A(n28), .ZN(n32) );
  NAND2_X1 U9 ( .A1(C), .A2(n29), .ZN(n28) );
  AOI22_X1 U10 ( .A1(n27), .A2(n5), .B1(D), .B2(n26), .ZN(n30) );
  NOR3_X1 U11 ( .A1(S[0]), .A2(S[2]), .A3(n2), .ZN(n29) );
  NAND4_X1 U12 ( .A1(n25), .A2(n24), .A3(n23), .A4(n22), .ZN(n27) );
  NAND4_X1 U13 ( .A1(E), .A2(S[2]), .A3(n1), .A4(n2), .ZN(n25) );
  NAND2_X1 U14 ( .A1(G), .A2(n21), .ZN(n23) );
  NAND2_X1 U15 ( .A1(n34), .A2(n33), .ZN(Y) );
  NOR2_X1 U16 ( .A1(n2), .A2(S[0]), .ZN(n21) );
  INV_X1 U17 ( .A(S[0]), .ZN(n1) );
  INV_X1 U18 ( .A(S[1]), .ZN(n2) );
  INV_X1 U19 ( .A(S[2]), .ZN(n3) );
endmodule


module MUX81_GENERIC_NBIT32 ( A, B, C, D, E, F, G, H, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [31:0] D;
  input [31:0] E;
  input [31:0] F;
  input [31:0] G;
  input [31:0] H;
  input [2:0] SEL;
  output [31:0] Y;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9;

  MUX81_0 MUXES_0 ( .A(A[0]), .B(B[0]), .C(C[0]), .D(D[0]), .E(E[0]), .F(F[0]), 
        .G(G[0]), .H(H[0]), .S({n9, n6, n3}), .Y(Y[0]) );
  MUX81_31 MUXES_1 ( .A(A[1]), .B(B[1]), .C(C[1]), .D(D[1]), .E(E[1]), .F(F[1]), .G(G[1]), .H(H[1]), .S({n7, n4, n1}), .Y(Y[1]) );
  MUX81_30 MUXES_2 ( .A(A[2]), .B(B[2]), .C(C[2]), .D(D[2]), .E(E[2]), .F(F[2]), .G(G[2]), .H(H[2]), .S({n7, n4, n1}), .Y(Y[2]) );
  MUX81_29 MUXES_3 ( .A(A[3]), .B(B[3]), .C(C[3]), .D(D[3]), .E(E[3]), .F(F[3]), .G(G[3]), .H(H[3]), .S({n7, n4, n1}), .Y(Y[3]) );
  MUX81_28 MUXES_4 ( .A(A[4]), .B(B[4]), .C(C[4]), .D(D[4]), .E(E[4]), .F(F[4]), .G(G[4]), .H(H[4]), .S({n7, n4, n1}), .Y(Y[4]) );
  MUX81_27 MUXES_5 ( .A(A[5]), .B(B[5]), .C(C[5]), .D(D[5]), .E(E[5]), .F(F[5]), .G(G[5]), .H(H[5]), .S({n7, n4, n1}), .Y(Y[5]) );
  MUX81_26 MUXES_6 ( .A(A[6]), .B(B[6]), .C(C[6]), .D(D[6]), .E(E[6]), .F(F[6]), .G(G[6]), .H(H[6]), .S({n7, n4, n1}), .Y(Y[6]) );
  MUX81_25 MUXES_7 ( .A(A[7]), .B(B[7]), .C(C[7]), .D(D[7]), .E(E[7]), .F(F[7]), .G(G[7]), .H(H[7]), .S({n7, n4, n1}), .Y(Y[7]) );
  MUX81_24 MUXES_8 ( .A(A[8]), .B(B[8]), .C(C[8]), .D(D[8]), .E(E[8]), .F(F[8]), .G(G[8]), .H(H[8]), .S({n7, n4, n1}), .Y(Y[8]) );
  MUX81_23 MUXES_9 ( .A(A[9]), .B(B[9]), .C(C[9]), .D(D[9]), .E(E[9]), .F(F[9]), .G(G[9]), .H(H[9]), .S({n7, n4, n1}), .Y(Y[9]) );
  MUX81_22 MUXES_10 ( .A(A[10]), .B(B[10]), .C(C[10]), .D(D[10]), .E(E[10]), 
        .F(F[10]), .G(G[10]), .H(H[10]), .S({n7, n4, n1}), .Y(Y[10]) );
  MUX81_21 MUXES_11 ( .A(A[11]), .B(B[11]), .C(C[11]), .D(D[11]), .E(E[11]), 
        .F(F[11]), .G(G[11]), .H(H[11]), .S({n7, n4, n1}), .Y(Y[11]) );
  MUX81_20 MUXES_12 ( .A(A[12]), .B(B[12]), .C(C[12]), .D(D[12]), .E(E[12]), 
        .F(F[12]), .G(G[12]), .H(H[12]), .S({n8, n4, n1}), .Y(Y[12]) );
  MUX81_19 MUXES_13 ( .A(A[13]), .B(B[13]), .C(C[13]), .D(D[13]), .E(E[13]), 
        .F(F[13]), .G(G[13]), .H(H[13]), .S({n8, n5, n2}), .Y(Y[13]) );
  MUX81_18 MUXES_14 ( .A(A[14]), .B(B[14]), .C(C[14]), .D(D[14]), .E(E[14]), 
        .F(F[14]), .G(G[14]), .H(H[14]), .S({n8, n5, n2}), .Y(Y[14]) );
  MUX81_17 MUXES_15 ( .A(A[15]), .B(B[15]), .C(C[15]), .D(D[15]), .E(E[15]), 
        .F(F[15]), .G(G[15]), .H(H[15]), .S({n8, n5, n2}), .Y(Y[15]) );
  MUX81_16 MUXES_16 ( .A(A[16]), .B(B[16]), .C(C[16]), .D(D[16]), .E(E[16]), 
        .F(F[16]), .G(G[16]), .H(H[16]), .S({n8, n5, n2}), .Y(Y[16]) );
  MUX81_15 MUXES_17 ( .A(A[17]), .B(B[17]), .C(C[17]), .D(D[17]), .E(E[17]), 
        .F(F[17]), .G(G[17]), .H(H[17]), .S({n8, n5, n2}), .Y(Y[17]) );
  MUX81_14 MUXES_18 ( .A(A[18]), .B(B[18]), .C(C[18]), .D(D[18]), .E(E[18]), 
        .F(F[18]), .G(G[18]), .H(H[18]), .S({n8, n5, n2}), .Y(Y[18]) );
  MUX81_13 MUXES_19 ( .A(A[19]), .B(B[19]), .C(C[19]), .D(D[19]), .E(E[19]), 
        .F(F[19]), .G(G[19]), .H(H[19]), .S({n8, n5, n2}), .Y(Y[19]) );
  MUX81_12 MUXES_20 ( .A(A[20]), .B(B[20]), .C(C[20]), .D(D[20]), .E(E[20]), 
        .F(F[20]), .G(G[20]), .H(H[20]), .S({n8, n5, n2}), .Y(Y[20]) );
  MUX81_11 MUXES_21 ( .A(A[21]), .B(B[21]), .C(C[21]), .D(D[21]), .E(E[21]), 
        .F(F[21]), .G(G[21]), .H(H[21]), .S({n8, n5, n2}), .Y(Y[21]) );
  MUX81_10 MUXES_22 ( .A(A[22]), .B(B[22]), .C(C[22]), .D(D[22]), .E(E[22]), 
        .F(F[22]), .G(G[22]), .H(H[22]), .S({n8, n5, n2}), .Y(Y[22]) );
  MUX81_9 MUXES_23 ( .A(A[23]), .B(B[23]), .C(C[23]), .D(D[23]), .E(E[23]), 
        .F(F[23]), .G(G[23]), .H(H[23]), .S({n9, n5, n2}), .Y(Y[23]) );
  MUX81_8 MUXES_24 ( .A(A[24]), .B(B[24]), .C(C[24]), .D(D[24]), .E(E[24]), 
        .F(F[24]), .G(G[24]), .H(H[24]), .S({n9, n5, n2}), .Y(Y[24]) );
  MUX81_7 MUXES_25 ( .A(A[25]), .B(B[25]), .C(C[25]), .D(D[25]), .E(E[25]), 
        .F(F[25]), .G(G[25]), .H(H[25]), .S({n9, n6, n3}), .Y(Y[25]) );
  MUX81_6 MUXES_26 ( .A(A[26]), .B(B[26]), .C(C[26]), .D(D[26]), .E(E[26]), 
        .F(F[26]), .G(G[26]), .H(H[26]), .S({n9, n6, n3}), .Y(Y[26]) );
  MUX81_5 MUXES_27 ( .A(A[27]), .B(B[27]), .C(C[27]), .D(D[27]), .E(E[27]), 
        .F(F[27]), .G(G[27]), .H(H[27]), .S({n9, n6, n3}), .Y(Y[27]) );
  MUX81_4 MUXES_28 ( .A(A[28]), .B(B[28]), .C(C[28]), .D(D[28]), .E(E[28]), 
        .F(F[28]), .G(G[28]), .H(H[28]), .S({n9, n6, n3}), .Y(Y[28]) );
  MUX81_3 MUXES_29 ( .A(A[29]), .B(B[29]), .C(C[29]), .D(D[29]), .E(E[29]), 
        .F(F[29]), .G(G[29]), .H(H[29]), .S({n9, n6, n3}), .Y(Y[29]) );
  MUX81_2 MUXES_30 ( .A(A[30]), .B(B[30]), .C(C[30]), .D(D[30]), .E(E[30]), 
        .F(F[30]), .G(G[30]), .H(H[30]), .S({n9, n6, n3}), .Y(Y[30]) );
  MUX81_1 MUXES_31 ( .A(A[31]), .B(B[31]), .C(C[31]), .D(D[31]), .E(E[31]), 
        .F(F[31]), .G(G[31]), .H(H[31]), .S({n9, n6, n3}), .Y(Y[31]) );
  BUF_X2 U1 ( .A(SEL[0]), .Z(n2) );
  BUF_X2 U2 ( .A(SEL[0]), .Z(n1) );
  BUF_X1 U3 ( .A(SEL[1]), .Z(n6) );
  BUF_X2 U4 ( .A(SEL[0]), .Z(n3) );
  BUF_X2 U5 ( .A(SEL[1]), .Z(n5) );
  BUF_X2 U6 ( .A(SEL[1]), .Z(n4) );
  BUF_X1 U7 ( .A(SEL[2]), .Z(n8) );
  BUF_X1 U8 ( .A(SEL[2]), .Z(n7) );
  BUF_X1 U9 ( .A(SEL[2]), .Z(n9) );
endmodule


module shifter_NBITS32 ( R1, R2, LnR, AnL, RnS, Rout );
  input [31:0] R1;
  input [31:0] R2;
  output [31:0] Rout;
  input LnR, AnL, RnS;
  wire   s_RnS, n1;
  wire   [39:0] s_mask0;
  wire   [39:0] s_mask8;
  wire   [39:0] s_mask16;
  wire   [39:0] s_mask24;
  wire   [39:0] s_selected_mask;
  wire   [31:0] s_sh0;
  wire   [31:0] s_sh1;
  wire   [31:0] s_sh2;
  wire   [31:0] s_sh3;
  wire   [31:0] s_sh4;
  wire   [31:0] s_sh5;
  wire   [31:0] s_sh6;
  wire   [31:0] s_sh7;

  mask_generator_NBITS32 mask_gen ( .R1(R1), .R2(R2), .LnR(LnR), .AnL(AnL), 
        .RnS(s_RnS), .mask0(s_mask0), .mask8(s_mask8), .mask16(s_mask16), 
        .mask24(s_mask24) );
  MUX41_GENERIC_NBIT40 MUX_mask_select ( .A(s_mask0), .B(s_mask8), .C(s_mask16), .D(s_mask24), .SEL(R2[4:3]), .Y(s_selected_mask) );
  mask_shifter_NBITS40 mask_shift ( .R1(s_selected_mask), .LnR(LnR), 
        .mask_sh0(s_sh0), .mask_sh1(s_sh1), .mask_sh2(s_sh2), .mask_sh3(s_sh3), 
        .mask_sh4(s_sh4), .mask_sh5(s_sh5), .mask_sh6(s_sh6), .mask_sh7(s_sh7)
         );
  MUX81_GENERIC_NBIT32 MUX_shift_select ( .A(s_sh0), .B(s_sh1), .C(s_sh2), .D(
        s_sh3), .E(s_sh4), .F(s_sh5), .G(s_sh6), .H(s_sh7), .SEL(R2[2:0]), .Y(
        Rout) );
  NOR2_X1 U1 ( .A1(LnR), .A2(n1), .ZN(s_RnS) );
  INV_X1 U2 ( .A(RnS), .ZN(n1) );
endmodule


module my_xor_224 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_223 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_222 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_221 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_220 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_219 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_218 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_217 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_216 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_215 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_214 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_213 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_212 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_211 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_210 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_209 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_208 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_207 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_206 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_205 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_204 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_203 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_202 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_201 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_200 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_199 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_198 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_197 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_196 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_195 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_194 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_193 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module pg_net_220 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_219 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_218 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_217 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_216 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_215 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_214 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_213 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_212 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_211 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_210 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_209 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_208 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_207 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_206 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_205 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_204 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_203 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_202 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_201 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_200 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_199 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_198 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_197 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_196 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_195 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_194 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_193 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_192 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_191 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_190 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_BLOCK_216 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_215 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_214 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_213 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_212 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_211 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_210 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_209 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_208 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_207 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_206 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_205 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_204 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_203 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_202 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_60 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_201 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AOI21_X1 U1 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_200 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_199 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_198 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_197 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_196 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_195 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_59 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_194 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_193 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_192 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_58 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_191 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_190 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_57 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_56 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_55 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_54 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_53 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_52 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_1 ( A, B, Cin, Co );
  input [31:0] A;
  input [31:0] B;
  output [7:0] Co;
  input Cin;
  wire   \g_vector[4][31] , \g_vector[4][27] , \g_vector[3][31] ,
         \g_vector[3][23] , \g_vector[3][15] , \g_vector[2][31] ,
         \g_vector[2][27] , \g_vector[2][23] , \g_vector[2][19] ,
         \g_vector[2][15] , \g_vector[2][11] , \g_vector[2][7] ,
         \g_vector[1][31] , \g_vector[1][29] , \g_vector[1][27] ,
         \g_vector[1][25] , \g_vector[1][23] , \g_vector[1][21] ,
         \g_vector[1][19] , \g_vector[1][17] , \g_vector[1][15] ,
         \g_vector[1][13] , \g_vector[1][11] , \g_vector[1][9] ,
         \g_vector[1][7] , \g_vector[1][5] , \g_vector[1][3] ,
         \g_vector[1][1] , \g_vector[0][31] , \g_vector[0][30] ,
         \g_vector[0][29] , \g_vector[0][28] , \g_vector[0][27] ,
         \g_vector[0][26] , \g_vector[0][25] , \g_vector[0][24] ,
         \g_vector[0][23] , \g_vector[0][22] , \g_vector[0][21] ,
         \g_vector[0][20] , \g_vector[0][19] , \g_vector[0][18] ,
         \g_vector[0][17] , \g_vector[0][16] , \g_vector[0][15] ,
         \g_vector[0][14] , \g_vector[0][13] , \g_vector[0][12] ,
         \g_vector[0][11] , \g_vector[0][10] , \g_vector[0][9] ,
         \g_vector[0][8] , \g_vector[0][7] , \g_vector[0][6] ,
         \g_vector[0][5] , \g_vector[0][4] , \g_vector[0][3] ,
         \g_vector[0][2] , \g_vector[0][1] , \g_vector[0][0] ,
         \p_vector[4][31] , \p_vector[4][27] , \p_vector[3][31] ,
         \p_vector[3][23] , \p_vector[3][15] , \p_vector[2][31] ,
         \p_vector[2][27] , \p_vector[2][23] , \p_vector[2][19] ,
         \p_vector[2][15] , \p_vector[2][11] , \p_vector[2][7] ,
         \p_vector[1][31] , \p_vector[1][29] , \p_vector[1][27] ,
         \p_vector[1][25] , \p_vector[1][23] , \p_vector[1][21] ,
         \p_vector[1][19] , \p_vector[1][17] , \p_vector[1][15] ,
         \p_vector[1][13] , \p_vector[1][11] , \p_vector[1][9] ,
         \p_vector[1][7] , \p_vector[1][5] , \p_vector[1][3] ,
         \p_vector[0][31] , \p_vector[0][30] , \p_vector[0][29] ,
         \p_vector[0][28] , \p_vector[0][27] , \p_vector[0][26] ,
         \p_vector[0][25] , \p_vector[0][24] , \p_vector[0][23] ,
         \p_vector[0][22] , \p_vector[0][21] , \p_vector[0][20] ,
         \p_vector[0][19] , \p_vector[0][18] , \p_vector[0][17] ,
         \p_vector[0][16] , \p_vector[0][15] , \p_vector[0][14] ,
         \p_vector[0][13] , \p_vector[0][12] , \p_vector[0][11] ,
         \p_vector[0][10] , \p_vector[0][9] , \p_vector[0][8] ,
         \p_vector[0][7] , \p_vector[0][6] , \p_vector[0][5] ,
         \p_vector[0][4] , \p_vector[0][3] , \p_vector[0][2] ,
         \p_vector[0][1] , n1, n2, n4;

  pg_net_220 pg_network_31 ( .a(A[31]), .b(B[31]), .p(\p_vector[0][31] ), .g(
        \g_vector[0][31] ) );
  pg_net_219 pg_network_30 ( .a(A[30]), .b(B[30]), .p(\p_vector[0][30] ), .g(
        \g_vector[0][30] ) );
  pg_net_218 pg_network_29 ( .a(A[29]), .b(B[29]), .p(\p_vector[0][29] ), .g(
        \g_vector[0][29] ) );
  pg_net_217 pg_network_28 ( .a(A[28]), .b(B[28]), .p(\p_vector[0][28] ), .g(
        \g_vector[0][28] ) );
  pg_net_216 pg_network_27 ( .a(A[27]), .b(B[27]), .p(\p_vector[0][27] ), .g(
        \g_vector[0][27] ) );
  pg_net_215 pg_network_26 ( .a(A[26]), .b(B[26]), .p(\p_vector[0][26] ), .g(
        \g_vector[0][26] ) );
  pg_net_214 pg_network_25 ( .a(A[25]), .b(B[25]), .p(\p_vector[0][25] ), .g(
        \g_vector[0][25] ) );
  pg_net_213 pg_network_24 ( .a(A[24]), .b(B[24]), .p(\p_vector[0][24] ), .g(
        \g_vector[0][24] ) );
  pg_net_212 pg_network_23 ( .a(A[23]), .b(B[23]), .p(\p_vector[0][23] ), .g(
        \g_vector[0][23] ) );
  pg_net_211 pg_network_22 ( .a(A[22]), .b(B[22]), .p(\p_vector[0][22] ), .g(
        \g_vector[0][22] ) );
  pg_net_210 pg_network_21 ( .a(A[21]), .b(B[21]), .p(\p_vector[0][21] ), .g(
        \g_vector[0][21] ) );
  pg_net_209 pg_network_20 ( .a(A[20]), .b(B[20]), .p(\p_vector[0][20] ), .g(
        \g_vector[0][20] ) );
  pg_net_208 pg_network_19 ( .a(A[19]), .b(B[19]), .p(\p_vector[0][19] ), .g(
        \g_vector[0][19] ) );
  pg_net_207 pg_network_18 ( .a(A[18]), .b(B[18]), .p(\p_vector[0][18] ), .g(
        \g_vector[0][18] ) );
  pg_net_206 pg_network_17 ( .a(A[17]), .b(B[17]), .p(\p_vector[0][17] ), .g(
        \g_vector[0][17] ) );
  pg_net_205 pg_network_16 ( .a(A[16]), .b(B[16]), .p(\p_vector[0][16] ), .g(
        \g_vector[0][16] ) );
  pg_net_204 pg_network_15 ( .a(A[15]), .b(B[15]), .p(\p_vector[0][15] ), .g(
        \g_vector[0][15] ) );
  pg_net_203 pg_network_14 ( .a(A[14]), .b(B[14]), .p(\p_vector[0][14] ), .g(
        \g_vector[0][14] ) );
  pg_net_202 pg_network_13 ( .a(A[13]), .b(B[13]), .p(\p_vector[0][13] ), .g(
        \g_vector[0][13] ) );
  pg_net_201 pg_network_12 ( .a(A[12]), .b(B[12]), .p(\p_vector[0][12] ), .g(
        \g_vector[0][12] ) );
  pg_net_200 pg_network_11 ( .a(A[11]), .b(B[11]), .p(\p_vector[0][11] ), .g(
        \g_vector[0][11] ) );
  pg_net_199 pg_network_10 ( .a(A[10]), .b(B[10]), .p(\p_vector[0][10] ), .g(
        \g_vector[0][10] ) );
  pg_net_198 pg_network_9 ( .a(A[9]), .b(B[9]), .p(\p_vector[0][9] ), .g(
        \g_vector[0][9] ) );
  pg_net_197 pg_network_8 ( .a(A[8]), .b(B[8]), .p(\p_vector[0][8] ), .g(
        \g_vector[0][8] ) );
  pg_net_196 pg_network_7 ( .a(A[7]), .b(B[7]), .p(\p_vector[0][7] ), .g(
        \g_vector[0][7] ) );
  pg_net_195 pg_network_6 ( .a(A[6]), .b(B[6]), .p(\p_vector[0][6] ), .g(
        \g_vector[0][6] ) );
  pg_net_194 pg_network_5 ( .a(A[5]), .b(B[5]), .p(\p_vector[0][5] ), .g(
        \g_vector[0][5] ) );
  pg_net_193 pg_network_4 ( .a(A[4]), .b(B[4]), .p(\p_vector[0][4] ), .g(
        \g_vector[0][4] ) );
  pg_net_192 pg_network_3 ( .a(A[3]), .b(B[3]), .p(\p_vector[0][3] ), .g(
        \g_vector[0][3] ) );
  pg_net_191 pg_network_2 ( .a(A[2]), .b(B[2]), .p(\p_vector[0][2] ), .g(
        \g_vector[0][2] ) );
  pg_net_190 pg_network_1 ( .a(A[1]), .b(B[1]), .p(\p_vector[0][1] ), .g(
        \g_vector[0][1] ) );
  PG_BLOCK_216 std_PG_1_31 ( .p2(\p_vector[0][31] ), .g2(\g_vector[0][31] ), 
        .p1(\p_vector[0][30] ), .g1(\g_vector[0][30] ), .PG_P(
        \p_vector[1][31] ), .PG_G(\g_vector[1][31] ) );
  PG_BLOCK_215 std_PG_1_29 ( .p2(\p_vector[0][29] ), .g2(\g_vector[0][29] ), 
        .p1(\p_vector[0][28] ), .g1(\g_vector[0][28] ), .PG_P(
        \p_vector[1][29] ), .PG_G(\g_vector[1][29] ) );
  PG_BLOCK_214 std_PG_1_27 ( .p2(\p_vector[0][27] ), .g2(\g_vector[0][27] ), 
        .p1(\p_vector[0][26] ), .g1(\g_vector[0][26] ), .PG_P(
        \p_vector[1][27] ), .PG_G(\g_vector[1][27] ) );
  PG_BLOCK_213 std_PG_1_25 ( .p2(\p_vector[0][25] ), .g2(\g_vector[0][25] ), 
        .p1(\p_vector[0][24] ), .g1(\g_vector[0][24] ), .PG_P(
        \p_vector[1][25] ), .PG_G(\g_vector[1][25] ) );
  PG_BLOCK_212 std_PG_1_23 ( .p2(\p_vector[0][23] ), .g2(\g_vector[0][23] ), 
        .p1(\p_vector[0][22] ), .g1(\g_vector[0][22] ), .PG_P(
        \p_vector[1][23] ), .PG_G(\g_vector[1][23] ) );
  PG_BLOCK_211 std_PG_1_21 ( .p2(\p_vector[0][21] ), .g2(\g_vector[0][21] ), 
        .p1(\p_vector[0][20] ), .g1(\g_vector[0][20] ), .PG_P(
        \p_vector[1][21] ), .PG_G(\g_vector[1][21] ) );
  PG_BLOCK_210 std_PG_1_19 ( .p2(\p_vector[0][19] ), .g2(\g_vector[0][19] ), 
        .p1(\p_vector[0][18] ), .g1(\g_vector[0][18] ), .PG_P(
        \p_vector[1][19] ), .PG_G(\g_vector[1][19] ) );
  PG_BLOCK_209 std_PG_1_17 ( .p2(\p_vector[0][17] ), .g2(\g_vector[0][17] ), 
        .p1(\p_vector[0][16] ), .g1(\g_vector[0][16] ), .PG_P(
        \p_vector[1][17] ), .PG_G(\g_vector[1][17] ) );
  PG_BLOCK_208 std_PG_1_15 ( .p2(\p_vector[0][15] ), .g2(\g_vector[0][15] ), 
        .p1(\p_vector[0][14] ), .g1(\g_vector[0][14] ), .PG_P(
        \p_vector[1][15] ), .PG_G(\g_vector[1][15] ) );
  PG_BLOCK_207 std_PG_1_13 ( .p2(\p_vector[0][13] ), .g2(\g_vector[0][13] ), 
        .p1(\p_vector[0][12] ), .g1(\g_vector[0][12] ), .PG_P(
        \p_vector[1][13] ), .PG_G(\g_vector[1][13] ) );
  PG_BLOCK_206 std_PG_1_11 ( .p2(\p_vector[0][11] ), .g2(\g_vector[0][11] ), 
        .p1(\p_vector[0][10] ), .g1(\g_vector[0][10] ), .PG_P(
        \p_vector[1][11] ), .PG_G(\g_vector[1][11] ) );
  PG_BLOCK_205 std_PG_1_9 ( .p2(\p_vector[0][9] ), .g2(\g_vector[0][9] ), .p1(
        \p_vector[0][8] ), .g1(\g_vector[0][8] ), .PG_P(\p_vector[1][9] ), 
        .PG_G(\g_vector[1][9] ) );
  PG_BLOCK_204 std_PG_1_7 ( .p2(\p_vector[0][7] ), .g2(\g_vector[0][7] ), .p1(
        \p_vector[0][6] ), .g1(\g_vector[0][6] ), .PG_P(\p_vector[1][7] ), 
        .PG_G(\g_vector[1][7] ) );
  PG_BLOCK_203 std_PG_1_5 ( .p2(\p_vector[0][5] ), .g2(\g_vector[0][5] ), .p1(
        \p_vector[0][4] ), .g1(\g_vector[0][4] ), .PG_P(\p_vector[1][5] ), 
        .PG_G(\g_vector[1][5] ) );
  PG_BLOCK_202 std_PG_1_3 ( .p2(\p_vector[0][3] ), .g2(\g_vector[0][3] ), .p1(
        \p_vector[0][2] ), .g1(\g_vector[0][2] ), .PG_P(\p_vector[1][3] ), 
        .PG_G(\g_vector[1][3] ) );
  G_BLOCK_60 std_G_1_1 ( .p2(\p_vector[0][1] ), .g2(\g_vector[0][1] ), .g1(
        \g_vector[0][0] ), .G(\g_vector[1][1] ) );
  PG_BLOCK_201 std_PG_2_31 ( .p2(\p_vector[1][31] ), .g2(\g_vector[1][31] ), 
        .p1(\p_vector[1][29] ), .g1(\g_vector[1][29] ), .PG_P(
        \p_vector[2][31] ), .PG_G(\g_vector[2][31] ) );
  PG_BLOCK_200 std_PG_2_27 ( .p2(\p_vector[1][27] ), .g2(\g_vector[1][27] ), 
        .p1(\p_vector[1][25] ), .g1(\g_vector[1][25] ), .PG_P(
        \p_vector[2][27] ), .PG_G(\g_vector[2][27] ) );
  PG_BLOCK_199 std_PG_2_23 ( .p2(\p_vector[1][23] ), .g2(\g_vector[1][23] ), 
        .p1(\p_vector[1][21] ), .g1(\g_vector[1][21] ), .PG_P(
        \p_vector[2][23] ), .PG_G(\g_vector[2][23] ) );
  PG_BLOCK_198 std_PG_2_19 ( .p2(\p_vector[1][19] ), .g2(\g_vector[1][19] ), 
        .p1(\p_vector[1][17] ), .g1(\g_vector[1][17] ), .PG_P(
        \p_vector[2][19] ), .PG_G(\g_vector[2][19] ) );
  PG_BLOCK_197 std_PG_2_15 ( .p2(\p_vector[1][15] ), .g2(\g_vector[1][15] ), 
        .p1(\p_vector[1][13] ), .g1(\g_vector[1][13] ), .PG_P(
        \p_vector[2][15] ), .PG_G(\g_vector[2][15] ) );
  PG_BLOCK_196 std_PG_2_11 ( .p2(\p_vector[1][11] ), .g2(\g_vector[1][11] ), 
        .p1(\p_vector[1][9] ), .g1(\g_vector[1][9] ), .PG_P(\p_vector[2][11] ), 
        .PG_G(\g_vector[2][11] ) );
  PG_BLOCK_195 std_PG_2_7 ( .p2(\p_vector[1][7] ), .g2(\g_vector[1][7] ), .p1(
        \p_vector[1][5] ), .g1(\g_vector[1][5] ), .PG_P(\p_vector[2][7] ), 
        .PG_G(\g_vector[2][7] ) );
  G_BLOCK_59 std_G_2_3 ( .p2(\p_vector[1][3] ), .g2(\g_vector[1][3] ), .g1(
        \g_vector[1][1] ), .G(Co[0]) );
  PG_BLOCK_194 std_PG_3_31 ( .p2(\p_vector[2][31] ), .g2(\g_vector[2][31] ), 
        .p1(\p_vector[2][27] ), .g1(\g_vector[2][27] ), .PG_P(
        \p_vector[3][31] ), .PG_G(\g_vector[3][31] ) );
  PG_BLOCK_193 std_PG_3_23 ( .p2(\p_vector[2][23] ), .g2(\g_vector[2][23] ), 
        .p1(\p_vector[2][19] ), .g1(\g_vector[2][19] ), .PG_P(
        \p_vector[3][23] ), .PG_G(\g_vector[3][23] ) );
  PG_BLOCK_192 std_PG_3_15 ( .p2(\p_vector[2][15] ), .g2(\g_vector[2][15] ), 
        .p1(\p_vector[2][11] ), .g1(\g_vector[2][11] ), .PG_P(
        \p_vector[3][15] ), .PG_G(\g_vector[3][15] ) );
  G_BLOCK_58 std_G_3_7 ( .p2(\p_vector[2][7] ), .g2(\g_vector[2][7] ), .g1(
        Co[0]), .G(Co[1]) );
  PG_BLOCK_191 std_PG_4_31 ( .p2(\p_vector[3][31] ), .g2(\g_vector[3][31] ), 
        .p1(\p_vector[3][23] ), .g1(\g_vector[3][23] ), .PG_P(
        \p_vector[4][31] ), .PG_G(\g_vector[4][31] ) );
  PG_BLOCK_190 add_PG_4_31_1 ( .p2(\p_vector[2][27] ), .g2(\g_vector[2][27] ), 
        .p1(\p_vector[3][23] ), .g1(\g_vector[3][23] ), .PG_P(
        \p_vector[4][27] ), .PG_G(\g_vector[4][27] ) );
  G_BLOCK_57 std_G_4_15 ( .p2(\p_vector[3][15] ), .g2(\g_vector[3][15] ), .g1(
        Co[1]), .G(Co[3]) );
  G_BLOCK_56 add_G_4_15_1 ( .p2(\p_vector[2][11] ), .g2(\g_vector[2][11] ), 
        .g1(Co[1]), .G(Co[2]) );
  G_BLOCK_55 std_G_5_31 ( .p2(\p_vector[4][31] ), .g2(\g_vector[4][31] ), .g1(
        Co[3]), .G(Co[7]) );
  G_BLOCK_54 add_G_5_31_1 ( .p2(\p_vector[4][27] ), .g2(\g_vector[4][27] ), 
        .g1(Co[3]), .G(Co[6]) );
  G_BLOCK_53 add_G_5_31_2 ( .p2(\p_vector[3][23] ), .g2(\g_vector[3][23] ), 
        .g1(Co[3]), .G(Co[5]) );
  G_BLOCK_52 add_G_5_31_3 ( .p2(\p_vector[2][19] ), .g2(\g_vector[2][19] ), 
        .g1(Co[3]), .G(Co[4]) );
  OAI21_X1 U1 ( .B1(n2), .B2(n1), .A(n4), .ZN(\g_vector[0][0] ) );
  INV_X1 U2 ( .A(A[0]), .ZN(n2) );
  INV_X1 U3 ( .A(B[0]), .ZN(n1) );
  OAI21_X1 U4 ( .B1(A[0]), .B2(B[0]), .A(Cin), .ZN(n4) );
endmodule


module FA_448 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_447 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_446 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_445 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_112 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_448 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_447 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_446 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_445 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_444 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_443 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_442 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_441 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_111 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_444 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_443 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_442 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_441 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_224 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_223 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_222 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_221 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_GENERIC_NBIT4_56 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_224 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_223 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_222 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_221 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_56 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_112 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_111 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_56 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module FA_440 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_439 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_438 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_437 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_110 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_440 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_439 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_438 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_437 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_436 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_435 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_434 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_433 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_109 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_436 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_435 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_434 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_433 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_220 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_219 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_218 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_217 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_GENERIC_NBIT4_55 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_220 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_219 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_218 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_217 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_55 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_110 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_109 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_55 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module FA_432 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_431 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_430 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_429 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_108 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_432 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_431 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_430 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_429 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_428 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_427 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_426 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_425 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_107 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_428 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_427 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_426 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_425 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_216 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_215 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_214 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_213 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_GENERIC_NBIT4_54 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_216 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_215 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_214 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_213 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_54 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_108 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_107 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_54 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module FA_424 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_423 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_422 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_421 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_106 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_424 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_423 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_422 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_421 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_420 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_419 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_418 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_417 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_105 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_420 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_419 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_418 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_417 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_212 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_211 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_210 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_209 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_GENERIC_NBIT4_53 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_212 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_211 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_210 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_209 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_53 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_106 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_105 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_53 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module FA_416 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_415 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_414 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_413 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_104 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_416 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_415 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_414 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_413 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_412 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_411 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_410 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_409 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_103 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_412 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_411 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_410 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_409 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_208 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_207 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_206 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_205 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_GENERIC_NBIT4_52 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_208 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_207 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_206 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_205 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_52 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_104 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_103 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_52 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module FA_408 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_407 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_406 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_405 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_102 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_408 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_407 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_406 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_405 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_404 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_403 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_402 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_401 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_101 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_404 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_403 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_402 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_401 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_204 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_203 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_202 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_201 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_GENERIC_NBIT4_51 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_204 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_203 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_202 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_201 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_51 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_102 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_101 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_51 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module FA_400 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_399 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_398 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_397 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_100 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_400 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_399 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_398 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_397 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_396 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_395 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_394 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_393 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_99 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_396 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_395 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_394 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_393 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_200 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_199 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_198 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_197 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_GENERIC_NBIT4_50 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_200 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_199 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_198 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_197 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_50 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_100 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_99 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_50 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module FA_392 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_391 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_390 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_389 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_98 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_392 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_391 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_390 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_389 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_388 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_387 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_386 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_385 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_97 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_388 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_387 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_386 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_385 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_196 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_195 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_194 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_193 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_GENERIC_NBIT4_49 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_196 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_195 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_194 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_193 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_49 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_98 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_97 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_49 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module sum_generator_n_bit32_n_CSB8_1 ( A, B, C_in, S );
  input [31:0] A;
  input [31:0] B;
  input [7:0] C_in;
  output [31:0] S;


  carry_select_block_n4_56 csb_0 ( .A(A[3:0]), .B(B[3:0]), .C_sel(C_in[0]), 
        .S(S[3:0]) );
  carry_select_block_n4_55 csb_1 ( .A(A[7:4]), .B(B[7:4]), .C_sel(C_in[1]), 
        .S(S[7:4]) );
  carry_select_block_n4_54 csb_2 ( .A(A[11:8]), .B(B[11:8]), .C_sel(C_in[2]), 
        .S(S[11:8]) );
  carry_select_block_n4_53 csb_3 ( .A(A[15:12]), .B(B[15:12]), .C_sel(C_in[3]), 
        .S(S[15:12]) );
  carry_select_block_n4_52 csb_4 ( .A(A[19:16]), .B(B[19:16]), .C_sel(C_in[4]), 
        .S(S[19:16]) );
  carry_select_block_n4_51 csb_5 ( .A(A[23:20]), .B(B[23:20]), .C_sel(C_in[5]), 
        .S(S[23:20]) );
  carry_select_block_n4_50 csb_6 ( .A(A[27:24]), .B(B[27:24]), .C_sel(C_in[6]), 
        .S(S[27:24]) );
  carry_select_block_n4_49 csb_7 ( .A(A[31:28]), .B(B[31:28]), .C_sel(C_in[7]), 
        .S(S[31:28]) );
endmodule


module P4_ADDER_NBIT32_1 ( A, B, Cin, S, Cout, ovf );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Cin;
  output Cout, ovf;
  wire   n3, n4, n5, n6;
  wire   [31:0] xor_b;
  wire   [6:0] carry;

  XOR2_X1 U3 ( .A(xor_b[31]), .B(A[31]), .Z(n5) );
  my_xor_224 bc_xor_31 ( .A(B[31]), .B(n3), .xor_out(xor_b[31]) );
  my_xor_223 bc_xor_30 ( .A(B[30]), .B(n3), .xor_out(xor_b[30]) );
  my_xor_222 bc_xor_29 ( .A(B[29]), .B(n3), .xor_out(xor_b[29]) );
  my_xor_221 bc_xor_28 ( .A(B[28]), .B(n3), .xor_out(xor_b[28]) );
  my_xor_220 bc_xor_27 ( .A(B[27]), .B(n3), .xor_out(xor_b[27]) );
  my_xor_219 bc_xor_26 ( .A(B[26]), .B(n3), .xor_out(xor_b[26]) );
  my_xor_218 bc_xor_25 ( .A(B[25]), .B(n3), .xor_out(xor_b[25]) );
  my_xor_217 bc_xor_24 ( .A(B[24]), .B(n3), .xor_out(xor_b[24]) );
  my_xor_216 bc_xor_23 ( .A(B[23]), .B(n3), .xor_out(xor_b[23]) );
  my_xor_215 bc_xor_22 ( .A(B[22]), .B(n3), .xor_out(xor_b[22]) );
  my_xor_214 bc_xor_21 ( .A(B[21]), .B(n3), .xor_out(xor_b[21]) );
  my_xor_213 bc_xor_20 ( .A(B[20]), .B(n3), .xor_out(xor_b[20]) );
  my_xor_212 bc_xor_19 ( .A(B[19]), .B(n3), .xor_out(xor_b[19]) );
  my_xor_211 bc_xor_18 ( .A(B[18]), .B(n3), .xor_out(xor_b[18]) );
  my_xor_210 bc_xor_17 ( .A(B[17]), .B(n3), .xor_out(xor_b[17]) );
  my_xor_209 bc_xor_16 ( .A(B[16]), .B(n4), .xor_out(xor_b[16]) );
  my_xor_208 bc_xor_15 ( .A(B[15]), .B(n4), .xor_out(xor_b[15]) );
  my_xor_207 bc_xor_14 ( .A(B[14]), .B(n4), .xor_out(xor_b[14]) );
  my_xor_206 bc_xor_13 ( .A(B[13]), .B(n4), .xor_out(xor_b[13]) );
  my_xor_205 bc_xor_12 ( .A(B[12]), .B(n4), .xor_out(xor_b[12]) );
  my_xor_204 bc_xor_11 ( .A(B[11]), .B(n4), .xor_out(xor_b[11]) );
  my_xor_203 bc_xor_10 ( .A(B[10]), .B(n4), .xor_out(xor_b[10]) );
  my_xor_202 bc_xor_9 ( .A(B[9]), .B(n4), .xor_out(xor_b[9]) );
  my_xor_201 bc_xor_8 ( .A(B[8]), .B(n4), .xor_out(xor_b[8]) );
  my_xor_200 bc_xor_7 ( .A(B[7]), .B(n4), .xor_out(xor_b[7]) );
  my_xor_199 bc_xor_6 ( .A(B[6]), .B(n4), .xor_out(xor_b[6]) );
  my_xor_198 bc_xor_5 ( .A(B[5]), .B(n4), .xor_out(xor_b[5]) );
  my_xor_197 bc_xor_4 ( .A(B[4]), .B(n4), .xor_out(xor_b[4]) );
  my_xor_196 bc_xor_3 ( .A(B[3]), .B(n4), .xor_out(xor_b[3]) );
  my_xor_195 bc_xor_2 ( .A(B[2]), .B(n4), .xor_out(xor_b[2]) );
  my_xor_194 bc_xor_1 ( .A(B[1]), .B(n4), .xor_out(xor_b[1]) );
  my_xor_193 bc_xor_0 ( .A(B[0]), .B(n4), .xor_out(xor_b[0]) );
  CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_1 CG ( .A(A), .B(xor_b), .Cin(n3), 
        .Co({Cout, carry}) );
  sum_generator_n_bit32_n_CSB8_1 SG ( .A(A), .B(xor_b), .C_in({carry, n3}), 
        .S(S) );
  NOR2_X1 U1 ( .A1(n6), .A2(n5), .ZN(ovf) );
  XNOR2_X1 U2 ( .A(A[31]), .B(S[31]), .ZN(n6) );
  BUF_X2 U4 ( .A(Cin), .Z(n3) );
  BUF_X1 U5 ( .A(Cin), .Z(n4) );
endmodule


module nand31_0 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_127 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_126 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_125 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_124 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_123 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_122 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_121 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_120 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_119 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_118 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_117 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_116 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_115 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_114 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_113 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_112 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_111 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_110 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_109 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_108 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_107 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_106 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_105 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_104 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_103 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_102 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_101 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_100 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_99 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_98 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_97 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_96 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_95 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_94 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_93 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_92 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_91 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_90 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_89 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_88 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_87 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_86 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_85 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_84 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_83 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_82 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_81 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_80 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_79 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_78 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_77 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_76 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_75 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_74 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_73 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_72 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_71 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_70 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_69 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_68 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_67 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_66 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_65 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_64 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_63 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_62 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_61 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_60 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_59 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_58 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_57 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_56 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_55 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_54 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_53 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_52 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_51 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_50 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_49 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_48 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_47 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_46 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_45 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_44 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_43 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_42 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_41 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_40 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_39 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_38 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_37 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_36 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_35 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_34 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_33 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_32 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_31 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_30 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_29 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_28 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_27 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_26 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_25 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_24 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_23 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_22 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_21 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_20 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_19 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_18 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_17 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_16 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_15 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_14 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_13 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_12 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_11 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_10 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_9 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_8 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_7 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_6 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_5 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_4 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_3 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_2 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand31_1 ( in1, in2, in3, o );
  input in1, in2, in3;
  output o;


  NAND3_X1 U1 ( .A1(in2), .A2(in1), .A3(in3), .ZN(o) );
endmodule


module nand41_0 ( in1, in2, in3, in4, o );
  input in1, in2, in3, in4;
  output o;


  NAND4_X1 U1 ( .A1(in4), .A2(in3), .A3(in2), .A4(in1), .ZN(o) );
endmodule


module nand41_31 ( in1, in2, in3, in4, o );
  input in1, in2, in3, in4;
  output o;


  NAND4_X1 U1 ( .A1(in4), .A2(in3), .A3(in2), .A4(in1), .ZN(o) );
endmodule


module nand41_30 ( in1, in2, in3, in4, o );
  input in1, in2, in3, in4;
  output o;


  NAND4_X1 U1 ( .A1(in4), .A2(in3), .A3(in2), .A4(in1), .ZN(o) );
endmodule


module nand41_29 ( in1, in2, in3, in4, o );
  input in1, in2, in3, in4;
  output o;


  NAND4_X1 U1 ( .A1(in4), .A2(in3), .A3(in2), .A4(in1), .ZN(o) );
endmodule


module nand41_28 ( in1, in2, in3, in4, o );
  input in1, in2, in3, in4;
  output o;


  NAND4_X1 U1 ( .A1(in4), .A2(in3), .A3(in2), .A4(in1), .ZN(o) );
endmodule


module nand41_27 ( in1, in2, in3, in4, o );
  input in1, in2, in3, in4;
  output o;


  NAND4_X1 U1 ( .A1(in4), .A2(in3), .A3(in2), .A4(in1), .ZN(o) );
endmodule


module nand41_26 ( in1, in2, in3, in4, o );
  input in1, in2, in3, in4;
  output o;


  NAND4_X1 U1 ( .A1(in4), .A2(in3), .A3(in2), .A4(in1), .ZN(o) );
endmodule


module nand41_25 ( in1, in2, in3, in4, o );
  input in1, in2, in3, in4;
  output o;


  NAND4_X1 U1 ( .A1(in4), .A2(in3), .A3(in2), .A4(in1), .ZN(o) );
endmodule


module nand41_24 ( in1, in2, in3, in4, o );
  input in1, in2, in3, in4;
  output o;


  NAND4_X1 U1 ( .A1(in4), .A2(in3), .A3(in2), .A4(in1), .ZN(o) );
endmodule


module nand41_23 ( in1, in2, in3, in4, o );
  input in1, in2, in3, in4;
  output o;


  NAND4_X1 U1 ( .A1(in4), .A2(in3), .A3(in2), .A4(in1), .ZN(o) );
endmodule


module nand41_22 ( in1, in2, in3, in4, o );
  input in1, in2, in3, in4;
  output o;


  NAND4_X1 U1 ( .A1(in4), .A2(in3), .A3(in2), .A4(in1), .ZN(o) );
endmodule


module nand41_21 ( in1, in2, in3, in4, o );
  input in1, in2, in3, in4;
  output o;


  NAND4_X1 U1 ( .A1(in4), .A2(in3), .A3(in2), .A4(in1), .ZN(o) );
endmodule


module nand41_20 ( in1, in2, in3, in4, o );
  input in1, in2, in3, in4;
  output o;


  NAND4_X1 U1 ( .A1(in4), .A2(in3), .A3(in2), .A4(in1), .ZN(o) );
endmodule


module nand41_19 ( in1, in2, in3, in4, o );
  input in1, in2, in3, in4;
  output o;


  NAND4_X1 U1 ( .A1(in4), .A2(in3), .A3(in2), .A4(in1), .ZN(o) );
endmodule


module nand41_18 ( in1, in2, in3, in4, o );
  input in1, in2, in3, in4;
  output o;


  NAND4_X1 U1 ( .A1(in4), .A2(in3), .A3(in2), .A4(in1), .ZN(o) );
endmodule


module nand41_17 ( in1, in2, in3, in4, o );
  input in1, in2, in3, in4;
  output o;


  NAND4_X1 U1 ( .A1(in4), .A2(in3), .A3(in2), .A4(in1), .ZN(o) );
endmodule


module nand41_16 ( in1, in2, in3, in4, o );
  input in1, in2, in3, in4;
  output o;


  NAND4_X1 U1 ( .A1(in4), .A2(in3), .A3(in2), .A4(in1), .ZN(o) );
endmodule


module nand41_15 ( in1, in2, in3, in4, o );
  input in1, in2, in3, in4;
  output o;


  NAND4_X1 U1 ( .A1(in4), .A2(in3), .A3(in2), .A4(in1), .ZN(o) );
endmodule


module nand41_14 ( in1, in2, in3, in4, o );
  input in1, in2, in3, in4;
  output o;


  NAND4_X1 U1 ( .A1(in4), .A2(in3), .A3(in2), .A4(in1), .ZN(o) );
endmodule


module nand41_13 ( in1, in2, in3, in4, o );
  input in1, in2, in3, in4;
  output o;


  NAND4_X1 U1 ( .A1(in4), .A2(in3), .A3(in2), .A4(in1), .ZN(o) );
endmodule


module nand41_12 ( in1, in2, in3, in4, o );
  input in1, in2, in3, in4;
  output o;


  NAND4_X1 U1 ( .A1(in4), .A2(in3), .A3(in2), .A4(in1), .ZN(o) );
endmodule


module nand41_11 ( in1, in2, in3, in4, o );
  input in1, in2, in3, in4;
  output o;


  NAND4_X1 U1 ( .A1(in4), .A2(in3), .A3(in2), .A4(in1), .ZN(o) );
endmodule


module nand41_10 ( in1, in2, in3, in4, o );
  input in1, in2, in3, in4;
  output o;


  NAND4_X1 U1 ( .A1(in4), .A2(in3), .A3(in2), .A4(in1), .ZN(o) );
endmodule


module nand41_9 ( in1, in2, in3, in4, o );
  input in1, in2, in3, in4;
  output o;


  NAND4_X1 U1 ( .A1(in4), .A2(in3), .A3(in2), .A4(in1), .ZN(o) );
endmodule


module nand41_8 ( in1, in2, in3, in4, o );
  input in1, in2, in3, in4;
  output o;


  NAND4_X1 U1 ( .A1(in4), .A2(in3), .A3(in2), .A4(in1), .ZN(o) );
endmodule


module nand41_7 ( in1, in2, in3, in4, o );
  input in1, in2, in3, in4;
  output o;


  NAND4_X1 U1 ( .A1(in4), .A2(in3), .A3(in2), .A4(in1), .ZN(o) );
endmodule


module nand41_6 ( in1, in2, in3, in4, o );
  input in1, in2, in3, in4;
  output o;


  NAND4_X1 U1 ( .A1(in4), .A2(in3), .A3(in2), .A4(in1), .ZN(o) );
endmodule


module nand41_5 ( in1, in2, in3, in4, o );
  input in1, in2, in3, in4;
  output o;


  NAND4_X1 U1 ( .A1(in4), .A2(in3), .A3(in2), .A4(in1), .ZN(o) );
endmodule


module nand41_4 ( in1, in2, in3, in4, o );
  input in1, in2, in3, in4;
  output o;


  NAND4_X1 U1 ( .A1(in4), .A2(in3), .A3(in2), .A4(in1), .ZN(o) );
endmodule


module nand41_3 ( in1, in2, in3, in4, o );
  input in1, in2, in3, in4;
  output o;


  NAND4_X1 U1 ( .A1(in4), .A2(in3), .A3(in2), .A4(in1), .ZN(o) );
endmodule


module nand41_2 ( in1, in2, in3, in4, o );
  input in1, in2, in3, in4;
  output o;


  NAND4_X1 U1 ( .A1(in4), .A2(in3), .A3(in2), .A4(in1), .ZN(o) );
endmodule


module nand41_1 ( in1, in2, in3, in4, o );
  input in1, in2, in3, in4;
  output o;


  NAND4_X1 U1 ( .A1(in4), .A2(in3), .A3(in2), .A4(in1), .ZN(o) );
endmodule


module logicals_nbit32 ( func, SN, in1, in2, o );
  input [3:0] func;
  input [31:0] in1;
  input [31:0] in2;
  output [31:0] o;
  input SN;
  wire   \s0[9] , \s2[9] , \s3[9] , n69, n70, n71, n72, n73, n74, n1, n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86;
  wire   [31:0] l0;
  wire   [31:0] l1;
  wire   [31:0] l2;
  wire   [31:0] l3;

  NAND3_X1 U77 ( .A1(n69), .A2(n71), .A3(n72), .ZN(\s2[9] ) );
  NAND3_X1 U78 ( .A1(n73), .A2(n86), .A3(func[0]), .ZN(n72) );
  NAND3_X1 U79 ( .A1(n73), .A2(n21), .A3(SN), .ZN(n71) );
  nand31_0 g1_a_31 ( .in1(n12), .in2(n18), .in3(n85), .o(l0[31]) );
  nand31_127 g1_b_31 ( .in1(n4), .in2(n18), .in3(in2[31]), .o(l1[31]) );
  nand31_126 g1_c_31 ( .in1(n4), .in2(in1[31]), .in3(n85), .o(l2[31]) );
  nand31_125 g1_d_31 ( .in1(n3), .in2(in1[31]), .in3(in2[31]), .o(l3[31]) );
  nand31_124 g1_a_30 ( .in1(n10), .in2(n51), .in3(n84), .o(l0[30]) );
  nand31_123 g1_b_30 ( .in1(n4), .in2(n51), .in3(in2[30]), .o(l1[30]) );
  nand31_122 g1_c_30 ( .in1(n4), .in2(in1[30]), .in3(n84), .o(l2[30]) );
  nand31_121 g1_d_30 ( .in1(n3), .in2(in1[30]), .in3(in2[30]), .o(l3[30]) );
  nand31_120 g1_a_29 ( .in1(n10), .in2(n50), .in3(n83), .o(l0[29]) );
  nand31_119 g1_b_29 ( .in1(n4), .in2(n50), .in3(in2[29]), .o(l1[29]) );
  nand31_118 g1_c_29 ( .in1(n4), .in2(in1[29]), .in3(n83), .o(l2[29]) );
  nand31_117 g1_d_29 ( .in1(n3), .in2(in1[29]), .in3(in2[29]), .o(l3[29]) );
  nand31_116 g1_a_28 ( .in1(n10), .in2(n49), .in3(n82), .o(l0[28]) );
  nand31_115 g1_b_28 ( .in1(n4), .in2(n49), .in3(in2[28]), .o(l1[28]) );
  nand31_114 g1_c_28 ( .in1(n4), .in2(in1[28]), .in3(n82), .o(l2[28]) );
  nand31_113 g1_d_28 ( .in1(n3), .in2(in1[28]), .in3(in2[28]), .o(l3[28]) );
  nand31_112 g1_a_27 ( .in1(n10), .in2(n48), .in3(n81), .o(l0[27]) );
  nand31_111 g1_b_27 ( .in1(n4), .in2(n48), .in3(in2[27]), .o(l1[27]) );
  nand31_110 g1_c_27 ( .in1(n4), .in2(in1[27]), .in3(n81), .o(l2[27]) );
  nand31_109 g1_d_27 ( .in1(n3), .in2(in1[27]), .in3(in2[27]), .o(l3[27]) );
  nand31_108 g1_a_26 ( .in1(n10), .in2(n47), .in3(n80), .o(l0[26]) );
  nand31_107 g1_b_26 ( .in1(n4), .in2(n47), .in3(in2[26]), .o(l1[26]) );
  nand31_106 g1_c_26 ( .in1(n5), .in2(in1[26]), .in3(n80), .o(l2[26]) );
  nand31_105 g1_d_26 ( .in1(n3), .in2(in1[26]), .in3(in2[26]), .o(l3[26]) );
  nand31_104 g1_a_25 ( .in1(n10), .in2(n46), .in3(n79), .o(l0[25]) );
  nand31_103 g1_b_25 ( .in1(n5), .in2(n46), .in3(in2[25]), .o(l1[25]) );
  nand31_102 g1_c_25 ( .in1(n5), .in2(in1[25]), .in3(n79), .o(l2[25]) );
  nand31_101 g1_d_25 ( .in1(n3), .in2(in1[25]), .in3(in2[25]), .o(l3[25]) );
  nand31_100 g1_a_24 ( .in1(n10), .in2(n45), .in3(n78), .o(l0[24]) );
  nand31_99 g1_b_24 ( .in1(n5), .in2(n45), .in3(in2[24]), .o(l1[24]) );
  nand31_98 g1_c_24 ( .in1(n5), .in2(in1[24]), .in3(n78), .o(l2[24]) );
  nand31_97 g1_d_24 ( .in1(n3), .in2(in1[24]), .in3(in2[24]), .o(l3[24]) );
  nand31_96 g1_a_23 ( .in1(n10), .in2(n44), .in3(n77), .o(l0[23]) );
  nand31_95 g1_b_23 ( .in1(n5), .in2(n44), .in3(in2[23]), .o(l1[23]) );
  nand31_94 g1_c_23 ( .in1(n5), .in2(in1[23]), .in3(n77), .o(l2[23]) );
  nand31_93 g1_d_23 ( .in1(n3), .in2(in1[23]), .in3(in2[23]), .o(l3[23]) );
  nand31_92 g1_a_22 ( .in1(n10), .in2(n43), .in3(n76), .o(l0[22]) );
  nand31_91 g1_b_22 ( .in1(n5), .in2(n43), .in3(in2[22]), .o(l1[22]) );
  nand31_90 g1_c_22 ( .in1(n5), .in2(in1[22]), .in3(n76), .o(l2[22]) );
  nand31_89 g1_d_22 ( .in1(n3), .in2(in1[22]), .in3(in2[22]), .o(l3[22]) );
  nand31_88 g1_a_21 ( .in1(n10), .in2(n42), .in3(n75), .o(l0[21]) );
  nand31_87 g1_b_21 ( .in1(n5), .in2(n42), .in3(in2[21]), .o(l1[21]) );
  nand31_86 g1_c_21 ( .in1(n5), .in2(in1[21]), .in3(n75), .o(l2[21]) );
  nand31_85 g1_d_21 ( .in1(n2), .in2(in1[21]), .in3(in2[21]), .o(l3[21]) );
  nand31_84 g1_a_20 ( .in1(n10), .in2(n41), .in3(n68), .o(l0[20]) );
  nand31_83 g1_b_20 ( .in1(n6), .in2(n41), .in3(in2[20]), .o(l1[20]) );
  nand31_82 g1_c_20 ( .in1(n6), .in2(in1[20]), .in3(n68), .o(l2[20]) );
  nand31_81 g1_d_20 ( .in1(n2), .in2(in1[20]), .in3(in2[20]), .o(l3[20]) );
  nand31_80 g1_a_19 ( .in1(n11), .in2(n40), .in3(n67), .o(l0[19]) );
  nand31_79 g1_b_19 ( .in1(n6), .in2(n40), .in3(in2[19]), .o(l1[19]) );
  nand31_78 g1_c_19 ( .in1(n6), .in2(in1[19]), .in3(n67), .o(l2[19]) );
  nand31_77 g1_d_19 ( .in1(n2), .in2(in1[19]), .in3(in2[19]), .o(l3[19]) );
  nand31_76 g1_a_18 ( .in1(n11), .in2(n39), .in3(n66), .o(l0[18]) );
  nand31_75 g1_b_18 ( .in1(n6), .in2(n39), .in3(in2[18]), .o(l1[18]) );
  nand31_74 g1_c_18 ( .in1(n6), .in2(in1[18]), .in3(n66), .o(l2[18]) );
  nand31_73 g1_d_18 ( .in1(n2), .in2(in1[18]), .in3(in2[18]), .o(l3[18]) );
  nand31_72 g1_a_17 ( .in1(n11), .in2(n38), .in3(n65), .o(l0[17]) );
  nand31_71 g1_b_17 ( .in1(n6), .in2(n38), .in3(in2[17]), .o(l1[17]) );
  nand31_70 g1_c_17 ( .in1(n6), .in2(in1[17]), .in3(n65), .o(l2[17]) );
  nand31_69 g1_d_17 ( .in1(n2), .in2(in1[17]), .in3(in2[17]), .o(l3[17]) );
  nand31_68 g1_a_16 ( .in1(n11), .in2(n37), .in3(n64), .o(l0[16]) );
  nand31_67 g1_b_16 ( .in1(n6), .in2(n37), .in3(in2[16]), .o(l1[16]) );
  nand31_66 g1_c_16 ( .in1(n6), .in2(in1[16]), .in3(n64), .o(l2[16]) );
  nand31_65 g1_d_16 ( .in1(n2), .in2(in1[16]), .in3(in2[16]), .o(l3[16]) );
  nand31_64 g1_a_15 ( .in1(n11), .in2(n36), .in3(n63), .o(l0[15]) );
  nand31_63 g1_b_15 ( .in1(n6), .in2(n36), .in3(in2[15]), .o(l1[15]) );
  nand31_62 g1_c_15 ( .in1(n7), .in2(in1[15]), .in3(n63), .o(l2[15]) );
  nand31_61 g1_d_15 ( .in1(n2), .in2(in1[15]), .in3(in2[15]), .o(l3[15]) );
  nand31_60 g1_a_14 ( .in1(n11), .in2(n35), .in3(n62), .o(l0[14]) );
  nand31_59 g1_b_14 ( .in1(n7), .in2(n35), .in3(in2[14]), .o(l1[14]) );
  nand31_58 g1_c_14 ( .in1(n7), .in2(in1[14]), .in3(n62), .o(l2[14]) );
  nand31_57 g1_d_14 ( .in1(n2), .in2(in1[14]), .in3(in2[14]), .o(l3[14]) );
  nand31_56 g1_a_13 ( .in1(n11), .in2(n34), .in3(n61), .o(l0[13]) );
  nand31_55 g1_b_13 ( .in1(n7), .in2(n34), .in3(in2[13]), .o(l1[13]) );
  nand31_54 g1_c_13 ( .in1(n7), .in2(in1[13]), .in3(n61), .o(l2[13]) );
  nand31_53 g1_d_13 ( .in1(n2), .in2(in1[13]), .in3(in2[13]), .o(l3[13]) );
  nand31_52 g1_a_12 ( .in1(n11), .in2(n33), .in3(n60), .o(l0[12]) );
  nand31_51 g1_b_12 ( .in1(n7), .in2(n33), .in3(in2[12]), .o(l1[12]) );
  nand31_50 g1_c_12 ( .in1(n7), .in2(in1[12]), .in3(n60), .o(l2[12]) );
  nand31_49 g1_d_12 ( .in1(n2), .in2(in1[12]), .in3(in2[12]), .o(l3[12]) );
  nand31_48 g1_a_11 ( .in1(n11), .in2(n32), .in3(n59), .o(l0[11]) );
  nand31_47 g1_b_11 ( .in1(n7), .in2(n32), .in3(in2[11]), .o(l1[11]) );
  nand31_46 g1_c_11 ( .in1(n7), .in2(in1[11]), .in3(n59), .o(l2[11]) );
  nand31_45 g1_d_11 ( .in1(n2), .in2(in1[11]), .in3(in2[11]), .o(l3[11]) );
  nand31_44 g1_a_10 ( .in1(n11), .in2(n31), .in3(n58), .o(l0[10]) );
  nand31_43 g1_b_10 ( .in1(n7), .in2(n31), .in3(in2[10]), .o(l1[10]) );
  nand31_42 g1_c_10 ( .in1(n7), .in2(in1[10]), .in3(n58), .o(l2[10]) );
  nand31_41 g1_d_10 ( .in1(n1), .in2(in1[10]), .in3(in2[10]), .o(l3[10]) );
  nand31_40 g1_a_9 ( .in1(n11), .in2(n30), .in3(n57), .o(l0[9]) );
  nand31_39 g1_b_9 ( .in1(n8), .in2(n30), .in3(in2[9]), .o(l1[9]) );
  nand31_38 g1_c_9 ( .in1(n8), .in2(in1[9]), .in3(n57), .o(l2[9]) );
  nand31_37 g1_d_9 ( .in1(n1), .in2(in1[9]), .in3(in2[9]), .o(l3[9]) );
  nand31_36 g1_a_8 ( .in1(n12), .in2(n29), .in3(n56), .o(l0[8]) );
  nand31_35 g1_b_8 ( .in1(n8), .in2(n29), .in3(in2[8]), .o(l1[8]) );
  nand31_34 g1_c_8 ( .in1(n8), .in2(in1[8]), .in3(n56), .o(l2[8]) );
  nand31_33 g1_d_8 ( .in1(n1), .in2(in1[8]), .in3(in2[8]), .o(l3[8]) );
  nand31_32 g1_a_7 ( .in1(n12), .in2(n28), .in3(n55), .o(l0[7]) );
  nand31_31 g1_b_7 ( .in1(n8), .in2(n28), .in3(in2[7]), .o(l1[7]) );
  nand31_30 g1_c_7 ( .in1(n8), .in2(in1[7]), .in3(n55), .o(l2[7]) );
  nand31_29 g1_d_7 ( .in1(n1), .in2(in1[7]), .in3(in2[7]), .o(l3[7]) );
  nand31_28 g1_a_6 ( .in1(n12), .in2(n27), .in3(n54), .o(l0[6]) );
  nand31_27 g1_b_6 ( .in1(n8), .in2(n27), .in3(in2[6]), .o(l1[6]) );
  nand31_26 g1_c_6 ( .in1(n8), .in2(in1[6]), .in3(n54), .o(l2[6]) );
  nand31_25 g1_d_6 ( .in1(n1), .in2(in1[6]), .in3(in2[6]), .o(l3[6]) );
  nand31_24 g1_a_5 ( .in1(n12), .in2(n26), .in3(n53), .o(l0[5]) );
  nand31_23 g1_b_5 ( .in1(n8), .in2(n26), .in3(in2[5]), .o(l1[5]) );
  nand31_22 g1_c_5 ( .in1(n8), .in2(in1[5]), .in3(n53), .o(l2[5]) );
  nand31_21 g1_d_5 ( .in1(n1), .in2(in1[5]), .in3(in2[5]), .o(l3[5]) );
  nand31_20 g1_a_4 ( .in1(n12), .in2(n25), .in3(n17), .o(l0[4]) );
  nand31_19 g1_b_4 ( .in1(n8), .in2(n25), .in3(in2[4]), .o(l1[4]) );
  nand31_18 g1_c_4 ( .in1(n9), .in2(in1[4]), .in3(n17), .o(l2[4]) );
  nand31_17 g1_d_4 ( .in1(n1), .in2(in1[4]), .in3(in2[4]), .o(l3[4]) );
  nand31_16 g1_a_3 ( .in1(n12), .in2(n24), .in3(n16), .o(l0[3]) );
  nand31_15 g1_b_3 ( .in1(n9), .in2(n24), .in3(in2[3]), .o(l1[3]) );
  nand31_14 g1_c_3 ( .in1(n9), .in2(in1[3]), .in3(n16), .o(l2[3]) );
  nand31_13 g1_d_3 ( .in1(n1), .in2(in1[3]), .in3(in2[3]), .o(l3[3]) );
  nand31_12 g1_a_2 ( .in1(n12), .in2(n23), .in3(n15), .o(l0[2]) );
  nand31_11 g1_b_2 ( .in1(n9), .in2(n23), .in3(in2[2]), .o(l1[2]) );
  nand31_10 g1_c_2 ( .in1(n9), .in2(in1[2]), .in3(n15), .o(l2[2]) );
  nand31_9 g1_d_2 ( .in1(n1), .in2(in1[2]), .in3(in2[2]), .o(l3[2]) );
  nand31_8 g1_a_1 ( .in1(n12), .in2(n22), .in3(n14), .o(l0[1]) );
  nand31_7 g1_b_1 ( .in1(n9), .in2(n22), .in3(in2[1]), .o(l1[1]) );
  nand31_6 g1_c_1 ( .in1(n9), .in2(in1[1]), .in3(n14), .o(l2[1]) );
  nand31_5 g1_d_1 ( .in1(n1), .in2(in1[1]), .in3(in2[1]), .o(l3[1]) );
  nand31_4 g1_a_0 ( .in1(n12), .in2(n52), .in3(n13), .o(l0[0]) );
  nand31_3 g1_b_0 ( .in1(n9), .in2(n52), .in3(in2[0]), .o(l1[0]) );
  nand31_2 g1_c_0 ( .in1(n9), .in2(in1[0]), .in3(n13), .o(l2[0]) );
  nand31_1 g1_d_0 ( .in1(n1), .in2(in1[0]), .in3(in2[0]), .o(l3[0]) );
  nand41_0 g2_a_31 ( .in1(l0[31]), .in2(l1[31]), .in3(l2[31]), .in4(l3[31]), 
        .o(o[31]) );
  nand41_31 g2_a_30 ( .in1(l0[30]), .in2(l1[30]), .in3(l2[30]), .in4(l3[30]), 
        .o(o[30]) );
  nand41_30 g2_a_29 ( .in1(l0[29]), .in2(l1[29]), .in3(l2[29]), .in4(l3[29]), 
        .o(o[29]) );
  nand41_29 g2_a_28 ( .in1(l0[28]), .in2(l1[28]), .in3(l2[28]), .in4(l3[28]), 
        .o(o[28]) );
  nand41_28 g2_a_27 ( .in1(l0[27]), .in2(l1[27]), .in3(l2[27]), .in4(l3[27]), 
        .o(o[27]) );
  nand41_27 g2_a_26 ( .in1(l0[26]), .in2(l1[26]), .in3(l2[26]), .in4(l3[26]), 
        .o(o[26]) );
  nand41_26 g2_a_25 ( .in1(l0[25]), .in2(l1[25]), .in3(l2[25]), .in4(l3[25]), 
        .o(o[25]) );
  nand41_25 g2_a_24 ( .in1(l0[24]), .in2(l1[24]), .in3(l2[24]), .in4(l3[24]), 
        .o(o[24]) );
  nand41_24 g2_a_23 ( .in1(l0[23]), .in2(l1[23]), .in3(l2[23]), .in4(l3[23]), 
        .o(o[23]) );
  nand41_23 g2_a_22 ( .in1(l0[22]), .in2(l1[22]), .in3(l2[22]), .in4(l3[22]), 
        .o(o[22]) );
  nand41_22 g2_a_21 ( .in1(l0[21]), .in2(l1[21]), .in3(l2[21]), .in4(l3[21]), 
        .o(o[21]) );
  nand41_21 g2_a_20 ( .in1(l0[20]), .in2(l1[20]), .in3(l2[20]), .in4(l3[20]), 
        .o(o[20]) );
  nand41_20 g2_a_19 ( .in1(l0[19]), .in2(l1[19]), .in3(l2[19]), .in4(l3[19]), 
        .o(o[19]) );
  nand41_19 g2_a_18 ( .in1(l0[18]), .in2(l1[18]), .in3(l2[18]), .in4(l3[18]), 
        .o(o[18]) );
  nand41_18 g2_a_17 ( .in1(l0[17]), .in2(l1[17]), .in3(l2[17]), .in4(l3[17]), 
        .o(o[17]) );
  nand41_17 g2_a_16 ( .in1(l0[16]), .in2(l1[16]), .in3(l2[16]), .in4(l3[16]), 
        .o(o[16]) );
  nand41_16 g2_a_15 ( .in1(l0[15]), .in2(l1[15]), .in3(l2[15]), .in4(l3[15]), 
        .o(o[15]) );
  nand41_15 g2_a_14 ( .in1(l0[14]), .in2(l1[14]), .in3(l2[14]), .in4(l3[14]), 
        .o(o[14]) );
  nand41_14 g2_a_13 ( .in1(l0[13]), .in2(l1[13]), .in3(l2[13]), .in4(l3[13]), 
        .o(o[13]) );
  nand41_13 g2_a_12 ( .in1(l0[12]), .in2(l1[12]), .in3(l2[12]), .in4(l3[12]), 
        .o(o[12]) );
  nand41_12 g2_a_11 ( .in1(l0[11]), .in2(l1[11]), .in3(l2[11]), .in4(l3[11]), 
        .o(o[11]) );
  nand41_11 g2_a_10 ( .in1(l0[10]), .in2(l1[10]), .in3(l2[10]), .in4(l3[10]), 
        .o(o[10]) );
  nand41_10 g2_a_9 ( .in1(l0[9]), .in2(l1[9]), .in3(l2[9]), .in4(l3[9]), .o(
        o[9]) );
  nand41_9 g2_a_8 ( .in1(l0[8]), .in2(l1[8]), .in3(l2[8]), .in4(l3[8]), .o(
        o[8]) );
  nand41_8 g2_a_7 ( .in1(l0[7]), .in2(l1[7]), .in3(l2[7]), .in4(l3[7]), .o(
        o[7]) );
  nand41_7 g2_a_6 ( .in1(l0[6]), .in2(l1[6]), .in3(l2[6]), .in4(l3[6]), .o(
        o[6]) );
  nand41_6 g2_a_5 ( .in1(l0[5]), .in2(l1[5]), .in3(l2[5]), .in4(l3[5]), .o(
        o[5]) );
  nand41_5 g2_a_4 ( .in1(l0[4]), .in2(l1[4]), .in3(l2[4]), .in4(l3[4]), .o(
        o[4]) );
  nand41_4 g2_a_3 ( .in1(l0[3]), .in2(l1[3]), .in3(l2[3]), .in4(l3[3]), .o(
        o[3]) );
  nand41_3 g2_a_2 ( .in1(l0[2]), .in2(l1[2]), .in3(l2[2]), .in4(l3[2]), .o(
        o[2]) );
  nand41_2 g2_a_1 ( .in1(l0[1]), .in2(l1[1]), .in3(l2[1]), .in4(l3[1]), .o(
        o[1]) );
  nand41_1 g2_a_0 ( .in1(l0[0]), .in2(l1[0]), .in3(l2[0]), .in4(l3[0]), .o(
        o[0]) );
  BUF_X1 U3 ( .A(\s0[9] ), .Z(n10) );
  BUF_X1 U4 ( .A(\s0[9] ), .Z(n11) );
  BUF_X1 U5 ( .A(\s3[9] ), .Z(n2) );
  BUF_X1 U6 ( .A(\s3[9] ), .Z(n1) );
  BUF_X1 U7 ( .A(\s0[9] ), .Z(n12) );
  BUF_X1 U8 ( .A(\s3[9] ), .Z(n3) );
  INV_X1 U9 ( .A(in1[0]), .ZN(n52) );
  INV_X1 U10 ( .A(in1[28]), .ZN(n49) );
  INV_X1 U11 ( .A(in1[27]), .ZN(n48) );
  INV_X1 U12 ( .A(in1[26]), .ZN(n47) );
  INV_X1 U13 ( .A(in1[25]), .ZN(n46) );
  INV_X1 U14 ( .A(in1[24]), .ZN(n45) );
  INV_X1 U15 ( .A(in1[7]), .ZN(n28) );
  INV_X1 U16 ( .A(in1[6]), .ZN(n27) );
  INV_X1 U17 ( .A(in1[5]), .ZN(n26) );
  INV_X1 U18 ( .A(in1[4]), .ZN(n25) );
  INV_X1 U19 ( .A(in1[3]), .ZN(n24) );
  INV_X1 U20 ( .A(in1[2]), .ZN(n23) );
  INV_X1 U21 ( .A(in1[1]), .ZN(n22) );
  INV_X1 U22 ( .A(in1[23]), .ZN(n44) );
  INV_X1 U23 ( .A(in1[22]), .ZN(n43) );
  INV_X1 U24 ( .A(in1[21]), .ZN(n42) );
  INV_X1 U25 ( .A(in1[20]), .ZN(n41) );
  INV_X1 U26 ( .A(in1[19]), .ZN(n40) );
  INV_X1 U27 ( .A(in1[18]), .ZN(n39) );
  INV_X1 U28 ( .A(in1[17]), .ZN(n38) );
  INV_X1 U29 ( .A(in1[16]), .ZN(n37) );
  INV_X1 U30 ( .A(in1[15]), .ZN(n36) );
  INV_X1 U31 ( .A(in1[14]), .ZN(n35) );
  INV_X1 U32 ( .A(in1[13]), .ZN(n34) );
  INV_X1 U33 ( .A(in1[12]), .ZN(n33) );
  INV_X1 U34 ( .A(in1[11]), .ZN(n32) );
  INV_X1 U35 ( .A(in1[10]), .ZN(n31) );
  INV_X1 U36 ( .A(in1[9]), .ZN(n30) );
  INV_X1 U37 ( .A(in1[8]), .ZN(n29) );
  INV_X1 U38 ( .A(in1[29]), .ZN(n50) );
  INV_X1 U39 ( .A(in1[30]), .ZN(n51) );
  INV_X1 U40 ( .A(in2[5]), .ZN(n53) );
  BUF_X1 U41 ( .A(\s2[9] ), .Z(n4) );
  BUF_X1 U42 ( .A(\s2[9] ), .Z(n5) );
  BUF_X1 U43 ( .A(\s2[9] ), .Z(n6) );
  BUF_X1 U44 ( .A(\s2[9] ), .Z(n7) );
  BUF_X1 U45 ( .A(\s2[9] ), .Z(n8) );
  BUF_X1 U46 ( .A(\s2[9] ), .Z(n9) );
  OAI21_X1 U47 ( .B1(n86), .B2(n74), .A(n70), .ZN(\s0[9] ) );
  INV_X1 U48 ( .A(in2[7]), .ZN(n55) );
  INV_X1 U49 ( .A(in2[6]), .ZN(n54) );
  INV_X1 U50 ( .A(in2[31]), .ZN(n85) );
  INV_X1 U51 ( .A(in2[8]), .ZN(n56) );
  INV_X1 U52 ( .A(in2[30]), .ZN(n84) );
  INV_X1 U53 ( .A(in2[29]), .ZN(n83) );
  INV_X1 U54 ( .A(in2[28]), .ZN(n82) );
  INV_X1 U55 ( .A(in2[27]), .ZN(n81) );
  INV_X1 U56 ( .A(in2[26]), .ZN(n80) );
  INV_X1 U57 ( .A(in2[25]), .ZN(n79) );
  INV_X1 U58 ( .A(in2[24]), .ZN(n78) );
  INV_X1 U59 ( .A(in2[23]), .ZN(n77) );
  INV_X1 U60 ( .A(in2[22]), .ZN(n76) );
  INV_X1 U61 ( .A(in2[21]), .ZN(n75) );
  INV_X1 U62 ( .A(in2[20]), .ZN(n68) );
  INV_X1 U63 ( .A(in2[19]), .ZN(n67) );
  INV_X1 U64 ( .A(in2[18]), .ZN(n66) );
  INV_X1 U65 ( .A(in2[17]), .ZN(n65) );
  INV_X1 U66 ( .A(in2[16]), .ZN(n64) );
  INV_X1 U67 ( .A(in2[15]), .ZN(n63) );
  INV_X1 U68 ( .A(in2[14]), .ZN(n62) );
  INV_X1 U69 ( .A(in2[13]), .ZN(n61) );
  INV_X1 U70 ( .A(in2[12]), .ZN(n60) );
  INV_X1 U71 ( .A(in2[11]), .ZN(n59) );
  INV_X1 U72 ( .A(in2[10]), .ZN(n58) );
  INV_X1 U73 ( .A(in2[9]), .ZN(n57) );
  AND2_X1 U74 ( .A1(n69), .A2(n70), .ZN(\s3[9] ) );
  NAND2_X1 U75 ( .A1(SN), .A2(n73), .ZN(n70) );
  INV_X1 U76 ( .A(SN), .ZN(n86) );
  OR2_X1 U80 ( .A1(n74), .A2(SN), .ZN(n69) );
  NOR3_X1 U81 ( .A1(func[2]), .A2(func[3]), .A3(n20), .ZN(n73) );
  NAND4_X1 U82 ( .A1(func[2]), .A2(n21), .A3(n20), .A4(n19), .ZN(n74) );
  INV_X1 U83 ( .A(func[3]), .ZN(n19) );
  INV_X1 U84 ( .A(func[1]), .ZN(n20) );
  INV_X1 U85 ( .A(func[0]), .ZN(n21) );
  INV_X1 U86 ( .A(in2[0]), .ZN(n13) );
  INV_X1 U87 ( .A(in2[1]), .ZN(n14) );
  INV_X1 U88 ( .A(in2[2]), .ZN(n15) );
  INV_X1 U89 ( .A(in2[3]), .ZN(n16) );
  INV_X1 U90 ( .A(in2[4]), .ZN(n17) );
  INV_X1 U91 ( .A(in1[31]), .ZN(n18) );
endmodule


module nor_generic_NBITS32 ( \input , result );
  input [31:0] \input ;
  output result;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10;

  NOR4_X1 U1 ( .A1(\input [1]), .A2(\input [19]), .A3(\input [18]), .A4(
        \input [17]), .ZN(n5) );
  NOR4_X1 U2 ( .A1(\input [9]), .A2(\input [8]), .A3(\input [7]), .A4(
        \input [6]), .ZN(n10) );
  NOR4_X1 U3 ( .A1(\input [23]), .A2(\input [22]), .A3(\input [21]), .A4(
        \input [20]), .ZN(n6) );
  NOR4_X1 U4 ( .A1(\input [5]), .A2(\input [4]), .A3(\input [3]), .A4(
        \input [31]), .ZN(n9) );
  NOR4_X1 U5 ( .A1(\input [30]), .A2(\input [2]), .A3(\input [29]), .A4(
        \input [28]), .ZN(n8) );
  NOR4_X1 U6 ( .A1(\input [16]), .A2(\input [15]), .A3(\input [14]), .A4(
        \input [13]), .ZN(n4) );
  NOR4_X1 U7 ( .A1(\input [27]), .A2(\input [26]), .A3(\input [25]), .A4(
        \input [24]), .ZN(n7) );
  NOR2_X1 U8 ( .A1(n1), .A2(n2), .ZN(result) );
  NAND4_X1 U9 ( .A1(n3), .A2(n4), .A3(n5), .A4(n6), .ZN(n2) );
  NAND4_X1 U10 ( .A1(n7), .A2(n8), .A3(n9), .A4(n10), .ZN(n1) );
  NOR4_X1 U11 ( .A1(\input [12]), .A2(\input [11]), .A3(\input [10]), .A4(
        \input [0]), .ZN(n3) );
endmodule


module comparator ( Z, cout, eq, neq, gt, lt, ge, le );
  input Z, cout;
  output eq, neq, gt, lt, ge, le;
  wire   Z, cout;
  assign eq = Z;
  assign ge = cout;

  INV_X1 U1 ( .A(le), .ZN(gt) );
  INV_X1 U2 ( .A(cout), .ZN(lt) );
  NAND2_X1 U3 ( .A1(cout), .A2(neq), .ZN(le) );
  INV_X1 U4 ( .A(Z), .ZN(neq) );
endmodule


module ALU_N32 ( DATA1, DATA2, FUNC, SN, OVF, OUTALU );
  input [31:0] DATA1;
  input [31:0] DATA2;
  input [3:0] FUNC;
  output [31:0] OUTALU;
  input SN;
  output OVF;
  wire   s_LnR, s_AnL, s_RnS, p4_cin, p4_cout, p4_ovf, is_zero, s_eq, s_neq,
         s_gt, s_lt, N74, N75, N76, N77, N78, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n42, n43, n100, n101, n102, n103, n104, n105, n106, n107
;
  wire   [31:0] shifter_out;
  wire   [31:0] p4_sum;
  wire   [3:0] logic_func;
  wire   [31:0] logic_out;

  DLH_X1 s_RnS_reg ( .G(n3), .D(n97), .Q(s_RnS) );
  DLH_X1 p4_cin_reg ( .G(N74), .D(N75), .Q(p4_cin) );
  DLH_X1 OVF_reg ( .G(n9), .D(p4_ovf), .Q(OVF) );
  DLH_X1 \logic_func_reg[3]  ( .G(n6), .D(FUNC[3]), .Q(logic_func[3]) );
  DLH_X1 \logic_func_reg[2]  ( .G(n6), .D(FUNC[2]), .Q(logic_func[2]) );
  DLH_X1 \logic_func_reg[1]  ( .G(n6), .D(FUNC[1]), .Q(logic_func[1]) );
  DLH_X1 \logic_func_reg[0]  ( .G(n6), .D(FUNC[0]), .Q(logic_func[0]) );
  DLH_X1 s_LnR_reg ( .G(n3), .D(n98), .Q(s_LnR) );
  DLH_X1 s_AnL_reg ( .G(n3), .D(n99), .Q(s_AnL) );
  NAND3_X1 U102 ( .A1(n78), .A2(n79), .A3(n80), .ZN(OUTALU[0]) );
  XOR2_X1 U103 ( .A(DATA2[31]), .B(n10), .Z(n94) );
  NAND3_X1 U104 ( .A1(FUNC[1]), .A2(n107), .A3(FUNC[2]), .ZN(n44) );
  OAI33_X1 U105 ( .A1(n106), .A2(FUNC[3]), .A3(FUNC[2]), .B1(n46), .B2(FUNC[1]), .B3(FUNC[0]), .ZN(N77) );
  NAND3_X1 U106 ( .A1(FUNC[3]), .A2(FUNC[2]), .A3(n105), .ZN(n88) );
  shifter_NBITS32 alu_shifter ( .R1({n10, DATA1[30:0]}), .R2(DATA2), .LnR(
        s_LnR), .AnL(s_AnL), .RnS(s_RnS), .Rout(shifter_out) );
  P4_ADDER_NBIT32_1 alu_adder ( .A({n10, DATA1[30:0]}), .B(DATA2), .Cin(p4_cin), .S(p4_sum), .Cout(p4_cout), .ovf(p4_ovf) );
  logicals_nbit32 alu_logicals ( .func(logic_func), .SN(SN), .in1({n10, 
        DATA1[30:0]}), .in2(DATA2), .o(logic_out) );
  nor_generic_NBITS32 nor_gen ( .\input (p4_sum), .result(is_zero) );
  comparator comp ( .Z(is_zero), .cout(p4_cout), .eq(s_eq), .neq(s_neq), .gt(
        s_gt), .lt(s_lt) );
  INV_X1 U2 ( .A(n64), .ZN(OUTALU[22]) );
  AOI222_X1 U3 ( .A1(shifter_out[22]), .A2(n2), .B1(p4_sum[22]), .B2(n8), .C1(
        logic_out[22]), .C2(n5), .ZN(n64) );
  INV_X1 U4 ( .A(n65), .ZN(OUTALU[21]) );
  AOI222_X1 U5 ( .A1(shifter_out[21]), .A2(n2), .B1(p4_sum[21]), .B2(n8), .C1(
        logic_out[21]), .C2(n5), .ZN(n65) );
  INV_X1 U6 ( .A(n68), .ZN(OUTALU[19]) );
  AOI222_X1 U7 ( .A1(shifter_out[19]), .A2(n2), .B1(p4_sum[19]), .B2(n8), .C1(
        logic_out[19]), .C2(n5), .ZN(n68) );
  INV_X1 U8 ( .A(n72), .ZN(OUTALU[15]) );
  AOI222_X1 U9 ( .A1(shifter_out[15]), .A2(n3), .B1(p4_sum[15]), .B2(n9), .C1(
        logic_out[15]), .C2(n6), .ZN(n72) );
  INV_X1 U10 ( .A(n73), .ZN(OUTALU[14]) );
  AOI222_X1 U11 ( .A1(shifter_out[14]), .A2(n3), .B1(p4_sum[14]), .B2(n9), 
        .C1(logic_out[14]), .C2(n6), .ZN(n73) );
  INV_X1 U12 ( .A(n74), .ZN(OUTALU[13]) );
  AOI222_X1 U13 ( .A1(shifter_out[13]), .A2(n3), .B1(p4_sum[13]), .B2(n9), 
        .C1(logic_out[13]), .C2(n6), .ZN(n74) );
  INV_X1 U14 ( .A(n76), .ZN(OUTALU[11]) );
  AOI222_X1 U15 ( .A1(shifter_out[11]), .A2(n3), .B1(p4_sum[11]), .B2(n9), 
        .C1(logic_out[11]), .C2(n6), .ZN(n76) );
  INV_X1 U16 ( .A(n77), .ZN(OUTALU[10]) );
  AOI222_X1 U17 ( .A1(shifter_out[10]), .A2(n3), .B1(p4_sum[10]), .B2(n9), 
        .C1(logic_out[10]), .C2(n6), .ZN(n77) );
  INV_X1 U18 ( .A(n54), .ZN(OUTALU[31]) );
  AOI222_X1 U19 ( .A1(shifter_out[31]), .A2(n1), .B1(p4_sum[31]), .B2(n7), 
        .C1(logic_out[31]), .C2(n4), .ZN(n54) );
  INV_X1 U20 ( .A(n55), .ZN(OUTALU[30]) );
  AOI222_X1 U21 ( .A1(shifter_out[30]), .A2(n1), .B1(p4_sum[30]), .B2(n7), 
        .C1(logic_out[30]), .C2(n4), .ZN(n55) );
  INV_X1 U22 ( .A(n57), .ZN(OUTALU[29]) );
  AOI222_X1 U23 ( .A1(shifter_out[29]), .A2(n1), .B1(p4_sum[29]), .B2(n7), 
        .C1(logic_out[29]), .C2(n4), .ZN(n57) );
  INV_X1 U24 ( .A(n59), .ZN(OUTALU[27]) );
  AOI222_X1 U25 ( .A1(shifter_out[27]), .A2(n2), .B1(p4_sum[27]), .B2(n8), 
        .C1(logic_out[27]), .C2(n5), .ZN(n59) );
  INV_X1 U26 ( .A(n60), .ZN(OUTALU[26]) );
  AOI222_X1 U27 ( .A1(shifter_out[26]), .A2(n2), .B1(p4_sum[26]), .B2(n8), 
        .C1(logic_out[26]), .C2(n5), .ZN(n60) );
  INV_X1 U28 ( .A(n61), .ZN(OUTALU[25]) );
  AOI222_X1 U29 ( .A1(shifter_out[25]), .A2(n2), .B1(p4_sum[25]), .B2(n8), 
        .C1(logic_out[25]), .C2(n5), .ZN(n61) );
  INV_X1 U30 ( .A(n63), .ZN(OUTALU[23]) );
  AOI222_X1 U31 ( .A1(shifter_out[23]), .A2(n2), .B1(p4_sum[23]), .B2(n8), 
        .C1(logic_out[23]), .C2(n5), .ZN(n63) );
  INV_X1 U32 ( .A(n69), .ZN(OUTALU[18]) );
  AOI222_X1 U33 ( .A1(shifter_out[18]), .A2(n2), .B1(p4_sum[18]), .B2(n8), 
        .C1(logic_out[18]), .C2(n5), .ZN(n69) );
  INV_X1 U34 ( .A(n47), .ZN(OUTALU[9]) );
  AOI222_X1 U35 ( .A1(shifter_out[9]), .A2(n2), .B1(p4_sum[9]), .B2(n8), .C1(
        logic_out[9]), .C2(n5), .ZN(n47) );
  INV_X1 U36 ( .A(n49), .ZN(OUTALU[7]) );
  AOI222_X1 U37 ( .A1(shifter_out[7]), .A2(n1), .B1(p4_sum[7]), .B2(n7), .C1(
        logic_out[7]), .C2(n4), .ZN(n49) );
  INV_X1 U38 ( .A(n50), .ZN(OUTALU[6]) );
  AOI222_X1 U39 ( .A1(shifter_out[6]), .A2(n1), .B1(p4_sum[6]), .B2(n7), .C1(
        logic_out[6]), .C2(n4), .ZN(n50) );
  INV_X1 U40 ( .A(n51), .ZN(OUTALU[5]) );
  AOI222_X1 U41 ( .A1(shifter_out[5]), .A2(n1), .B1(p4_sum[5]), .B2(n7), .C1(
        logic_out[5]), .C2(n4), .ZN(n51) );
  INV_X1 U42 ( .A(n53), .ZN(OUTALU[3]) );
  AOI222_X1 U43 ( .A1(shifter_out[3]), .A2(n1), .B1(p4_sum[3]), .B2(n7), .C1(
        logic_out[3]), .C2(n4), .ZN(n53) );
  INV_X1 U44 ( .A(n56), .ZN(OUTALU[2]) );
  AOI222_X1 U45 ( .A1(shifter_out[2]), .A2(n1), .B1(p4_sum[2]), .B2(n7), .C1(
        logic_out[2]), .C2(n4), .ZN(n56) );
  INV_X1 U46 ( .A(n67), .ZN(OUTALU[1]) );
  AOI222_X1 U47 ( .A1(shifter_out[1]), .A2(n2), .B1(p4_sum[1]), .B2(n8), .C1(
        logic_out[1]), .C2(n5), .ZN(n67) );
  INV_X1 U48 ( .A(n70), .ZN(OUTALU[17]) );
  AOI222_X1 U49 ( .A1(shifter_out[17]), .A2(n3), .B1(p4_sum[17]), .B2(n9), 
        .C1(logic_out[17]), .C2(n6), .ZN(n70) );
  BUF_X1 U50 ( .A(N78), .Z(n1) );
  BUF_X1 U51 ( .A(N78), .Z(n2) );
  BUF_X1 U52 ( .A(N78), .Z(n3) );
  INV_X1 U53 ( .A(n93), .ZN(n100) );
  OR2_X1 U54 ( .A1(n9), .A2(N75), .ZN(N74) );
  INV_X1 U55 ( .A(n62), .ZN(OUTALU[24]) );
  AOI222_X1 U56 ( .A1(shifter_out[24]), .A2(n2), .B1(p4_sum[24]), .B2(n8), 
        .C1(logic_out[24]), .C2(n5), .ZN(n62) );
  INV_X1 U57 ( .A(n66), .ZN(OUTALU[20]) );
  AOI222_X1 U58 ( .A1(shifter_out[20]), .A2(n2), .B1(p4_sum[20]), .B2(n8), 
        .C1(logic_out[20]), .C2(n5), .ZN(n66) );
  INV_X1 U59 ( .A(n71), .ZN(OUTALU[16]) );
  AOI222_X1 U60 ( .A1(shifter_out[16]), .A2(n3), .B1(p4_sum[16]), .B2(n9), 
        .C1(logic_out[16]), .C2(n6), .ZN(n71) );
  INV_X1 U61 ( .A(n75), .ZN(OUTALU[12]) );
  AOI222_X1 U62 ( .A1(shifter_out[12]), .A2(n3), .B1(p4_sum[12]), .B2(n9), 
        .C1(logic_out[12]), .C2(n6), .ZN(n75) );
  OAI222_X1 U63 ( .A1(s_lt), .A2(n88), .B1(s_eq), .B2(n90), .C1(s_gt), .C2(n91), .ZN(n81) );
  AOI22_X1 U64 ( .A1(n92), .A2(s_gt), .B1(n93), .B2(s_lt), .ZN(n90) );
  BUF_X1 U65 ( .A(DATA1[31]), .Z(n10) );
  OAI21_X1 U66 ( .B1(n42), .B2(n84), .A(n85), .ZN(n83) );
  OAI21_X1 U67 ( .B1(s_eq), .B2(n86), .A(n87), .ZN(n85) );
  AOI22_X1 U68 ( .A1(s_lt), .A2(n103), .B1(s_gt), .B2(n102), .ZN(n84) );
  OAI22_X1 U69 ( .A1(n100), .A2(s_lt), .B1(n101), .B2(s_gt), .ZN(n87) );
  AOI22_X1 U70 ( .A1(logic_out[0]), .A2(n4), .B1(shifter_out[0]), .B2(n1), 
        .ZN(n78) );
  AOI22_X1 U71 ( .A1(s_eq), .A2(n95), .B1(p4_sum[0]), .B2(n7), .ZN(n79) );
  AOI221_X1 U72 ( .B1(n42), .B2(n81), .C1(n82), .C2(s_neq), .A(n83), .ZN(n80)
         );
  INV_X1 U73 ( .A(n58), .ZN(OUTALU[28]) );
  AOI222_X1 U74 ( .A1(shifter_out[28]), .A2(n1), .B1(p4_sum[28]), .B2(n7), 
        .C1(logic_out[28]), .C2(n4), .ZN(n58) );
  INV_X1 U75 ( .A(n48), .ZN(OUTALU[8]) );
  AOI222_X1 U76 ( .A1(shifter_out[8]), .A2(n1), .B1(p4_sum[8]), .B2(n7), .C1(
        logic_out[8]), .C2(n4), .ZN(n48) );
  INV_X1 U77 ( .A(n52), .ZN(OUTALU[4]) );
  AOI222_X1 U78 ( .A1(shifter_out[4]), .A2(n1), .B1(p4_sum[4]), .B2(n7), .C1(
        logic_out[4]), .C2(n4), .ZN(n52) );
  INV_X1 U79 ( .A(n86), .ZN(n42) );
  BUF_X1 U80 ( .A(N76), .Z(n7) );
  BUF_X1 U81 ( .A(N76), .Z(n8) );
  NOR3_X1 U82 ( .A1(n107), .A2(n106), .A3(n89), .ZN(n93) );
  BUF_X1 U83 ( .A(N77), .Z(n6) );
  BUF_X1 U84 ( .A(N76), .Z(n9) );
  BUF_X1 U85 ( .A(N77), .Z(n4) );
  BUF_X1 U86 ( .A(N77), .Z(n5) );
  OAI21_X1 U87 ( .B1(n107), .B2(n46), .A(n44), .ZN(N78) );
  NOR2_X1 U88 ( .A1(n45), .A2(n89), .ZN(n82) );
  INV_X1 U89 ( .A(n91), .ZN(n102) );
  INV_X1 U90 ( .A(n88), .ZN(n103) );
  INV_X1 U91 ( .A(n92), .ZN(n101) );
  INV_X1 U92 ( .A(n45), .ZN(n105) );
  NOR3_X1 U93 ( .A1(n46), .A2(n106), .A3(n107), .ZN(n99) );
  NAND4_X1 U94 ( .A1(n100), .A2(n88), .A3(n101), .A4(n96), .ZN(N75) );
  AOI211_X1 U95 ( .C1(n105), .C2(n104), .A(n102), .B(n95), .ZN(n96) );
  NOR2_X1 U96 ( .A1(n44), .A2(n43), .ZN(n97) );
  NOR2_X1 U97 ( .A1(n45), .A2(n46), .ZN(n98) );
  NAND2_X1 U98 ( .A1(SN), .A2(n94), .ZN(n86) );
  NOR3_X1 U99 ( .A1(FUNC[0]), .A2(FUNC[1]), .A3(n89), .ZN(n95) );
  NOR3_X1 U100 ( .A1(n106), .A2(FUNC[0]), .A3(n89), .ZN(n92) );
  NOR3_X1 U101 ( .A1(FUNC[2]), .A2(FUNC[3]), .A3(FUNC[1]), .ZN(N76) );
  NAND4_X1 U107 ( .A1(FUNC[3]), .A2(FUNC[2]), .A3(n107), .A4(n106), .ZN(n91)
         );
  INV_X1 U108 ( .A(FUNC[1]), .ZN(n106) );
  NAND2_X1 U109 ( .A1(FUNC[2]), .A2(n43), .ZN(n46) );
  NAND2_X1 U110 ( .A1(FUNC[3]), .A2(n104), .ZN(n89) );
  NAND2_X1 U111 ( .A1(FUNC[0]), .A2(n106), .ZN(n45) );
  INV_X1 U112 ( .A(FUNC[0]), .ZN(n107) );
  INV_X1 U113 ( .A(FUNC[2]), .ZN(n104) );
  INV_X1 U114 ( .A(FUNC[3]), .ZN(n43) );
endmodule


module enc33_0 ( A, Y );
  input [2:0] A;
  output [2:0] Y;
  wire   n3, n4, n5, n1, n2;

  XOR2_X1 U8 ( .A(A[0]), .B(A[1]), .Z(n4) );
  OAI21_X1 U1 ( .B1(n2), .B2(n1), .A(n5), .ZN(Y[1]) );
  NOR3_X1 U2 ( .A1(n1), .A2(n3), .A3(n4), .ZN(Y[2]) );
  OAI21_X1 U3 ( .B1(A[2]), .B2(n2), .A(n5), .ZN(Y[0]) );
  INV_X1 U4 ( .A(n4), .ZN(n2) );
  NAND2_X1 U5 ( .A1(n3), .A2(n1), .ZN(n5) );
  AND2_X1 U6 ( .A1(A[1]), .A2(A[0]), .ZN(n3) );
  INV_X1 U7 ( .A(A[2]), .ZN(n1) );
endmodule


module enc33_3 ( A, Y );
  input [2:0] A;
  output [2:0] Y;
  wire   n1, n2, n7, n8, n9;

  XOR2_X1 U8 ( .A(A[0]), .B(A[1]), .Z(n8) );
  NOR3_X1 U1 ( .A1(n1), .A2(n9), .A3(n8), .ZN(Y[2]) );
  OAI21_X1 U2 ( .B1(n2), .B2(n1), .A(n7), .ZN(Y[1]) );
  NAND2_X1 U3 ( .A1(n9), .A2(n1), .ZN(n7) );
  INV_X1 U4 ( .A(n8), .ZN(n2) );
  OAI21_X1 U5 ( .B1(A[2]), .B2(n2), .A(n7), .ZN(Y[0]) );
  AND2_X1 U6 ( .A1(A[1]), .A2(A[0]), .ZN(n9) );
  INV_X1 U7 ( .A(A[2]), .ZN(n1) );
endmodule


module enc33_2 ( A, Y );
  input [2:0] A;
  output [2:0] Y;
  wire   n1, n2, n7, n8, n9;

  XOR2_X1 U8 ( .A(A[0]), .B(A[1]), .Z(n8) );
  NOR3_X1 U1 ( .A1(n2), .A2(n9), .A3(n8), .ZN(Y[2]) );
  INV_X1 U2 ( .A(n8), .ZN(n1) );
  NAND2_X1 U3 ( .A1(n9), .A2(n2), .ZN(n7) );
  OAI21_X1 U4 ( .B1(n1), .B2(n2), .A(n7), .ZN(Y[1]) );
  INV_X1 U5 ( .A(A[2]), .ZN(n2) );
  OAI21_X1 U6 ( .B1(A[2]), .B2(n1), .A(n7), .ZN(Y[0]) );
  AND2_X1 U7 ( .A1(A[1]), .A2(A[0]), .ZN(n9) );
endmodule


module enc33_1 ( A, Y );
  input [2:0] A;
  output [2:0] Y;
  wire   n1, n2, n7, n8, n9;

  XOR2_X1 U8 ( .A(A[0]), .B(A[1]), .Z(n8) );
  NOR3_X1 U1 ( .A1(n2), .A2(n9), .A3(n8), .ZN(Y[2]) );
  INV_X1 U2 ( .A(n8), .ZN(n1) );
  OAI21_X1 U3 ( .B1(n1), .B2(n2), .A(n7), .ZN(Y[1]) );
  NAND2_X1 U4 ( .A1(n9), .A2(n2), .ZN(n7) );
  INV_X1 U5 ( .A(A[2]), .ZN(n2) );
  OAI21_X1 U6 ( .B1(A[2]), .B2(n1), .A(n7), .ZN(Y[0]) );
  AND2_X1 U7 ( .A1(A[1]), .A2(A[0]), .ZN(n9) );
endmodule


module shl1_NBIT32_0 ( A, Y );
  input [31:0] A;
  output [31:0] Y;
  wire   \A[30] , \A[29] , \A[28] , \A[27] , \A[26] , \A[25] , \A[24] ,
         \A[23] , \A[22] , \A[21] , \A[20] , \A[19] , \A[18] , \A[17] ,
         \A[16] , \A[15] , \A[14] , \A[13] , \A[12] , \A[11] , \A[10] , \A[9] ,
         \A[8] , \A[7] , \A[6] , \A[5] , \A[4] , \A[3] , \A[2] , \A[1] ,
         \A[0] ;
  assign Y[0] = 1'b0;
  assign Y[31] = \A[30] ;
  assign \A[30]  = A[30];
  assign Y[30] = \A[29] ;
  assign \A[29]  = A[29];
  assign Y[29] = \A[28] ;
  assign \A[28]  = A[28];
  assign Y[28] = \A[27] ;
  assign \A[27]  = A[27];
  assign Y[27] = \A[26] ;
  assign \A[26]  = A[26];
  assign Y[26] = \A[25] ;
  assign \A[25]  = A[25];
  assign Y[25] = \A[24] ;
  assign \A[24]  = A[24];
  assign Y[24] = \A[23] ;
  assign \A[23]  = A[23];
  assign Y[23] = \A[22] ;
  assign \A[22]  = A[22];
  assign Y[22] = \A[21] ;
  assign \A[21]  = A[21];
  assign Y[21] = \A[20] ;
  assign \A[20]  = A[20];
  assign Y[20] = \A[19] ;
  assign \A[19]  = A[19];
  assign Y[19] = \A[18] ;
  assign \A[18]  = A[18];
  assign Y[18] = \A[17] ;
  assign \A[17]  = A[17];
  assign Y[17] = \A[16] ;
  assign \A[16]  = A[16];
  assign Y[16] = \A[15] ;
  assign \A[15]  = A[15];
  assign Y[15] = \A[14] ;
  assign \A[14]  = A[14];
  assign Y[14] = \A[13] ;
  assign \A[13]  = A[13];
  assign Y[13] = \A[12] ;
  assign \A[12]  = A[12];
  assign Y[12] = \A[11] ;
  assign \A[11]  = A[11];
  assign Y[11] = \A[10] ;
  assign \A[10]  = A[10];
  assign Y[10] = \A[9] ;
  assign \A[9]  = A[9];
  assign Y[9] = \A[8] ;
  assign \A[8]  = A[8];
  assign Y[8] = \A[7] ;
  assign \A[7]  = A[7];
  assign Y[7] = \A[6] ;
  assign \A[6]  = A[6];
  assign Y[6] = \A[5] ;
  assign \A[5]  = A[5];
  assign Y[5] = \A[4] ;
  assign \A[4]  = A[4];
  assign Y[4] = \A[3] ;
  assign \A[3]  = A[3];
  assign Y[3] = \A[2] ;
  assign \A[2]  = A[2];
  assign Y[2] = \A[1] ;
  assign \A[1]  = A[1];
  assign Y[1] = \A[0] ;
  assign \A[0]  = A[0];

endmodule


module shl2_NBIT32_0 ( A, Y );
  input [31:0] A;
  output [31:0] Y;
  wire   \A[29] , \A[28] , \A[27] , \A[26] , \A[25] , \A[24] , \A[23] ,
         \A[22] , \A[21] , \A[20] , \A[19] , \A[18] , \A[17] , \A[16] ,
         \A[15] , \A[14] , \A[13] , \A[12] , \A[11] , \A[10] , \A[9] , \A[8] ,
         \A[7] , \A[6] , \A[5] , \A[4] , \A[3] , \A[2] , \A[1] , \A[0] ;
  assign Y[0] = 1'b0;
  assign Y[1] = 1'b0;
  assign Y[31] = \A[29] ;
  assign \A[29]  = A[29];
  assign Y[30] = \A[28] ;
  assign \A[28]  = A[28];
  assign Y[29] = \A[27] ;
  assign \A[27]  = A[27];
  assign Y[28] = \A[26] ;
  assign \A[26]  = A[26];
  assign Y[27] = \A[25] ;
  assign \A[25]  = A[25];
  assign Y[26] = \A[24] ;
  assign \A[24]  = A[24];
  assign Y[25] = \A[23] ;
  assign \A[23]  = A[23];
  assign Y[24] = \A[22] ;
  assign \A[22]  = A[22];
  assign Y[23] = \A[21] ;
  assign \A[21]  = A[21];
  assign Y[22] = \A[20] ;
  assign \A[20]  = A[20];
  assign Y[21] = \A[19] ;
  assign \A[19]  = A[19];
  assign Y[20] = \A[18] ;
  assign \A[18]  = A[18];
  assign Y[19] = \A[17] ;
  assign \A[17]  = A[17];
  assign Y[18] = \A[16] ;
  assign \A[16]  = A[16];
  assign Y[17] = \A[15] ;
  assign \A[15]  = A[15];
  assign Y[16] = \A[14] ;
  assign \A[14]  = A[14];
  assign Y[15] = \A[13] ;
  assign \A[13]  = A[13];
  assign Y[14] = \A[12] ;
  assign \A[12]  = A[12];
  assign Y[13] = \A[11] ;
  assign \A[11]  = A[11];
  assign Y[12] = \A[10] ;
  assign \A[10]  = A[10];
  assign Y[11] = \A[9] ;
  assign \A[9]  = A[9];
  assign Y[10] = \A[8] ;
  assign \A[8]  = A[8];
  assign Y[9] = \A[7] ;
  assign \A[7]  = A[7];
  assign Y[8] = \A[6] ;
  assign \A[6]  = A[6];
  assign Y[7] = \A[5] ;
  assign \A[5]  = A[5];
  assign Y[6] = \A[4] ;
  assign \A[4]  = A[4];
  assign Y[5] = \A[3] ;
  assign \A[3]  = A[3];
  assign Y[4] = \A[2] ;
  assign \A[2]  = A[2];
  assign Y[3] = \A[1] ;
  assign \A[1]  = A[1];
  assign Y[2] = \A[0] ;
  assign \A[0]  = A[0];

endmodule


module shl3_NBIT32 ( A, Y );
  input [31:0] A;
  output [31:0] Y;
  wire   \A[28] , \A[27] , \A[26] , \A[25] , \A[24] , \A[23] , \A[22] ,
         \A[21] , \A[20] , \A[19] , \A[18] , \A[17] , \A[16] , \A[15] ,
         \A[14] , \A[13] , \A[12] , \A[11] , \A[10] , \A[9] , \A[8] , \A[7] ,
         \A[6] , \A[5] , \A[4] , \A[3] , \A[2] , \A[1] , \A[0] ;
  assign Y[0] = 1'b0;
  assign Y[1] = 1'b0;
  assign Y[2] = 1'b0;
  assign Y[31] = \A[28] ;
  assign \A[28]  = A[28];
  assign Y[30] = \A[27] ;
  assign \A[27]  = A[27];
  assign Y[29] = \A[26] ;
  assign \A[26]  = A[26];
  assign Y[28] = \A[25] ;
  assign \A[25]  = A[25];
  assign Y[27] = \A[24] ;
  assign \A[24]  = A[24];
  assign Y[26] = \A[23] ;
  assign \A[23]  = A[23];
  assign Y[25] = \A[22] ;
  assign \A[22]  = A[22];
  assign Y[24] = \A[21] ;
  assign \A[21]  = A[21];
  assign Y[23] = \A[20] ;
  assign \A[20]  = A[20];
  assign Y[22] = \A[19] ;
  assign \A[19]  = A[19];
  assign Y[21] = \A[18] ;
  assign \A[18]  = A[18];
  assign Y[20] = \A[17] ;
  assign \A[17]  = A[17];
  assign Y[19] = \A[16] ;
  assign \A[16]  = A[16];
  assign Y[18] = \A[15] ;
  assign \A[15]  = A[15];
  assign Y[17] = \A[14] ;
  assign \A[14]  = A[14];
  assign Y[16] = \A[13] ;
  assign \A[13]  = A[13];
  assign Y[15] = \A[12] ;
  assign \A[12]  = A[12];
  assign Y[14] = \A[11] ;
  assign \A[11]  = A[11];
  assign Y[13] = \A[10] ;
  assign \A[10]  = A[10];
  assign Y[12] = \A[9] ;
  assign \A[9]  = A[9];
  assign Y[11] = \A[8] ;
  assign \A[8]  = A[8];
  assign Y[10] = \A[7] ;
  assign \A[7]  = A[7];
  assign Y[9] = \A[6] ;
  assign \A[6]  = A[6];
  assign Y[8] = \A[5] ;
  assign \A[5]  = A[5];
  assign Y[7] = \A[4] ;
  assign \A[4]  = A[4];
  assign Y[6] = \A[3] ;
  assign \A[3]  = A[3];
  assign Y[5] = \A[2] ;
  assign \A[2]  = A[2];
  assign Y[4] = \A[1] ;
  assign \A[1]  = A[1];
  assign Y[3] = \A[0] ;
  assign \A[0]  = A[0];

endmodule


module negate_NBIT32_0_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U1 ( .A(n63), .B(n7), .Z(DIFF[2]) );
  XOR2_X1 U2 ( .A(n64), .B(n8), .Z(DIFF[3]) );
  XOR2_X1 U3 ( .A(n65), .B(n9), .Z(DIFF[4]) );
  XOR2_X1 U4 ( .A(n62), .B(n92), .Z(DIFF[1]) );
  AND2_X1 U5 ( .A1(n73), .A2(n22), .ZN(n5) );
  AND2_X1 U6 ( .A1(n74), .A2(n5), .ZN(n6) );
  AND2_X1 U7 ( .A1(n62), .A2(n92), .ZN(n7) );
  AND2_X1 U8 ( .A1(n63), .A2(n7), .ZN(n8) );
  AND2_X1 U9 ( .A1(n64), .A2(n8), .ZN(n9) );
  AND2_X1 U10 ( .A1(n65), .A2(n9), .ZN(n10) );
  AND2_X1 U11 ( .A1(n66), .A2(n10), .ZN(n11) );
  AND2_X1 U12 ( .A1(n67), .A2(n11), .ZN(n12) );
  AND2_X1 U13 ( .A1(n68), .A2(n12), .ZN(n13) );
  AND2_X1 U14 ( .A1(n85), .A2(n32), .ZN(n14) );
  AND2_X1 U15 ( .A1(n86), .A2(n14), .ZN(n15) );
  AND2_X1 U16 ( .A1(n87), .A2(n15), .ZN(n16) );
  AND2_X1 U17 ( .A1(n88), .A2(n16), .ZN(n17) );
  AND2_X1 U18 ( .A1(n89), .A2(n17), .ZN(n18) );
  AND2_X1 U19 ( .A1(n69), .A2(n13), .ZN(n19) );
  AND2_X1 U20 ( .A1(n70), .A2(n19), .ZN(n20) );
  AND2_X1 U21 ( .A1(n71), .A2(n20), .ZN(n21) );
  AND2_X1 U22 ( .A1(n72), .A2(n21), .ZN(n22) );
  AND2_X1 U23 ( .A1(n75), .A2(n6), .ZN(n23) );
  AND2_X1 U24 ( .A1(n76), .A2(n23), .ZN(n24) );
  AND2_X1 U25 ( .A1(n77), .A2(n24), .ZN(n25) );
  AND2_X1 U26 ( .A1(n78), .A2(n25), .ZN(n26) );
  AND2_X1 U27 ( .A1(n79), .A2(n26), .ZN(n27) );
  AND2_X1 U28 ( .A1(n80), .A2(n27), .ZN(n28) );
  AND2_X1 U29 ( .A1(n81), .A2(n28), .ZN(n29) );
  AND2_X1 U30 ( .A1(n82), .A2(n29), .ZN(n30) );
  AND2_X1 U31 ( .A1(n83), .A2(n30), .ZN(n31) );
  AND2_X1 U32 ( .A1(n84), .A2(n31), .ZN(n32) );
  AND2_X1 U33 ( .A1(n90), .A2(n18), .ZN(n33) );
  NAND2_X1 U34 ( .A1(n91), .A2(n33), .ZN(n61) );
  XOR2_X1 U35 ( .A(n85), .B(n32), .Z(DIFF[24]) );
  XOR2_X1 U36 ( .A(n86), .B(n14), .Z(DIFF[25]) );
  XOR2_X1 U37 ( .A(n87), .B(n15), .Z(DIFF[26]) );
  XOR2_X1 U38 ( .A(n88), .B(n16), .Z(DIFF[27]) );
  XOR2_X1 U39 ( .A(n89), .B(n17), .Z(DIFF[28]) );
  XOR2_X1 U40 ( .A(n84), .B(n31), .Z(DIFF[23]) );
  XOR2_X1 U41 ( .A(n90), .B(n18), .Z(DIFF[29]) );
  XOR2_X1 U42 ( .A(n91), .B(n33), .Z(DIFF[30]) );
  XOR2_X1 U43 ( .A(B[31]), .B(n61), .Z(DIFF[31]) );
  XOR2_X1 U44 ( .A(n73), .B(n22), .Z(DIFF[12]) );
  XOR2_X1 U45 ( .A(n74), .B(n5), .Z(DIFF[13]) );
  XOR2_X1 U46 ( .A(n75), .B(n6), .Z(DIFF[14]) );
  XOR2_X1 U47 ( .A(n76), .B(n23), .Z(DIFF[15]) );
  XOR2_X1 U48 ( .A(n77), .B(n24), .Z(DIFF[16]) );
  XOR2_X1 U49 ( .A(n78), .B(n25), .Z(DIFF[17]) );
  XOR2_X1 U50 ( .A(n79), .B(n26), .Z(DIFF[18]) );
  XOR2_X1 U51 ( .A(n80), .B(n27), .Z(DIFF[19]) );
  XOR2_X1 U52 ( .A(n81), .B(n28), .Z(DIFF[20]) );
  XOR2_X1 U53 ( .A(n82), .B(n29), .Z(DIFF[21]) );
  XOR2_X1 U54 ( .A(n83), .B(n30), .Z(DIFF[22]) );
  XOR2_X1 U55 ( .A(n66), .B(n10), .Z(DIFF[5]) );
  XOR2_X1 U56 ( .A(n67), .B(n11), .Z(DIFF[6]) );
  XOR2_X1 U57 ( .A(n68), .B(n12), .Z(DIFF[7]) );
  XOR2_X1 U58 ( .A(n69), .B(n13), .Z(DIFF[8]) );
  XOR2_X1 U59 ( .A(n70), .B(n19), .Z(DIFF[9]) );
  XOR2_X1 U60 ( .A(n71), .B(n20), .Z(DIFF[10]) );
  XOR2_X1 U61 ( .A(n72), .B(n21), .Z(DIFF[11]) );
  INV_X1 U62 ( .A(\B[0] ), .ZN(n92) );
  INV_X1 U63 ( .A(B[1]), .ZN(n62) );
  INV_X1 U64 ( .A(B[2]), .ZN(n63) );
  INV_X1 U65 ( .A(B[3]), .ZN(n64) );
  INV_X1 U66 ( .A(B[4]), .ZN(n65) );
  INV_X1 U67 ( .A(B[5]), .ZN(n66) );
  INV_X1 U68 ( .A(B[6]), .ZN(n67) );
  INV_X1 U69 ( .A(B[7]), .ZN(n68) );
  INV_X1 U70 ( .A(B[8]), .ZN(n69) );
  INV_X1 U71 ( .A(B[9]), .ZN(n70) );
  INV_X1 U72 ( .A(B[10]), .ZN(n71) );
  INV_X1 U73 ( .A(B[11]), .ZN(n72) );
  INV_X1 U74 ( .A(B[12]), .ZN(n73) );
  INV_X1 U75 ( .A(B[13]), .ZN(n74) );
  INV_X1 U76 ( .A(B[14]), .ZN(n75) );
  INV_X1 U77 ( .A(B[15]), .ZN(n76) );
  INV_X1 U78 ( .A(B[16]), .ZN(n77) );
  INV_X1 U79 ( .A(B[17]), .ZN(n78) );
  INV_X1 U80 ( .A(B[18]), .ZN(n79) );
  INV_X1 U81 ( .A(B[19]), .ZN(n80) );
  INV_X1 U82 ( .A(B[20]), .ZN(n81) );
  INV_X1 U83 ( .A(B[24]), .ZN(n85) );
  INV_X1 U84 ( .A(B[25]), .ZN(n86) );
  INV_X1 U85 ( .A(B[26]), .ZN(n87) );
  INV_X1 U86 ( .A(B[27]), .ZN(n88) );
  INV_X1 U87 ( .A(B[28]), .ZN(n89) );
  INV_X1 U88 ( .A(B[21]), .ZN(n82) );
  INV_X1 U89 ( .A(B[22]), .ZN(n83) );
  INV_X1 U90 ( .A(B[23]), .ZN(n84) );
  INV_X1 U91 ( .A(B[29]), .ZN(n90) );
  INV_X1 U92 ( .A(B[30]), .ZN(n91) );
endmodule


module negate_NBIT32_0 ( A, Y );
  input [31:0] A;
  output [31:0] Y;


  negate_NBIT32_0_DW01_sub_0 sub_add_14_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .B(A), .CI(1'b0), .DIFF(Y) );
endmodule


module negate_NBIT32_7_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n59, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U1 ( .A(B[31]), .B(n61), .Z(DIFF[31]) );
  XOR2_X1 U2 ( .A(n91), .B(n41), .Z(DIFF[30]) );
  XOR2_X1 U3 ( .A(n84), .B(n53), .Z(DIFF[23]) );
  XOR2_X1 U4 ( .A(n85), .B(n54), .Z(DIFF[24]) );
  XOR2_X1 U5 ( .A(n90), .B(n40), .Z(DIFF[29]) );
  XOR2_X1 U6 ( .A(n86), .B(n55), .Z(DIFF[25]) );
  XOR2_X1 U7 ( .A(n87), .B(n37), .Z(DIFF[26]) );
  XOR2_X1 U8 ( .A(n88), .B(n38), .Z(DIFF[27]) );
  XOR2_X1 U9 ( .A(n89), .B(n39), .Z(DIFF[28]) );
  XOR2_X1 U10 ( .A(n73), .B(n44), .Z(DIFF[12]) );
  XOR2_X1 U11 ( .A(n74), .B(n28), .Z(DIFF[13]) );
  XOR2_X1 U12 ( .A(n75), .B(n29), .Z(DIFF[14]) );
  XOR2_X1 U13 ( .A(n76), .B(n45), .Z(DIFF[15]) );
  XOR2_X1 U14 ( .A(n77), .B(n46), .Z(DIFF[16]) );
  XOR2_X1 U15 ( .A(n78), .B(n47), .Z(DIFF[17]) );
  XOR2_X1 U16 ( .A(n79), .B(n48), .Z(DIFF[18]) );
  XOR2_X1 U17 ( .A(n80), .B(n49), .Z(DIFF[19]) );
  XOR2_X1 U18 ( .A(n81), .B(n50), .Z(DIFF[20]) );
  XOR2_X1 U19 ( .A(n82), .B(n51), .Z(DIFF[21]) );
  XOR2_X1 U20 ( .A(n83), .B(n52), .Z(DIFF[22]) );
  XOR2_X1 U21 ( .A(n70), .B(n36), .Z(DIFF[9]) );
  XOR2_X1 U22 ( .A(n71), .B(n42), .Z(DIFF[10]) );
  XOR2_X1 U23 ( .A(n72), .B(n43), .Z(DIFF[11]) );
  XOR2_X1 U24 ( .A(n69), .B(n35), .Z(DIFF[8]) );
  XOR2_X1 U25 ( .A(n66), .B(n32), .Z(DIFF[5]) );
  XOR2_X1 U26 ( .A(n67), .B(n33), .Z(DIFF[6]) );
  XOR2_X1 U27 ( .A(n68), .B(n34), .Z(DIFF[7]) );
  AND2_X1 U28 ( .A1(n73), .A2(n44), .ZN(n28) );
  AND2_X1 U29 ( .A1(n74), .A2(n28), .ZN(n29) );
  AND2_X1 U30 ( .A1(n63), .A2(n59), .ZN(n30) );
  AND2_X1 U31 ( .A1(n64), .A2(n30), .ZN(n31) );
  AND2_X1 U32 ( .A1(n65), .A2(n31), .ZN(n32) );
  AND2_X1 U33 ( .A1(n66), .A2(n32), .ZN(n33) );
  AND2_X1 U34 ( .A1(n67), .A2(n33), .ZN(n34) );
  AND2_X1 U35 ( .A1(n68), .A2(n34), .ZN(n35) );
  AND2_X1 U36 ( .A1(n69), .A2(n35), .ZN(n36) );
  AND2_X1 U37 ( .A1(n86), .A2(n55), .ZN(n37) );
  AND2_X1 U38 ( .A1(n87), .A2(n37), .ZN(n38) );
  AND2_X1 U39 ( .A1(n88), .A2(n38), .ZN(n39) );
  AND2_X1 U40 ( .A1(n89), .A2(n39), .ZN(n40) );
  AND2_X1 U41 ( .A1(n90), .A2(n40), .ZN(n41) );
  AND2_X1 U42 ( .A1(n70), .A2(n36), .ZN(n42) );
  AND2_X1 U43 ( .A1(n71), .A2(n42), .ZN(n43) );
  AND2_X1 U44 ( .A1(n72), .A2(n43), .ZN(n44) );
  AND2_X1 U45 ( .A1(n75), .A2(n29), .ZN(n45) );
  AND2_X1 U46 ( .A1(n76), .A2(n45), .ZN(n46) );
  AND2_X1 U47 ( .A1(n77), .A2(n46), .ZN(n47) );
  AND2_X1 U48 ( .A1(n78), .A2(n47), .ZN(n48) );
  AND2_X1 U49 ( .A1(n79), .A2(n48), .ZN(n49) );
  AND2_X1 U50 ( .A1(n80), .A2(n49), .ZN(n50) );
  AND2_X1 U51 ( .A1(n81), .A2(n50), .ZN(n51) );
  AND2_X1 U52 ( .A1(n82), .A2(n51), .ZN(n52) );
  AND2_X1 U53 ( .A1(n83), .A2(n52), .ZN(n53) );
  AND2_X1 U54 ( .A1(n84), .A2(n53), .ZN(n54) );
  AND2_X1 U55 ( .A1(n85), .A2(n54), .ZN(n55) );
  XOR2_X1 U56 ( .A(n63), .B(n59), .Z(DIFF[2]) );
  XOR2_X1 U57 ( .A(n64), .B(n30), .Z(DIFF[3]) );
  XOR2_X1 U58 ( .A(n65), .B(n31), .Z(DIFF[4]) );
  INV_X1 U59 ( .A(B[1]), .ZN(n92) );
  INV_X1 U60 ( .A(B[2]), .ZN(n63) );
  INV_X1 U61 ( .A(B[3]), .ZN(n64) );
  INV_X1 U62 ( .A(B[4]), .ZN(n65) );
  INV_X1 U63 ( .A(B[5]), .ZN(n66) );
  INV_X1 U64 ( .A(B[6]), .ZN(n67) );
  INV_X1 U65 ( .A(B[7]), .ZN(n68) );
  INV_X1 U66 ( .A(B[8]), .ZN(n69) );
  INV_X1 U67 ( .A(B[9]), .ZN(n70) );
  NAND2_X1 U68 ( .A1(n91), .A2(n41), .ZN(n61) );
  AND2_X1 U69 ( .A1(n92), .A2(n62), .ZN(n59) );
  INV_X1 U70 ( .A(B[10]), .ZN(n71) );
  INV_X1 U71 ( .A(B[11]), .ZN(n72) );
  INV_X1 U72 ( .A(B[12]), .ZN(n73) );
  INV_X1 U73 ( .A(B[13]), .ZN(n74) );
  INV_X1 U74 ( .A(B[14]), .ZN(n75) );
  INV_X1 U75 ( .A(B[15]), .ZN(n76) );
  INV_X1 U76 ( .A(B[16]), .ZN(n77) );
  INV_X1 U77 ( .A(B[17]), .ZN(n78) );
  INV_X1 U78 ( .A(B[18]), .ZN(n79) );
  INV_X1 U79 ( .A(B[19]), .ZN(n80) );
  INV_X1 U80 ( .A(B[25]), .ZN(n86) );
  INV_X1 U81 ( .A(B[26]), .ZN(n87) );
  INV_X1 U82 ( .A(B[27]), .ZN(n88) );
  INV_X1 U83 ( .A(B[28]), .ZN(n89) );
  INV_X1 U84 ( .A(B[29]), .ZN(n90) );
  INV_X1 U85 ( .A(B[20]), .ZN(n81) );
  INV_X1 U86 ( .A(B[21]), .ZN(n82) );
  INV_X1 U87 ( .A(B[22]), .ZN(n83) );
  INV_X1 U88 ( .A(B[23]), .ZN(n84) );
  INV_X1 U89 ( .A(B[24]), .ZN(n85) );
  INV_X1 U90 ( .A(B[30]), .ZN(n91) );
  XOR2_X1 U91 ( .A(n92), .B(n62), .Z(DIFF[1]) );
  INV_X1 U92 ( .A(\B[0] ), .ZN(n62) );
endmodule


module negate_NBIT32_7 ( A, Y );
  input [31:0] A;
  output [31:0] Y;


  negate_NBIT32_7_DW01_sub_0 sub_add_14_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .B(A), .CI(1'b0), .DIFF(Y) );
endmodule


module negate_NBIT32_6_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n59, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U1 ( .A(n65), .B(n8), .Z(DIFF[4]) );
  XOR2_X1 U2 ( .A(n66), .B(n9), .Z(DIFF[5]) );
  XOR2_X1 U3 ( .A(n64), .B(n7), .Z(DIFF[3]) );
  NAND2_X1 U4 ( .A1(n91), .A2(n18), .ZN(n61) );
  AND2_X1 U5 ( .A1(n73), .A2(n20), .ZN(n4) );
  AND2_X1 U6 ( .A1(n74), .A2(n4), .ZN(n5) );
  AND2_X1 U7 ( .A1(n75), .A2(n5), .ZN(n6) );
  AND2_X1 U8 ( .A1(n92), .A2(n59), .ZN(n7) );
  AND2_X1 U9 ( .A1(n64), .A2(n7), .ZN(n8) );
  AND2_X1 U10 ( .A1(n65), .A2(n8), .ZN(n9) );
  AND2_X1 U11 ( .A1(n66), .A2(n9), .ZN(n10) );
  AND2_X1 U12 ( .A1(n67), .A2(n10), .ZN(n11) );
  AND2_X1 U13 ( .A1(n68), .A2(n11), .ZN(n12) );
  AND2_X1 U14 ( .A1(n69), .A2(n12), .ZN(n13) );
  AND2_X1 U15 ( .A1(n70), .A2(n13), .ZN(n14) );
  AND2_X1 U16 ( .A1(n87), .A2(n31), .ZN(n15) );
  AND2_X1 U17 ( .A1(n88), .A2(n15), .ZN(n16) );
  AND2_X1 U18 ( .A1(n89), .A2(n16), .ZN(n17) );
  AND2_X1 U19 ( .A1(n90), .A2(n17), .ZN(n18) );
  AND2_X1 U20 ( .A1(n71), .A2(n14), .ZN(n19) );
  AND2_X1 U21 ( .A1(n72), .A2(n19), .ZN(n20) );
  AND2_X1 U22 ( .A1(n76), .A2(n6), .ZN(n21) );
  AND2_X1 U23 ( .A1(n77), .A2(n21), .ZN(n22) );
  AND2_X1 U24 ( .A1(n78), .A2(n22), .ZN(n23) );
  AND2_X1 U25 ( .A1(n79), .A2(n23), .ZN(n24) );
  AND2_X1 U26 ( .A1(n80), .A2(n24), .ZN(n25) );
  AND2_X1 U27 ( .A1(n81), .A2(n25), .ZN(n26) );
  AND2_X1 U28 ( .A1(n82), .A2(n26), .ZN(n27) );
  AND2_X1 U29 ( .A1(n83), .A2(n27), .ZN(n28) );
  AND2_X1 U30 ( .A1(n84), .A2(n28), .ZN(n29) );
  AND2_X1 U31 ( .A1(n85), .A2(n29), .ZN(n30) );
  AND2_X1 U32 ( .A1(n86), .A2(n30), .ZN(n31) );
  XOR2_X1 U33 ( .A(n87), .B(n31), .Z(DIFF[26]) );
  XOR2_X1 U34 ( .A(n88), .B(n15), .Z(DIFF[27]) );
  XOR2_X1 U35 ( .A(n89), .B(n16), .Z(DIFF[28]) );
  XOR2_X1 U36 ( .A(n90), .B(n17), .Z(DIFF[29]) );
  XOR2_X1 U37 ( .A(n91), .B(n18), .Z(DIFF[30]) );
  XOR2_X1 U38 ( .A(n85), .B(n29), .Z(DIFF[24]) );
  XOR2_X1 U39 ( .A(n86), .B(n30), .Z(DIFF[25]) );
  XOR2_X1 U40 ( .A(n74), .B(n4), .Z(DIFF[13]) );
  XOR2_X1 U41 ( .A(n75), .B(n5), .Z(DIFF[14]) );
  XOR2_X1 U42 ( .A(n76), .B(n6), .Z(DIFF[15]) );
  XOR2_X1 U43 ( .A(n77), .B(n21), .Z(DIFF[16]) );
  XOR2_X1 U44 ( .A(n78), .B(n22), .Z(DIFF[17]) );
  XOR2_X1 U45 ( .A(n79), .B(n23), .Z(DIFF[18]) );
  XOR2_X1 U46 ( .A(n80), .B(n24), .Z(DIFF[19]) );
  XOR2_X1 U47 ( .A(n81), .B(n25), .Z(DIFF[20]) );
  XOR2_X1 U48 ( .A(n82), .B(n26), .Z(DIFF[21]) );
  XOR2_X1 U49 ( .A(n83), .B(n27), .Z(DIFF[22]) );
  XOR2_X1 U50 ( .A(n84), .B(n28), .Z(DIFF[23]) );
  XOR2_X1 U51 ( .A(n67), .B(n10), .Z(DIFF[6]) );
  XOR2_X1 U52 ( .A(n68), .B(n11), .Z(DIFF[7]) );
  XOR2_X1 U53 ( .A(n69), .B(n12), .Z(DIFF[8]) );
  XOR2_X1 U54 ( .A(n70), .B(n13), .Z(DIFF[9]) );
  XOR2_X1 U55 ( .A(n71), .B(n14), .Z(DIFF[10]) );
  XOR2_X1 U56 ( .A(n72), .B(n19), .Z(DIFF[11]) );
  XOR2_X1 U57 ( .A(n73), .B(n20), .Z(DIFF[12]) );
  XOR2_X1 U58 ( .A(n92), .B(n59), .Z(DIFF[2]) );
  INV_X1 U59 ( .A(B[2]), .ZN(n92) );
  INV_X1 U60 ( .A(B[3]), .ZN(n64) );
  INV_X1 U61 ( .A(B[4]), .ZN(n65) );
  INV_X1 U62 ( .A(B[5]), .ZN(n66) );
  INV_X1 U63 ( .A(B[6]), .ZN(n67) );
  INV_X1 U64 ( .A(B[7]), .ZN(n68) );
  INV_X1 U65 ( .A(B[8]), .ZN(n69) );
  INV_X1 U66 ( .A(B[9]), .ZN(n70) );
  XOR2_X1 U67 ( .A(B[31]), .B(n61), .Z(DIFF[31]) );
  INV_X1 U68 ( .A(B[10]), .ZN(n71) );
  INV_X1 U69 ( .A(B[11]), .ZN(n72) );
  INV_X1 U70 ( .A(B[12]), .ZN(n73) );
  INV_X1 U71 ( .A(B[13]), .ZN(n74) );
  INV_X1 U72 ( .A(B[14]), .ZN(n75) );
  INV_X1 U73 ( .A(B[15]), .ZN(n76) );
  INV_X1 U74 ( .A(B[16]), .ZN(n77) );
  INV_X1 U75 ( .A(B[17]), .ZN(n78) );
  INV_X1 U76 ( .A(B[18]), .ZN(n79) );
  INV_X1 U77 ( .A(B[19]), .ZN(n80) );
  INV_X1 U78 ( .A(B[20]), .ZN(n81) );
  INV_X1 U79 ( .A(B[26]), .ZN(n87) );
  INV_X1 U80 ( .A(B[27]), .ZN(n88) );
  INV_X1 U81 ( .A(B[28]), .ZN(n89) );
  INV_X1 U82 ( .A(B[29]), .ZN(n90) );
  INV_X1 U83 ( .A(B[30]), .ZN(n91) );
  INV_X1 U84 ( .A(B[21]), .ZN(n82) );
  INV_X1 U85 ( .A(B[22]), .ZN(n83) );
  INV_X1 U86 ( .A(B[23]), .ZN(n84) );
  INV_X1 U87 ( .A(B[24]), .ZN(n85) );
  INV_X1 U88 ( .A(B[25]), .ZN(n86) );
  AND2_X1 U89 ( .A1(n63), .A2(n62), .ZN(n59) );
  XOR2_X1 U90 ( .A(n63), .B(n62), .Z(DIFF[1]) );
  INV_X1 U91 ( .A(\B[0] ), .ZN(n62) );
  INV_X1 U92 ( .A(B[1]), .ZN(n63) );
endmodule


module negate_NBIT32_6 ( A, Y );
  input [31:0] A;
  output [31:0] Y;


  negate_NBIT32_6_DW01_sub_0 sub_add_14_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .B(A), .CI(1'b0), .DIFF(Y) );
endmodule


module negate_NBIT32_5_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U1 ( .A(B[31]), .B(n61), .Z(DIFF[31]) );
  XOR2_X1 U2 ( .A(n86), .B(n53), .Z(DIFF[25]) );
  XOR2_X1 U3 ( .A(n87), .B(n54), .Z(DIFF[26]) );
  XOR2_X1 U4 ( .A(n91), .B(n43), .Z(DIFF[30]) );
  XOR2_X1 U5 ( .A(n88), .B(n55), .Z(DIFF[27]) );
  XOR2_X1 U6 ( .A(n89), .B(n41), .Z(DIFF[28]) );
  XOR2_X1 U7 ( .A(n90), .B(n42), .Z(DIFF[29]) );
  XOR2_X1 U8 ( .A(n85), .B(n52), .Z(DIFF[24]) );
  XOR2_X1 U9 ( .A(n74), .B(n29), .Z(DIFF[13]) );
  XOR2_X1 U10 ( .A(n75), .B(n30), .Z(DIFF[14]) );
  XOR2_X1 U11 ( .A(n76), .B(n31), .Z(DIFF[15]) );
  XOR2_X1 U12 ( .A(n77), .B(n32), .Z(DIFF[16]) );
  XOR2_X1 U13 ( .A(n78), .B(n45), .Z(DIFF[17]) );
  XOR2_X1 U14 ( .A(n79), .B(n46), .Z(DIFF[18]) );
  XOR2_X1 U15 ( .A(n80), .B(n47), .Z(DIFF[19]) );
  XOR2_X1 U16 ( .A(n81), .B(n48), .Z(DIFF[20]) );
  XOR2_X1 U17 ( .A(n82), .B(n49), .Z(DIFF[21]) );
  XOR2_X1 U18 ( .A(n83), .B(n50), .Z(DIFF[22]) );
  XOR2_X1 U19 ( .A(n84), .B(n51), .Z(DIFF[23]) );
  XOR2_X1 U20 ( .A(n72), .B(n40), .Z(DIFF[11]) );
  XOR2_X1 U21 ( .A(n73), .B(n44), .Z(DIFF[12]) );
  XOR2_X1 U22 ( .A(n71), .B(n39), .Z(DIFF[10]) );
  XOR2_X1 U23 ( .A(n67), .B(n35), .Z(DIFF[6]) );
  XOR2_X1 U24 ( .A(n68), .B(n36), .Z(DIFF[7]) );
  XOR2_X1 U25 ( .A(n69), .B(n37), .Z(DIFF[8]) );
  XOR2_X1 U26 ( .A(n70), .B(n38), .Z(DIFF[9]) );
  XOR2_X1 U27 ( .A(n64), .B(n60), .Z(DIFF[2]) );
  XOR2_X1 U28 ( .A(n63), .B(n62), .Z(DIFF[1]) );
  AND2_X1 U29 ( .A1(n73), .A2(n44), .ZN(n29) );
  AND2_X1 U30 ( .A1(n74), .A2(n29), .ZN(n30) );
  AND2_X1 U31 ( .A1(n75), .A2(n30), .ZN(n31) );
  AND2_X1 U32 ( .A1(n76), .A2(n31), .ZN(n32) );
  AND2_X1 U33 ( .A1(n92), .A2(n59), .ZN(n33) );
  AND2_X1 U34 ( .A1(n65), .A2(n33), .ZN(n34) );
  AND2_X1 U35 ( .A1(n66), .A2(n34), .ZN(n35) );
  AND2_X1 U36 ( .A1(n67), .A2(n35), .ZN(n36) );
  AND2_X1 U37 ( .A1(n68), .A2(n36), .ZN(n37) );
  AND2_X1 U38 ( .A1(n69), .A2(n37), .ZN(n38) );
  AND2_X1 U39 ( .A1(n70), .A2(n38), .ZN(n39) );
  AND2_X1 U40 ( .A1(n71), .A2(n39), .ZN(n40) );
  AND2_X1 U41 ( .A1(n88), .A2(n55), .ZN(n41) );
  AND2_X1 U42 ( .A1(n89), .A2(n41), .ZN(n42) );
  AND2_X1 U43 ( .A1(n90), .A2(n42), .ZN(n43) );
  AND2_X1 U44 ( .A1(n72), .A2(n40), .ZN(n44) );
  AND2_X1 U45 ( .A1(n77), .A2(n32), .ZN(n45) );
  AND2_X1 U46 ( .A1(n78), .A2(n45), .ZN(n46) );
  AND2_X1 U47 ( .A1(n79), .A2(n46), .ZN(n47) );
  AND2_X1 U48 ( .A1(n80), .A2(n47), .ZN(n48) );
  AND2_X1 U49 ( .A1(n81), .A2(n48), .ZN(n49) );
  AND2_X1 U50 ( .A1(n82), .A2(n49), .ZN(n50) );
  AND2_X1 U51 ( .A1(n83), .A2(n50), .ZN(n51) );
  AND2_X1 U52 ( .A1(n84), .A2(n51), .ZN(n52) );
  AND2_X1 U53 ( .A1(n85), .A2(n52), .ZN(n53) );
  AND2_X1 U54 ( .A1(n86), .A2(n53), .ZN(n54) );
  AND2_X1 U55 ( .A1(n87), .A2(n54), .ZN(n55) );
  XOR2_X1 U56 ( .A(n65), .B(n33), .Z(DIFF[4]) );
  XOR2_X1 U57 ( .A(n66), .B(n34), .Z(DIFF[5]) );
  XOR2_X1 U58 ( .A(n92), .B(n59), .Z(DIFF[3]) );
  INV_X1 U59 ( .A(B[3]), .ZN(n92) );
  INV_X1 U60 ( .A(B[4]), .ZN(n65) );
  INV_X1 U61 ( .A(B[5]), .ZN(n66) );
  INV_X1 U62 ( .A(B[6]), .ZN(n67) );
  INV_X1 U63 ( .A(B[7]), .ZN(n68) );
  INV_X1 U64 ( .A(B[8]), .ZN(n69) );
  INV_X1 U65 ( .A(B[9]), .ZN(n70) );
  NAND2_X1 U66 ( .A1(n91), .A2(n43), .ZN(n61) );
  INV_X1 U67 ( .A(B[10]), .ZN(n71) );
  INV_X1 U68 ( .A(B[11]), .ZN(n72) );
  INV_X1 U69 ( .A(B[12]), .ZN(n73) );
  INV_X1 U70 ( .A(B[13]), .ZN(n74) );
  INV_X1 U71 ( .A(B[14]), .ZN(n75) );
  INV_X1 U72 ( .A(B[15]), .ZN(n76) );
  INV_X1 U73 ( .A(B[16]), .ZN(n77) );
  INV_X1 U74 ( .A(B[17]), .ZN(n78) );
  INV_X1 U75 ( .A(B[18]), .ZN(n79) );
  INV_X1 U76 ( .A(B[19]), .ZN(n80) );
  INV_X1 U77 ( .A(B[27]), .ZN(n88) );
  INV_X1 U78 ( .A(B[28]), .ZN(n89) );
  INV_X1 U79 ( .A(B[29]), .ZN(n90) );
  INV_X1 U80 ( .A(B[30]), .ZN(n91) );
  INV_X1 U81 ( .A(B[20]), .ZN(n81) );
  INV_X1 U82 ( .A(B[21]), .ZN(n82) );
  INV_X1 U83 ( .A(B[22]), .ZN(n83) );
  INV_X1 U84 ( .A(B[23]), .ZN(n84) );
  INV_X1 U85 ( .A(B[24]), .ZN(n85) );
  INV_X1 U86 ( .A(B[25]), .ZN(n86) );
  INV_X1 U87 ( .A(B[26]), .ZN(n87) );
  AND2_X1 U88 ( .A1(n64), .A2(n60), .ZN(n59) );
  AND2_X1 U89 ( .A1(n63), .A2(n62), .ZN(n60) );
  INV_X1 U90 ( .A(\B[0] ), .ZN(n62) );
  INV_X1 U91 ( .A(B[1]), .ZN(n63) );
  INV_X1 U92 ( .A(B[2]), .ZN(n64) );
endmodule


module negate_NBIT32_5 ( A, Y );
  input [31:0] A;
  output [31:0] Y;


  negate_NBIT32_5_DW01_sub_0 sub_add_14_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .B(A), .CI(1'b0), .DIFF(Y) );
endmodule


module mux51_gen_NBIT32_0 ( A0, A1, A2, A3, A4, SEL, Y );
  input [31:0] A0;
  input [31:0] A1;
  input [31:0] A2;
  input [31:0] A3;
  input [31:0] A4;
  input [2:0] SEL;
  output [31:0] Y;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n1, n2,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86;

  BUF_X1 U2 ( .A(n8), .Z(n73) );
  BUF_X1 U3 ( .A(n8), .Z(n74) );
  BUF_X1 U4 ( .A(n9), .Z(n1) );
  BUF_X1 U5 ( .A(n5), .Z(n82) );
  BUF_X1 U6 ( .A(n5), .Z(n83) );
  BUF_X1 U7 ( .A(n5), .Z(n84) );
  BUF_X1 U8 ( .A(n6), .Z(n79) );
  BUF_X1 U9 ( .A(n6), .Z(n80) );
  BUF_X1 U10 ( .A(n7), .Z(n76) );
  BUF_X1 U11 ( .A(n7), .Z(n77) );
  BUF_X1 U12 ( .A(n8), .Z(n75) );
  BUF_X1 U13 ( .A(n6), .Z(n81) );
  BUF_X1 U14 ( .A(n7), .Z(n78) );
  INV_X1 U15 ( .A(SEL[1]), .ZN(n85) );
  BUF_X1 U16 ( .A(n9), .Z(n2) );
  BUF_X1 U17 ( .A(n9), .Z(n72) );
  NOR3_X1 U18 ( .A1(SEL[0]), .A2(SEL[2]), .A3(n85), .ZN(n5) );
  NOR3_X1 U19 ( .A1(SEL[0]), .A2(SEL[1]), .A3(n1), .ZN(n8) );
  NOR3_X1 U20 ( .A1(SEL[1]), .A2(SEL[2]), .A3(SEL[0]), .ZN(n9) );
  AND3_X1 U21 ( .A1(SEL[0]), .A2(n86), .A3(SEL[1]), .ZN(n7) );
  AND3_X1 U22 ( .A1(n85), .A2(n86), .A3(SEL[0]), .ZN(n6) );
  INV_X1 U23 ( .A(SEL[2]), .ZN(n86) );
  NAND2_X1 U24 ( .A1(n28), .A2(n29), .ZN(Y[29]) );
  AOI22_X1 U25 ( .A1(A4[29]), .A2(n74), .B1(A0[29]), .B2(n2), .ZN(n28) );
  AOI222_X1 U26 ( .A1(A2[29]), .A2(n83), .B1(A1[29]), .B2(n80), .C1(A3[29]), 
        .C2(n77), .ZN(n29) );
  NAND2_X1 U27 ( .A1(n24), .A2(n25), .ZN(Y[30]) );
  AOI22_X1 U28 ( .A1(A4[30]), .A2(n74), .B1(A0[30]), .B2(n72), .ZN(n24) );
  AOI222_X1 U29 ( .A1(A2[30]), .A2(n84), .B1(A1[30]), .B2(n80), .C1(A3[30]), 
        .C2(n77), .ZN(n25) );
  NAND2_X1 U30 ( .A1(n36), .A2(n37), .ZN(Y[25]) );
  AOI22_X1 U31 ( .A1(A4[25]), .A2(n74), .B1(A0[25]), .B2(n2), .ZN(n36) );
  AOI222_X1 U32 ( .A1(A2[25]), .A2(n83), .B1(A1[25]), .B2(n80), .C1(A3[25]), 
        .C2(n77), .ZN(n37) );
  NAND2_X1 U33 ( .A1(n34), .A2(n35), .ZN(Y[26]) );
  AOI22_X1 U34 ( .A1(A4[26]), .A2(n74), .B1(A0[26]), .B2(n2), .ZN(n34) );
  AOI222_X1 U35 ( .A1(A2[26]), .A2(n83), .B1(A1[26]), .B2(n80), .C1(A3[26]), 
        .C2(n77), .ZN(n35) );
  NAND2_X1 U36 ( .A1(n32), .A2(n33), .ZN(Y[27]) );
  AOI22_X1 U37 ( .A1(A4[27]), .A2(n74), .B1(A0[27]), .B2(n2), .ZN(n32) );
  AOI222_X1 U38 ( .A1(A2[27]), .A2(n83), .B1(A1[27]), .B2(n80), .C1(A3[27]), 
        .C2(n77), .ZN(n33) );
  NAND2_X1 U39 ( .A1(n30), .A2(n31), .ZN(Y[28]) );
  AOI22_X1 U40 ( .A1(A4[28]), .A2(n74), .B1(A0[28]), .B2(n2), .ZN(n30) );
  AOI222_X1 U41 ( .A1(A2[28]), .A2(n83), .B1(A1[28]), .B2(n80), .C1(A3[28]), 
        .C2(n77), .ZN(n31) );
  NAND2_X1 U42 ( .A1(n40), .A2(n41), .ZN(Y[23]) );
  AOI22_X1 U43 ( .A1(A4[23]), .A2(n74), .B1(A0[23]), .B2(n2), .ZN(n40) );
  AOI222_X1 U44 ( .A1(A2[23]), .A2(n83), .B1(A1[23]), .B2(n80), .C1(A3[23]), 
        .C2(n77), .ZN(n41) );
  NAND2_X1 U45 ( .A1(n38), .A2(n39), .ZN(Y[24]) );
  AOI22_X1 U46 ( .A1(A4[24]), .A2(n74), .B1(A0[24]), .B2(n2), .ZN(n38) );
  AOI222_X1 U47 ( .A1(A2[24]), .A2(n83), .B1(A1[24]), .B2(n80), .C1(A3[24]), 
        .C2(n77), .ZN(n39) );
  NAND2_X1 U48 ( .A1(n22), .A2(n23), .ZN(Y[31]) );
  AOI22_X1 U49 ( .A1(A4[31]), .A2(n75), .B1(A0[31]), .B2(n72), .ZN(n22) );
  AOI222_X1 U50 ( .A1(A2[31]), .A2(n84), .B1(A1[31]), .B2(n81), .C1(A3[31]), 
        .C2(n78), .ZN(n23) );
  NAND2_X1 U51 ( .A1(n64), .A2(n65), .ZN(Y[12]) );
  AOI22_X1 U52 ( .A1(A4[12]), .A2(n73), .B1(A0[12]), .B2(n1), .ZN(n64) );
  AOI222_X1 U53 ( .A1(A2[12]), .A2(n82), .B1(A1[12]), .B2(n79), .C1(A3[12]), 
        .C2(n76), .ZN(n65) );
  NAND2_X1 U54 ( .A1(n62), .A2(n63), .ZN(Y[13]) );
  AOI22_X1 U55 ( .A1(A4[13]), .A2(n73), .B1(A0[13]), .B2(n1), .ZN(n62) );
  AOI222_X1 U56 ( .A1(A2[13]), .A2(n82), .B1(A1[13]), .B2(n79), .C1(A3[13]), 
        .C2(n76), .ZN(n63) );
  NAND2_X1 U57 ( .A1(n60), .A2(n61), .ZN(Y[14]) );
  AOI22_X1 U58 ( .A1(A4[14]), .A2(n73), .B1(A0[14]), .B2(n1), .ZN(n60) );
  AOI222_X1 U59 ( .A1(A2[14]), .A2(n82), .B1(A1[14]), .B2(n79), .C1(A3[14]), 
        .C2(n76), .ZN(n61) );
  NAND2_X1 U60 ( .A1(n58), .A2(n59), .ZN(Y[15]) );
  AOI22_X1 U61 ( .A1(A4[15]), .A2(n73), .B1(A0[15]), .B2(n1), .ZN(n58) );
  AOI222_X1 U62 ( .A1(A2[15]), .A2(n82), .B1(A1[15]), .B2(n79), .C1(A3[15]), 
        .C2(n76), .ZN(n59) );
  NAND2_X1 U63 ( .A1(n56), .A2(n57), .ZN(Y[16]) );
  AOI22_X1 U64 ( .A1(A4[16]), .A2(n73), .B1(A0[16]), .B2(n1), .ZN(n56) );
  AOI222_X1 U65 ( .A1(A2[16]), .A2(n82), .B1(A1[16]), .B2(n79), .C1(A3[16]), 
        .C2(n76), .ZN(n57) );
  NAND2_X1 U66 ( .A1(n54), .A2(n55), .ZN(Y[17]) );
  AOI22_X1 U67 ( .A1(A4[17]), .A2(n73), .B1(A0[17]), .B2(n1), .ZN(n54) );
  AOI222_X1 U68 ( .A1(A2[17]), .A2(n82), .B1(A1[17]), .B2(n79), .C1(A3[17]), 
        .C2(n76), .ZN(n55) );
  NAND2_X1 U69 ( .A1(n52), .A2(n53), .ZN(Y[18]) );
  AOI22_X1 U70 ( .A1(A4[18]), .A2(n73), .B1(A0[18]), .B2(n1), .ZN(n52) );
  AOI222_X1 U71 ( .A1(A2[18]), .A2(n82), .B1(A1[18]), .B2(n79), .C1(A3[18]), 
        .C2(n76), .ZN(n53) );
  NAND2_X1 U72 ( .A1(n50), .A2(n51), .ZN(Y[19]) );
  AOI22_X1 U73 ( .A1(A4[19]), .A2(n73), .B1(A0[19]), .B2(n1), .ZN(n50) );
  AOI222_X1 U74 ( .A1(A2[19]), .A2(n82), .B1(A1[19]), .B2(n79), .C1(A3[19]), 
        .C2(n76), .ZN(n51) );
  NAND2_X1 U75 ( .A1(n46), .A2(n47), .ZN(Y[20]) );
  AOI22_X1 U76 ( .A1(A4[20]), .A2(n74), .B1(A0[20]), .B2(n2), .ZN(n46) );
  AOI222_X1 U77 ( .A1(A2[20]), .A2(n83), .B1(A1[20]), .B2(n80), .C1(A3[20]), 
        .C2(n77), .ZN(n47) );
  NAND2_X1 U78 ( .A1(n44), .A2(n45), .ZN(Y[21]) );
  AOI22_X1 U79 ( .A1(A4[21]), .A2(n74), .B1(A0[21]), .B2(n2), .ZN(n44) );
  AOI222_X1 U80 ( .A1(A2[21]), .A2(n83), .B1(A1[21]), .B2(n80), .C1(A3[21]), 
        .C2(n77), .ZN(n45) );
  NAND2_X1 U81 ( .A1(n42), .A2(n43), .ZN(Y[22]) );
  AOI22_X1 U82 ( .A1(A4[22]), .A2(n74), .B1(A0[22]), .B2(n2), .ZN(n42) );
  AOI222_X1 U83 ( .A1(A2[22]), .A2(n83), .B1(A1[22]), .B2(n80), .C1(A3[22]), 
        .C2(n77), .ZN(n43) );
  NAND2_X1 U84 ( .A1(n10), .A2(n11), .ZN(Y[8]) );
  AOI22_X1 U85 ( .A1(A4[8]), .A2(n75), .B1(A0[8]), .B2(n72), .ZN(n10) );
  AOI222_X1 U86 ( .A1(A2[8]), .A2(n84), .B1(A1[8]), .B2(n81), .C1(A3[8]), .C2(
        n78), .ZN(n11) );
  NAND2_X1 U87 ( .A1(n3), .A2(n4), .ZN(Y[9]) );
  AOI22_X1 U88 ( .A1(A4[9]), .A2(n75), .B1(A0[9]), .B2(n72), .ZN(n3) );
  AOI222_X1 U89 ( .A1(A2[9]), .A2(n84), .B1(A1[9]), .B2(n81), .C1(A3[9]), .C2(
        n78), .ZN(n4) );
  NAND2_X1 U90 ( .A1(n68), .A2(n69), .ZN(Y[10]) );
  AOI22_X1 U91 ( .A1(A4[10]), .A2(n73), .B1(A0[10]), .B2(n1), .ZN(n68) );
  AOI222_X1 U92 ( .A1(A2[10]), .A2(n82), .B1(A1[10]), .B2(n79), .C1(A3[10]), 
        .C2(n76), .ZN(n69) );
  NAND2_X1 U93 ( .A1(n66), .A2(n67), .ZN(Y[11]) );
  AOI22_X1 U94 ( .A1(A4[11]), .A2(n73), .B1(A0[11]), .B2(n1), .ZN(n66) );
  AOI222_X1 U95 ( .A1(A2[11]), .A2(n82), .B1(A1[11]), .B2(n79), .C1(A3[11]), 
        .C2(n76), .ZN(n67) );
  NAND2_X1 U96 ( .A1(n48), .A2(n49), .ZN(Y[1]) );
  AOI222_X1 U97 ( .A1(A2[1]), .A2(n83), .B1(A1[1]), .B2(n79), .C1(A3[1]), .C2(
        n76), .ZN(n49) );
  AOI22_X1 U98 ( .A1(A4[1]), .A2(n73), .B1(A0[1]), .B2(n2), .ZN(n48) );
  NAND2_X1 U99 ( .A1(n26), .A2(n27), .ZN(Y[2]) );
  AOI222_X1 U100 ( .A1(A2[2]), .A2(n84), .B1(A1[2]), .B2(n80), .C1(A3[2]), 
        .C2(n77), .ZN(n27) );
  AOI22_X1 U101 ( .A1(A4[2]), .A2(n74), .B1(A0[2]), .B2(n2), .ZN(n26) );
  NAND2_X1 U102 ( .A1(n20), .A2(n21), .ZN(Y[3]) );
  AOI222_X1 U103 ( .A1(A2[3]), .A2(n84), .B1(A1[3]), .B2(n81), .C1(A3[3]), 
        .C2(n78), .ZN(n21) );
  AOI22_X1 U104 ( .A1(A4[3]), .A2(n75), .B1(A0[3]), .B2(n72), .ZN(n20) );
  NAND2_X1 U105 ( .A1(n18), .A2(n19), .ZN(Y[4]) );
  AOI222_X1 U106 ( .A1(A2[4]), .A2(n84), .B1(A1[4]), .B2(n81), .C1(A3[4]), 
        .C2(n78), .ZN(n19) );
  AOI22_X1 U107 ( .A1(A4[4]), .A2(n75), .B1(A0[4]), .B2(n72), .ZN(n18) );
  NAND2_X1 U108 ( .A1(n16), .A2(n17), .ZN(Y[5]) );
  AOI22_X1 U109 ( .A1(A4[5]), .A2(n75), .B1(A0[5]), .B2(n72), .ZN(n16) );
  AOI222_X1 U110 ( .A1(A2[5]), .A2(n84), .B1(A1[5]), .B2(n81), .C1(A3[5]), 
        .C2(n78), .ZN(n17) );
  NAND2_X1 U111 ( .A1(n14), .A2(n15), .ZN(Y[6]) );
  AOI22_X1 U112 ( .A1(A4[6]), .A2(n75), .B1(A0[6]), .B2(n72), .ZN(n14) );
  AOI222_X1 U113 ( .A1(A2[6]), .A2(n84), .B1(A1[6]), .B2(n81), .C1(A3[6]), 
        .C2(n78), .ZN(n15) );
  NAND2_X1 U114 ( .A1(n12), .A2(n13), .ZN(Y[7]) );
  AOI22_X1 U115 ( .A1(A4[7]), .A2(n75), .B1(A0[7]), .B2(n72), .ZN(n12) );
  AOI222_X1 U116 ( .A1(A2[7]), .A2(n84), .B1(A1[7]), .B2(n81), .C1(A3[7]), 
        .C2(n78), .ZN(n13) );
  NAND2_X1 U117 ( .A1(n70), .A2(n71), .ZN(Y[0]) );
  AOI22_X1 U118 ( .A1(A4[0]), .A2(n73), .B1(A0[0]), .B2(n1), .ZN(n70) );
  AOI222_X1 U119 ( .A1(A2[0]), .A2(n82), .B1(A1[0]), .B2(n79), .C1(A3[0]), 
        .C2(n76), .ZN(n71) );
endmodule


module mux51_gen_NBIT32_3 ( A0, A1, A2, A3, A4, SEL, Y );
  input [31:0] A0;
  input [31:0] A1;
  input [31:0] A2;
  input [31:0] A3;
  input [31:0] A4;
  input [2:0] SEL;
  output [31:0] Y;
  wire   n1, n2, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155;

  BUF_X1 U2 ( .A(n150), .Z(n73) );
  BUF_X1 U3 ( .A(n150), .Z(n74) );
  BUF_X1 U4 ( .A(n149), .Z(n1) );
  BUF_X1 U5 ( .A(n153), .Z(n82) );
  BUF_X1 U6 ( .A(n153), .Z(n83) );
  BUF_X1 U7 ( .A(n153), .Z(n84) );
  BUF_X1 U8 ( .A(n152), .Z(n79) );
  BUF_X1 U9 ( .A(n152), .Z(n80) );
  BUF_X1 U10 ( .A(n151), .Z(n76) );
  BUF_X1 U11 ( .A(n151), .Z(n77) );
  BUF_X1 U12 ( .A(n150), .Z(n75) );
  BUF_X1 U13 ( .A(n152), .Z(n81) );
  BUF_X1 U14 ( .A(n151), .Z(n78) );
  INV_X1 U15 ( .A(SEL[2]), .ZN(n86) );
  INV_X1 U16 ( .A(SEL[1]), .ZN(n85) );
  BUF_X1 U17 ( .A(n149), .Z(n2) );
  BUF_X1 U18 ( .A(n149), .Z(n72) );
  NOR3_X1 U19 ( .A1(SEL[0]), .A2(SEL[2]), .A3(n85), .ZN(n153) );
  NOR3_X1 U20 ( .A1(SEL[0]), .A2(SEL[1]), .A3(n1), .ZN(n150) );
  NOR3_X1 U21 ( .A1(SEL[1]), .A2(SEL[2]), .A3(SEL[0]), .ZN(n149) );
  AND3_X1 U22 ( .A1(SEL[0]), .A2(n86), .A3(SEL[1]), .ZN(n151) );
  AND3_X1 U23 ( .A1(n85), .A2(n86), .A3(SEL[0]), .ZN(n152) );
  NAND2_X1 U24 ( .A1(n126), .A2(n125), .ZN(Y[27]) );
  AOI22_X1 U25 ( .A1(A4[27]), .A2(n74), .B1(A0[27]), .B2(n2), .ZN(n126) );
  AOI222_X1 U26 ( .A1(A2[27]), .A2(n83), .B1(A1[27]), .B2(n80), .C1(A3[27]), 
        .C2(n77), .ZN(n125) );
  NAND2_X1 U27 ( .A1(n128), .A2(n127), .ZN(Y[28]) );
  AOI22_X1 U28 ( .A1(A4[28]), .A2(n74), .B1(A0[28]), .B2(n2), .ZN(n128) );
  AOI222_X1 U29 ( .A1(A2[28]), .A2(n83), .B1(A1[28]), .B2(n80), .C1(A3[28]), 
        .C2(n77), .ZN(n127) );
  NAND2_X1 U30 ( .A1(n130), .A2(n129), .ZN(Y[29]) );
  AOI22_X1 U31 ( .A1(A4[29]), .A2(n74), .B1(A0[29]), .B2(n2), .ZN(n130) );
  AOI222_X1 U32 ( .A1(A2[29]), .A2(n83), .B1(A1[29]), .B2(n80), .C1(A3[29]), 
        .C2(n77), .ZN(n129) );
  NAND2_X1 U33 ( .A1(n134), .A2(n133), .ZN(Y[30]) );
  AOI22_X1 U34 ( .A1(A4[30]), .A2(n74), .B1(A0[30]), .B2(n72), .ZN(n134) );
  AOI222_X1 U35 ( .A1(A2[30]), .A2(n84), .B1(A1[30]), .B2(n80), .C1(A3[30]), 
        .C2(n77), .ZN(n133) );
  NAND2_X1 U36 ( .A1(n136), .A2(n135), .ZN(Y[31]) );
  AOI22_X1 U37 ( .A1(A4[31]), .A2(n75), .B1(A0[31]), .B2(n72), .ZN(n136) );
  AOI222_X1 U38 ( .A1(A2[31]), .A2(n84), .B1(A1[31]), .B2(n81), .C1(A3[31]), 
        .C2(n78), .ZN(n135) );
  NAND2_X1 U39 ( .A1(n120), .A2(n119), .ZN(Y[24]) );
  AOI22_X1 U40 ( .A1(A4[24]), .A2(n74), .B1(A0[24]), .B2(n2), .ZN(n120) );
  AOI222_X1 U41 ( .A1(A2[24]), .A2(n83), .B1(A1[24]), .B2(n80), .C1(A3[24]), 
        .C2(n77), .ZN(n119) );
  NAND2_X1 U42 ( .A1(n122), .A2(n121), .ZN(Y[25]) );
  AOI22_X1 U43 ( .A1(A4[25]), .A2(n74), .B1(A0[25]), .B2(n2), .ZN(n122) );
  AOI222_X1 U44 ( .A1(A2[25]), .A2(n83), .B1(A1[25]), .B2(n80), .C1(A3[25]), 
        .C2(n77), .ZN(n121) );
  NAND2_X1 U45 ( .A1(n124), .A2(n123), .ZN(Y[26]) );
  AOI22_X1 U46 ( .A1(A4[26]), .A2(n74), .B1(A0[26]), .B2(n2), .ZN(n124) );
  AOI222_X1 U47 ( .A1(A2[26]), .A2(n83), .B1(A1[26]), .B2(n80), .C1(A3[26]), 
        .C2(n77), .ZN(n123) );
  NAND2_X1 U48 ( .A1(n96), .A2(n95), .ZN(Y[13]) );
  AOI22_X1 U49 ( .A1(A4[13]), .A2(n73), .B1(A0[13]), .B2(n1), .ZN(n96) );
  AOI222_X1 U50 ( .A1(A2[13]), .A2(n82), .B1(A1[13]), .B2(n79), .C1(A3[13]), 
        .C2(n76), .ZN(n95) );
  NAND2_X1 U51 ( .A1(n98), .A2(n97), .ZN(Y[14]) );
  AOI22_X1 U52 ( .A1(A4[14]), .A2(n73), .B1(A0[14]), .B2(n1), .ZN(n98) );
  AOI222_X1 U53 ( .A1(A2[14]), .A2(n82), .B1(A1[14]), .B2(n79), .C1(A3[14]), 
        .C2(n76), .ZN(n97) );
  NAND2_X1 U54 ( .A1(n100), .A2(n99), .ZN(Y[15]) );
  AOI22_X1 U55 ( .A1(A4[15]), .A2(n73), .B1(A0[15]), .B2(n1), .ZN(n100) );
  AOI222_X1 U56 ( .A1(A2[15]), .A2(n82), .B1(A1[15]), .B2(n79), .C1(A3[15]), 
        .C2(n76), .ZN(n99) );
  NAND2_X1 U57 ( .A1(n102), .A2(n101), .ZN(Y[16]) );
  AOI22_X1 U58 ( .A1(A4[16]), .A2(n73), .B1(A0[16]), .B2(n1), .ZN(n102) );
  AOI222_X1 U59 ( .A1(A2[16]), .A2(n82), .B1(A1[16]), .B2(n79), .C1(A3[16]), 
        .C2(n76), .ZN(n101) );
  NAND2_X1 U60 ( .A1(n104), .A2(n103), .ZN(Y[17]) );
  AOI22_X1 U61 ( .A1(A4[17]), .A2(n73), .B1(A0[17]), .B2(n1), .ZN(n104) );
  AOI222_X1 U62 ( .A1(A2[17]), .A2(n82), .B1(A1[17]), .B2(n79), .C1(A3[17]), 
        .C2(n76), .ZN(n103) );
  NAND2_X1 U63 ( .A1(n106), .A2(n105), .ZN(Y[18]) );
  AOI22_X1 U64 ( .A1(A4[18]), .A2(n73), .B1(A0[18]), .B2(n1), .ZN(n106) );
  AOI222_X1 U65 ( .A1(A2[18]), .A2(n82), .B1(A1[18]), .B2(n79), .C1(A3[18]), 
        .C2(n76), .ZN(n105) );
  NAND2_X1 U66 ( .A1(n108), .A2(n107), .ZN(Y[19]) );
  AOI22_X1 U67 ( .A1(A4[19]), .A2(n73), .B1(A0[19]), .B2(n1), .ZN(n108) );
  AOI222_X1 U68 ( .A1(A2[19]), .A2(n82), .B1(A1[19]), .B2(n79), .C1(A3[19]), 
        .C2(n76), .ZN(n107) );
  NAND2_X1 U69 ( .A1(n112), .A2(n111), .ZN(Y[20]) );
  AOI22_X1 U70 ( .A1(A4[20]), .A2(n74), .B1(A0[20]), .B2(n2), .ZN(n112) );
  AOI222_X1 U71 ( .A1(A2[20]), .A2(n83), .B1(A1[20]), .B2(n80), .C1(A3[20]), 
        .C2(n77), .ZN(n111) );
  NAND2_X1 U72 ( .A1(n114), .A2(n113), .ZN(Y[21]) );
  AOI22_X1 U73 ( .A1(A4[21]), .A2(n74), .B1(A0[21]), .B2(n2), .ZN(n114) );
  AOI222_X1 U74 ( .A1(A2[21]), .A2(n83), .B1(A1[21]), .B2(n80), .C1(A3[21]), 
        .C2(n77), .ZN(n113) );
  NAND2_X1 U75 ( .A1(n116), .A2(n115), .ZN(Y[22]) );
  AOI22_X1 U76 ( .A1(A4[22]), .A2(n74), .B1(A0[22]), .B2(n2), .ZN(n116) );
  AOI222_X1 U77 ( .A1(A2[22]), .A2(n83), .B1(A1[22]), .B2(n80), .C1(A3[22]), 
        .C2(n77), .ZN(n115) );
  NAND2_X1 U78 ( .A1(n118), .A2(n117), .ZN(Y[23]) );
  AOI22_X1 U79 ( .A1(A4[23]), .A2(n74), .B1(A0[23]), .B2(n2), .ZN(n118) );
  AOI222_X1 U80 ( .A1(A2[23]), .A2(n83), .B1(A1[23]), .B2(n80), .C1(A3[23]), 
        .C2(n77), .ZN(n117) );
  NAND2_X1 U81 ( .A1(n90), .A2(n89), .ZN(Y[10]) );
  AOI22_X1 U82 ( .A1(A4[10]), .A2(n73), .B1(A0[10]), .B2(n1), .ZN(n90) );
  AOI222_X1 U83 ( .A1(A2[10]), .A2(n82), .B1(A1[10]), .B2(n79), .C1(A3[10]), 
        .C2(n76), .ZN(n89) );
  NAND2_X1 U84 ( .A1(n92), .A2(n91), .ZN(Y[11]) );
  AOI22_X1 U85 ( .A1(A4[11]), .A2(n73), .B1(A0[11]), .B2(n1), .ZN(n92) );
  AOI222_X1 U86 ( .A1(A2[11]), .A2(n82), .B1(A1[11]), .B2(n79), .C1(A3[11]), 
        .C2(n76), .ZN(n91) );
  NAND2_X1 U87 ( .A1(n94), .A2(n93), .ZN(Y[12]) );
  AOI22_X1 U88 ( .A1(A4[12]), .A2(n73), .B1(A0[12]), .B2(n1), .ZN(n94) );
  AOI222_X1 U89 ( .A1(A2[12]), .A2(n82), .B1(A1[12]), .B2(n79), .C1(A3[12]), 
        .C2(n76), .ZN(n93) );
  NAND2_X1 U90 ( .A1(n138), .A2(n137), .ZN(Y[3]) );
  AOI222_X1 U91 ( .A1(A2[3]), .A2(n84), .B1(A1[3]), .B2(n81), .C1(A3[3]), .C2(
        n78), .ZN(n137) );
  AOI22_X1 U92 ( .A1(A4[3]), .A2(n75), .B1(A0[3]), .B2(n72), .ZN(n138) );
  NAND2_X1 U93 ( .A1(n140), .A2(n139), .ZN(Y[4]) );
  AOI222_X1 U94 ( .A1(A2[4]), .A2(n84), .B1(A1[4]), .B2(n81), .C1(A3[4]), .C2(
        n78), .ZN(n139) );
  AOI22_X1 U95 ( .A1(A4[4]), .A2(n75), .B1(A0[4]), .B2(n72), .ZN(n140) );
  NAND2_X1 U96 ( .A1(n142), .A2(n141), .ZN(Y[5]) );
  AOI222_X1 U97 ( .A1(A2[5]), .A2(n84), .B1(A1[5]), .B2(n81), .C1(A3[5]), .C2(
        n78), .ZN(n141) );
  AOI22_X1 U98 ( .A1(A4[5]), .A2(n75), .B1(A0[5]), .B2(n72), .ZN(n142) );
  NAND2_X1 U99 ( .A1(n144), .A2(n143), .ZN(Y[6]) );
  AOI22_X1 U100 ( .A1(A4[6]), .A2(n75), .B1(A0[6]), .B2(n72), .ZN(n144) );
  AOI222_X1 U101 ( .A1(A2[6]), .A2(n84), .B1(A1[6]), .B2(n81), .C1(A3[6]), 
        .C2(n78), .ZN(n143) );
  NAND2_X1 U102 ( .A1(n146), .A2(n145), .ZN(Y[7]) );
  AOI22_X1 U103 ( .A1(A4[7]), .A2(n75), .B1(A0[7]), .B2(n72), .ZN(n146) );
  AOI222_X1 U104 ( .A1(A2[7]), .A2(n84), .B1(A1[7]), .B2(n81), .C1(A3[7]), 
        .C2(n78), .ZN(n145) );
  NAND2_X1 U105 ( .A1(n148), .A2(n147), .ZN(Y[8]) );
  AOI22_X1 U106 ( .A1(A4[8]), .A2(n75), .B1(A0[8]), .B2(n72), .ZN(n148) );
  AOI222_X1 U107 ( .A1(A2[8]), .A2(n84), .B1(A1[8]), .B2(n81), .C1(A3[8]), 
        .C2(n78), .ZN(n147) );
  NAND2_X1 U108 ( .A1(n155), .A2(n154), .ZN(Y[9]) );
  AOI22_X1 U109 ( .A1(A4[9]), .A2(n75), .B1(A0[9]), .B2(n72), .ZN(n155) );
  AOI222_X1 U110 ( .A1(A2[9]), .A2(n84), .B1(A1[9]), .B2(n81), .C1(A3[9]), 
        .C2(n78), .ZN(n154) );
  NAND2_X1 U111 ( .A1(n132), .A2(n131), .ZN(Y[2]) );
  AOI22_X1 U112 ( .A1(A4[2]), .A2(n74), .B1(A0[2]), .B2(n2), .ZN(n132) );
  AOI222_X1 U113 ( .A1(A2[2]), .A2(n84), .B1(A1[2]), .B2(n80), .C1(A3[2]), 
        .C2(n77), .ZN(n131) );
  NAND2_X1 U114 ( .A1(n110), .A2(n109), .ZN(Y[1]) );
  AOI22_X1 U115 ( .A1(A4[1]), .A2(n73), .B1(A0[1]), .B2(n2), .ZN(n110) );
  AOI222_X1 U116 ( .A1(A2[1]), .A2(n83), .B1(A1[1]), .B2(n79), .C1(A3[1]), 
        .C2(n76), .ZN(n109) );
  NAND2_X1 U117 ( .A1(n88), .A2(n87), .ZN(Y[0]) );
  AOI22_X1 U118 ( .A1(A4[0]), .A2(n73), .B1(A0[0]), .B2(n1), .ZN(n88) );
  AOI222_X1 U119 ( .A1(A2[0]), .A2(n82), .B1(A1[0]), .B2(n79), .C1(A3[0]), 
        .C2(n76), .ZN(n87) );
endmodule


module shl1_NBIT32_2 ( A, Y );
  input [31:0] A;
  output [31:0] Y;
  wire   \A[30] , \A[29] , \A[28] , \A[27] , \A[26] , \A[25] , \A[24] ,
         \A[23] , \A[22] , \A[21] , \A[20] , \A[19] , \A[18] , \A[17] ,
         \A[16] , \A[15] , \A[14] , \A[13] , \A[12] , \A[11] , \A[10] , \A[9] ,
         \A[8] , \A[7] , \A[6] , \A[5] , \A[4] , \A[3] , \A[2] , \A[1] ,
         \A[0] ;
  assign Y[0] = 1'b0;
  assign Y[31] = \A[30] ;
  assign \A[30]  = A[30];
  assign Y[30] = \A[29] ;
  assign \A[29]  = A[29];
  assign Y[29] = \A[28] ;
  assign \A[28]  = A[28];
  assign Y[28] = \A[27] ;
  assign \A[27]  = A[27];
  assign Y[27] = \A[26] ;
  assign \A[26]  = A[26];
  assign Y[26] = \A[25] ;
  assign \A[25]  = A[25];
  assign Y[25] = \A[24] ;
  assign \A[24]  = A[24];
  assign Y[24] = \A[23] ;
  assign \A[23]  = A[23];
  assign Y[23] = \A[22] ;
  assign \A[22]  = A[22];
  assign Y[22] = \A[21] ;
  assign \A[21]  = A[21];
  assign Y[21] = \A[20] ;
  assign \A[20]  = A[20];
  assign Y[20] = \A[19] ;
  assign \A[19]  = A[19];
  assign Y[19] = \A[18] ;
  assign \A[18]  = A[18];
  assign Y[18] = \A[17] ;
  assign \A[17]  = A[17];
  assign Y[17] = \A[16] ;
  assign \A[16]  = A[16];
  assign Y[16] = \A[15] ;
  assign \A[15]  = A[15];
  assign Y[15] = \A[14] ;
  assign \A[14]  = A[14];
  assign Y[14] = \A[13] ;
  assign \A[13]  = A[13];
  assign Y[13] = \A[12] ;
  assign \A[12]  = A[12];
  assign Y[12] = \A[11] ;
  assign \A[11]  = A[11];
  assign Y[11] = \A[10] ;
  assign \A[10]  = A[10];
  assign Y[10] = \A[9] ;
  assign \A[9]  = A[9];
  assign Y[9] = \A[8] ;
  assign \A[8]  = A[8];
  assign Y[8] = \A[7] ;
  assign \A[7]  = A[7];
  assign Y[7] = \A[6] ;
  assign \A[6]  = A[6];
  assign Y[6] = \A[5] ;
  assign \A[5]  = A[5];
  assign Y[5] = \A[4] ;
  assign \A[4]  = A[4];
  assign Y[4] = \A[3] ;
  assign \A[3]  = A[3];
  assign Y[3] = \A[2] ;
  assign \A[2]  = A[2];
  assign Y[2] = \A[1] ;
  assign \A[1]  = A[1];
  assign Y[1] = \A[0] ;
  assign \A[0]  = A[0];

endmodule


module shl2_NBIT32_2 ( A, Y );
  input [31:0] A;
  output [31:0] Y;
  wire   \A[29] , \A[28] , \A[27] , \A[26] , \A[25] , \A[24] , \A[23] ,
         \A[22] , \A[21] , \A[20] , \A[19] , \A[18] , \A[17] , \A[16] ,
         \A[15] , \A[14] , \A[13] , \A[12] , \A[11] , \A[10] , \A[9] , \A[8] ,
         \A[7] , \A[6] , \A[5] , \A[4] , \A[3] , \A[2] , \A[1] , \A[0] ;
  assign Y[0] = 1'b0;
  assign Y[1] = 1'b0;
  assign Y[31] = \A[29] ;
  assign \A[29]  = A[29];
  assign Y[30] = \A[28] ;
  assign \A[28]  = A[28];
  assign Y[29] = \A[27] ;
  assign \A[27]  = A[27];
  assign Y[28] = \A[26] ;
  assign \A[26]  = A[26];
  assign Y[27] = \A[25] ;
  assign \A[25]  = A[25];
  assign Y[26] = \A[24] ;
  assign \A[24]  = A[24];
  assign Y[25] = \A[23] ;
  assign \A[23]  = A[23];
  assign Y[24] = \A[22] ;
  assign \A[22]  = A[22];
  assign Y[23] = \A[21] ;
  assign \A[21]  = A[21];
  assign Y[22] = \A[20] ;
  assign \A[20]  = A[20];
  assign Y[21] = \A[19] ;
  assign \A[19]  = A[19];
  assign Y[20] = \A[18] ;
  assign \A[18]  = A[18];
  assign Y[19] = \A[17] ;
  assign \A[17]  = A[17];
  assign Y[18] = \A[16] ;
  assign \A[16]  = A[16];
  assign Y[17] = \A[15] ;
  assign \A[15]  = A[15];
  assign Y[16] = \A[14] ;
  assign \A[14]  = A[14];
  assign Y[15] = \A[13] ;
  assign \A[13]  = A[13];
  assign Y[14] = \A[12] ;
  assign \A[12]  = A[12];
  assign Y[13] = \A[11] ;
  assign \A[11]  = A[11];
  assign Y[12] = \A[10] ;
  assign \A[10]  = A[10];
  assign Y[11] = \A[9] ;
  assign \A[9]  = A[9];
  assign Y[10] = \A[8] ;
  assign \A[8]  = A[8];
  assign Y[9] = \A[7] ;
  assign \A[7]  = A[7];
  assign Y[8] = \A[6] ;
  assign \A[6]  = A[6];
  assign Y[7] = \A[5] ;
  assign \A[5]  = A[5];
  assign Y[6] = \A[4] ;
  assign \A[4]  = A[4];
  assign Y[5] = \A[3] ;
  assign \A[3]  = A[3];
  assign Y[4] = \A[2] ;
  assign \A[2]  = A[2];
  assign Y[3] = \A[1] ;
  assign \A[1]  = A[1];
  assign Y[2] = \A[0] ;
  assign \A[0]  = A[0];

endmodule


module negate_NBIT32_4_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n54, n55,
         n56, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U1 ( .A(n87), .B(n4), .Z(DIFF[6]) );
  XOR2_X1 U2 ( .A(n88), .B(n3), .Z(DIFF[5]) );
  AND2_X1 U3 ( .A1(n89), .A2(n54), .ZN(n3) );
  AND2_X1 U4 ( .A1(n88), .A2(n3), .ZN(n4) );
  AND2_X1 U5 ( .A1(n87), .A2(n4), .ZN(n5) );
  AND2_X1 U6 ( .A1(n85), .A2(n28), .ZN(n6) );
  AND2_X1 U7 ( .A1(n84), .A2(n6), .ZN(n7) );
  AND2_X1 U8 ( .A1(n83), .A2(n7), .ZN(n8) );
  AND2_X1 U9 ( .A1(n82), .A2(n8), .ZN(n9) );
  AND2_X1 U10 ( .A1(n81), .A2(n9), .ZN(n10) );
  AND2_X1 U11 ( .A1(n80), .A2(n10), .ZN(n11) );
  AND2_X1 U12 ( .A1(n79), .A2(n11), .ZN(n12) );
  AND2_X1 U13 ( .A1(n78), .A2(n12), .ZN(n13) );
  AND2_X1 U14 ( .A1(n77), .A2(n13), .ZN(n14) );
  AND2_X1 U15 ( .A1(n76), .A2(n14), .ZN(n15) );
  AND2_X1 U16 ( .A1(n75), .A2(n15), .ZN(n16) );
  AND2_X1 U17 ( .A1(n74), .A2(n16), .ZN(n17) );
  AND2_X1 U18 ( .A1(n73), .A2(n17), .ZN(n18) );
  AND2_X1 U19 ( .A1(n72), .A2(n18), .ZN(n19) );
  AND2_X1 U20 ( .A1(n71), .A2(n19), .ZN(n20) );
  AND2_X1 U21 ( .A1(n70), .A2(n20), .ZN(n21) );
  AND2_X1 U22 ( .A1(n69), .A2(n21), .ZN(n22) );
  AND2_X1 U23 ( .A1(n68), .A2(n22), .ZN(n23) );
  AND2_X1 U24 ( .A1(n67), .A2(n23), .ZN(n24) );
  AND2_X1 U25 ( .A1(n66), .A2(n24), .ZN(n25) );
  AND2_X1 U26 ( .A1(n65), .A2(n25), .ZN(n26) );
  AND2_X1 U27 ( .A1(n64), .A2(n26), .ZN(n27) );
  AND2_X1 U28 ( .A1(n86), .A2(n5), .ZN(n28) );
  NAND2_X1 U29 ( .A1(n63), .A2(n27), .ZN(n61) );
  XOR2_X1 U30 ( .A(n63), .B(n27), .Z(DIFF[30]) );
  XOR2_X1 U31 ( .A(n64), .B(n26), .Z(DIFF[29]) );
  XOR2_X1 U32 ( .A(n65), .B(n25), .Z(DIFF[28]) );
  XOR2_X1 U33 ( .A(n66), .B(n24), .Z(DIFF[27]) );
  XOR2_X1 U34 ( .A(n67), .B(n23), .Z(DIFF[26]) );
  XOR2_X1 U35 ( .A(n68), .B(n22), .Z(DIFF[25]) );
  XOR2_X1 U36 ( .A(n69), .B(n21), .Z(DIFF[24]) );
  XOR2_X1 U37 ( .A(n70), .B(n20), .Z(DIFF[23]) );
  XOR2_X1 U38 ( .A(n71), .B(n19), .Z(DIFF[22]) );
  XOR2_X1 U39 ( .A(n72), .B(n18), .Z(DIFF[21]) );
  XOR2_X1 U40 ( .A(n73), .B(n17), .Z(DIFF[20]) );
  XOR2_X1 U41 ( .A(n74), .B(n16), .Z(DIFF[19]) );
  XOR2_X1 U42 ( .A(n75), .B(n15), .Z(DIFF[18]) );
  XOR2_X1 U43 ( .A(n76), .B(n14), .Z(DIFF[17]) );
  XOR2_X1 U44 ( .A(n77), .B(n13), .Z(DIFF[16]) );
  XOR2_X1 U45 ( .A(n78), .B(n12), .Z(DIFF[15]) );
  XOR2_X1 U46 ( .A(n79), .B(n11), .Z(DIFF[14]) );
  XOR2_X1 U47 ( .A(n80), .B(n10), .Z(DIFF[13]) );
  XOR2_X1 U48 ( .A(n81), .B(n9), .Z(DIFF[12]) );
  XOR2_X1 U49 ( .A(n82), .B(n8), .Z(DIFF[11]) );
  XOR2_X1 U50 ( .A(n83), .B(n7), .Z(DIFF[10]) );
  XOR2_X1 U51 ( .A(n84), .B(n6), .Z(DIFF[9]) );
  XOR2_X1 U52 ( .A(n85), .B(n28), .Z(DIFF[8]) );
  XOR2_X1 U53 ( .A(n86), .B(n5), .Z(DIFF[7]) );
  XOR2_X1 U54 ( .A(n89), .B(n54), .Z(DIFF[4]) );
  AND2_X1 U55 ( .A1(n90), .A2(n55), .ZN(n54) );
  AND2_X1 U56 ( .A1(n91), .A2(n56), .ZN(n55) );
  AND2_X1 U57 ( .A1(n92), .A2(n62), .ZN(n56) );
  XOR2_X1 U58 ( .A(n90), .B(n55), .Z(DIFF[3]) );
  XOR2_X1 U59 ( .A(n91), .B(n56), .Z(DIFF[2]) );
  XOR2_X1 U60 ( .A(n92), .B(n62), .Z(DIFF[1]) );
  INV_X1 U61 ( .A(B[4]), .ZN(n89) );
  INV_X1 U62 ( .A(B[5]), .ZN(n88) );
  INV_X1 U63 ( .A(B[6]), .ZN(n87) );
  INV_X1 U64 ( .A(B[7]), .ZN(n86) );
  INV_X1 U65 ( .A(B[8]), .ZN(n85) );
  INV_X1 U66 ( .A(B[9]), .ZN(n84) );
  INV_X1 U67 ( .A(B[10]), .ZN(n83) );
  INV_X1 U68 ( .A(B[11]), .ZN(n82) );
  INV_X1 U69 ( .A(B[12]), .ZN(n81) );
  INV_X1 U70 ( .A(B[13]), .ZN(n80) );
  XOR2_X1 U71 ( .A(B[31]), .B(n61), .Z(DIFF[31]) );
  INV_X1 U72 ( .A(B[14]), .ZN(n79) );
  INV_X1 U73 ( .A(B[15]), .ZN(n78) );
  INV_X1 U74 ( .A(B[16]), .ZN(n77) );
  INV_X1 U75 ( .A(B[17]), .ZN(n76) );
  INV_X1 U76 ( .A(B[18]), .ZN(n75) );
  INV_X1 U77 ( .A(B[19]), .ZN(n74) );
  INV_X1 U78 ( .A(B[20]), .ZN(n73) );
  INV_X1 U79 ( .A(B[21]), .ZN(n72) );
  INV_X1 U80 ( .A(B[22]), .ZN(n71) );
  INV_X1 U81 ( .A(B[23]), .ZN(n70) );
  INV_X1 U82 ( .A(B[24]), .ZN(n69) );
  INV_X1 U83 ( .A(B[25]), .ZN(n68) );
  INV_X1 U84 ( .A(B[26]), .ZN(n67) );
  INV_X1 U85 ( .A(B[27]), .ZN(n66) );
  INV_X1 U86 ( .A(B[28]), .ZN(n65) );
  INV_X1 U87 ( .A(B[29]), .ZN(n64) );
  INV_X1 U88 ( .A(B[30]), .ZN(n63) );
  INV_X1 U89 ( .A(\B[0] ), .ZN(n62) );
  INV_X1 U90 ( .A(B[1]), .ZN(n92) );
  INV_X1 U91 ( .A(B[2]), .ZN(n91) );
  INV_X1 U92 ( .A(B[3]), .ZN(n90) );
endmodule


module negate_NBIT32_4 ( A, Y );
  input [31:0] A;
  output [31:0] Y;


  negate_NBIT32_4_DW01_sub_0 sub_add_14_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .B(A), .CI(1'b0), .DIFF(Y) );
endmodule


module negate_NBIT32_3_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U1 ( .A(B[31]), .B(n61), .Z(DIFF[31]) );
  XOR2_X1 U2 ( .A(n64), .B(n54), .Z(DIFF[30]) );
  XOR2_X1 U3 ( .A(n65), .B(n53), .Z(DIFF[29]) );
  XOR2_X1 U4 ( .A(n66), .B(n52), .Z(DIFF[28]) );
  XOR2_X1 U5 ( .A(n67), .B(n51), .Z(DIFF[27]) );
  XOR2_X1 U6 ( .A(n68), .B(n50), .Z(DIFF[26]) );
  XOR2_X1 U7 ( .A(n69), .B(n49), .Z(DIFF[25]) );
  XOR2_X1 U8 ( .A(n70), .B(n48), .Z(DIFF[24]) );
  XOR2_X1 U9 ( .A(n71), .B(n47), .Z(DIFF[23]) );
  XOR2_X1 U10 ( .A(n72), .B(n46), .Z(DIFF[22]) );
  XOR2_X1 U11 ( .A(n73), .B(n45), .Z(DIFF[21]) );
  XOR2_X1 U12 ( .A(n74), .B(n44), .Z(DIFF[20]) );
  XOR2_X1 U13 ( .A(n75), .B(n43), .Z(DIFF[19]) );
  XOR2_X1 U14 ( .A(n76), .B(n42), .Z(DIFF[18]) );
  XOR2_X1 U15 ( .A(n77), .B(n41), .Z(DIFF[17]) );
  XOR2_X1 U16 ( .A(n78), .B(n40), .Z(DIFF[16]) );
  XOR2_X1 U17 ( .A(n79), .B(n39), .Z(DIFF[15]) );
  XOR2_X1 U18 ( .A(n80), .B(n38), .Z(DIFF[14]) );
  XOR2_X1 U19 ( .A(n81), .B(n37), .Z(DIFF[13]) );
  XOR2_X1 U20 ( .A(n82), .B(n36), .Z(DIFF[12]) );
  XOR2_X1 U21 ( .A(n83), .B(n35), .Z(DIFF[11]) );
  XOR2_X1 U22 ( .A(n85), .B(n33), .Z(DIFF[9]) );
  XOR2_X1 U23 ( .A(n86), .B(n32), .Z(DIFF[8]) );
  XOR2_X1 U24 ( .A(n84), .B(n34), .Z(DIFF[10]) );
  XOR2_X1 U25 ( .A(n87), .B(n31), .Z(DIFF[7]) );
  XOR2_X1 U26 ( .A(n90), .B(n57), .Z(DIFF[4]) );
  XOR2_X1 U27 ( .A(n91), .B(n59), .Z(DIFF[3]) );
  XOR2_X1 U28 ( .A(n92), .B(n60), .Z(DIFF[2]) );
  XOR2_X1 U29 ( .A(n63), .B(n62), .Z(DIFF[1]) );
  AND2_X1 U30 ( .A1(n89), .A2(n58), .ZN(n30) );
  AND2_X1 U31 ( .A1(n88), .A2(n30), .ZN(n31) );
  AND2_X1 U32 ( .A1(n87), .A2(n31), .ZN(n32) );
  AND2_X1 U33 ( .A1(n86), .A2(n32), .ZN(n33) );
  AND2_X1 U34 ( .A1(n85), .A2(n33), .ZN(n34) );
  AND2_X1 U35 ( .A1(n84), .A2(n34), .ZN(n35) );
  AND2_X1 U36 ( .A1(n83), .A2(n35), .ZN(n36) );
  AND2_X1 U37 ( .A1(n82), .A2(n36), .ZN(n37) );
  AND2_X1 U38 ( .A1(n81), .A2(n37), .ZN(n38) );
  AND2_X1 U39 ( .A1(n80), .A2(n38), .ZN(n39) );
  AND2_X1 U40 ( .A1(n79), .A2(n39), .ZN(n40) );
  AND2_X1 U41 ( .A1(n78), .A2(n40), .ZN(n41) );
  AND2_X1 U42 ( .A1(n77), .A2(n41), .ZN(n42) );
  AND2_X1 U43 ( .A1(n76), .A2(n42), .ZN(n43) );
  AND2_X1 U44 ( .A1(n75), .A2(n43), .ZN(n44) );
  AND2_X1 U45 ( .A1(n74), .A2(n44), .ZN(n45) );
  AND2_X1 U46 ( .A1(n73), .A2(n45), .ZN(n46) );
  AND2_X1 U47 ( .A1(n72), .A2(n46), .ZN(n47) );
  AND2_X1 U48 ( .A1(n71), .A2(n47), .ZN(n48) );
  AND2_X1 U49 ( .A1(n70), .A2(n48), .ZN(n49) );
  AND2_X1 U50 ( .A1(n69), .A2(n49), .ZN(n50) );
  AND2_X1 U51 ( .A1(n68), .A2(n50), .ZN(n51) );
  AND2_X1 U52 ( .A1(n67), .A2(n51), .ZN(n52) );
  AND2_X1 U53 ( .A1(n66), .A2(n52), .ZN(n53) );
  AND2_X1 U54 ( .A1(n65), .A2(n53), .ZN(n54) );
  XOR2_X1 U55 ( .A(n88), .B(n30), .Z(DIFF[6]) );
  XOR2_X1 U56 ( .A(n89), .B(n58), .Z(DIFF[5]) );
  AND2_X1 U57 ( .A1(n91), .A2(n59), .ZN(n57) );
  AND2_X1 U58 ( .A1(n90), .A2(n57), .ZN(n58) );
  AND2_X1 U59 ( .A1(n92), .A2(n60), .ZN(n59) );
  AND2_X1 U60 ( .A1(n63), .A2(n62), .ZN(n60) );
  NAND2_X1 U61 ( .A1(n64), .A2(n54), .ZN(n61) );
  INV_X1 U62 ( .A(B[5]), .ZN(n89) );
  INV_X1 U63 ( .A(B[6]), .ZN(n88) );
  INV_X1 U64 ( .A(B[7]), .ZN(n87) );
  INV_X1 U65 ( .A(B[8]), .ZN(n86) );
  INV_X1 U66 ( .A(B[9]), .ZN(n85) );
  INV_X1 U67 ( .A(B[10]), .ZN(n84) );
  INV_X1 U68 ( .A(B[11]), .ZN(n83) );
  INV_X1 U69 ( .A(B[12]), .ZN(n82) );
  INV_X1 U70 ( .A(B[13]), .ZN(n81) );
  INV_X1 U71 ( .A(B[14]), .ZN(n80) );
  INV_X1 U72 ( .A(B[15]), .ZN(n79) );
  INV_X1 U73 ( .A(B[16]), .ZN(n78) );
  INV_X1 U74 ( .A(B[17]), .ZN(n77) );
  INV_X1 U75 ( .A(B[18]), .ZN(n76) );
  INV_X1 U76 ( .A(B[19]), .ZN(n75) );
  INV_X1 U77 ( .A(B[20]), .ZN(n74) );
  INV_X1 U78 ( .A(B[21]), .ZN(n73) );
  INV_X1 U79 ( .A(B[22]), .ZN(n72) );
  INV_X1 U80 ( .A(B[23]), .ZN(n71) );
  INV_X1 U81 ( .A(B[24]), .ZN(n70) );
  INV_X1 U82 ( .A(B[25]), .ZN(n69) );
  INV_X1 U83 ( .A(B[26]), .ZN(n68) );
  INV_X1 U84 ( .A(B[27]), .ZN(n67) );
  INV_X1 U85 ( .A(B[28]), .ZN(n66) );
  INV_X1 U86 ( .A(B[29]), .ZN(n65) );
  INV_X1 U87 ( .A(B[30]), .ZN(n64) );
  INV_X1 U88 ( .A(\B[0] ), .ZN(n62) );
  INV_X1 U89 ( .A(B[1]), .ZN(n63) );
  INV_X1 U90 ( .A(B[2]), .ZN(n92) );
  INV_X1 U91 ( .A(B[3]), .ZN(n91) );
  INV_X1 U92 ( .A(B[4]), .ZN(n90) );
endmodule


module negate_NBIT32_3 ( A, Y );
  input [31:0] A;
  output [31:0] Y;


  negate_NBIT32_3_DW01_sub_0 sub_add_14_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .B(A), .CI(1'b0), .DIFF(Y) );
endmodule


module mux51_gen_NBIT32_2 ( A0, A1, A2, A3, A4, SEL, Y );
  input [31:0] A0;
  input [31:0] A1;
  input [31:0] A2;
  input [31:0] A3;
  input [31:0] A4;
  input [2:0] SEL;
  output [31:0] Y;
  wire   n1, n2, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155;

  BUF_X1 U2 ( .A(n150), .Z(n74) );
  BUF_X1 U3 ( .A(n150), .Z(n73) );
  BUF_X1 U4 ( .A(n149), .Z(n1) );
  BUF_X1 U5 ( .A(n153), .Z(n83) );
  BUF_X1 U6 ( .A(n153), .Z(n82) );
  BUF_X1 U7 ( .A(n153), .Z(n84) );
  BUF_X1 U8 ( .A(n152), .Z(n80) );
  BUF_X1 U9 ( .A(n152), .Z(n79) );
  BUF_X1 U10 ( .A(n151), .Z(n77) );
  BUF_X1 U11 ( .A(n151), .Z(n76) );
  BUF_X1 U12 ( .A(n150), .Z(n75) );
  BUF_X1 U13 ( .A(n152), .Z(n81) );
  BUF_X1 U14 ( .A(n151), .Z(n78) );
  BUF_X1 U15 ( .A(n149), .Z(n2) );
  BUF_X1 U16 ( .A(n149), .Z(n72) );
  NAND2_X1 U17 ( .A1(n134), .A2(n133), .ZN(Y[30]) );
  AOI22_X1 U18 ( .A1(A4[30]), .A2(n74), .B1(A0[30]), .B2(n72), .ZN(n134) );
  AOI222_X1 U19 ( .A1(A2[30]), .A2(n84), .B1(A1[30]), .B2(n80), .C1(A3[30]), 
        .C2(n77), .ZN(n133) );
  NAND2_X1 U20 ( .A1(n130), .A2(n129), .ZN(Y[29]) );
  AOI22_X1 U21 ( .A1(A4[29]), .A2(n74), .B1(A0[29]), .B2(n2), .ZN(n130) );
  AOI222_X1 U22 ( .A1(A2[29]), .A2(n83), .B1(A1[29]), .B2(n80), .C1(A3[29]), 
        .C2(n77), .ZN(n129) );
  NAND2_X1 U23 ( .A1(n128), .A2(n127), .ZN(Y[28]) );
  AOI22_X1 U24 ( .A1(A4[28]), .A2(n74), .B1(A0[28]), .B2(n2), .ZN(n128) );
  AOI222_X1 U25 ( .A1(A2[28]), .A2(n83), .B1(A1[28]), .B2(n80), .C1(A3[28]), 
        .C2(n77), .ZN(n127) );
  NAND2_X1 U26 ( .A1(n126), .A2(n125), .ZN(Y[27]) );
  AOI22_X1 U27 ( .A1(A4[27]), .A2(n74), .B1(A0[27]), .B2(n2), .ZN(n126) );
  AOI222_X1 U28 ( .A1(A2[27]), .A2(n83), .B1(A1[27]), .B2(n80), .C1(A3[27]), 
        .C2(n77), .ZN(n125) );
  NAND2_X1 U29 ( .A1(n124), .A2(n123), .ZN(Y[26]) );
  AOI22_X1 U30 ( .A1(A4[26]), .A2(n74), .B1(A0[26]), .B2(n2), .ZN(n124) );
  AOI222_X1 U31 ( .A1(A2[26]), .A2(n83), .B1(A1[26]), .B2(n80), .C1(A3[26]), 
        .C2(n77), .ZN(n123) );
  NAND2_X1 U32 ( .A1(n122), .A2(n121), .ZN(Y[25]) );
  AOI22_X1 U33 ( .A1(A4[25]), .A2(n74), .B1(A0[25]), .B2(n2), .ZN(n122) );
  AOI222_X1 U34 ( .A1(A2[25]), .A2(n83), .B1(A1[25]), .B2(n80), .C1(A3[25]), 
        .C2(n77), .ZN(n121) );
  NAND2_X1 U35 ( .A1(n120), .A2(n119), .ZN(Y[24]) );
  AOI22_X1 U36 ( .A1(A4[24]), .A2(n74), .B1(A0[24]), .B2(n2), .ZN(n120) );
  AOI222_X1 U37 ( .A1(A2[24]), .A2(n83), .B1(A1[24]), .B2(n80), .C1(A3[24]), 
        .C2(n77), .ZN(n119) );
  NAND2_X1 U38 ( .A1(n118), .A2(n117), .ZN(Y[23]) );
  AOI22_X1 U39 ( .A1(A4[23]), .A2(n74), .B1(A0[23]), .B2(n2), .ZN(n118) );
  AOI222_X1 U40 ( .A1(A2[23]), .A2(n83), .B1(A1[23]), .B2(n80), .C1(A3[23]), 
        .C2(n77), .ZN(n117) );
  NAND2_X1 U41 ( .A1(n116), .A2(n115), .ZN(Y[22]) );
  AOI22_X1 U42 ( .A1(A4[22]), .A2(n74), .B1(A0[22]), .B2(n2), .ZN(n116) );
  AOI222_X1 U43 ( .A1(A2[22]), .A2(n83), .B1(A1[22]), .B2(n80), .C1(A3[22]), 
        .C2(n77), .ZN(n115) );
  NAND2_X1 U44 ( .A1(n136), .A2(n135), .ZN(Y[31]) );
  AOI22_X1 U45 ( .A1(A4[31]), .A2(n75), .B1(A0[31]), .B2(n72), .ZN(n136) );
  AOI222_X1 U46 ( .A1(A2[31]), .A2(n84), .B1(A1[31]), .B2(n81), .C1(A3[31]), 
        .C2(n78), .ZN(n135) );
  NAND2_X1 U47 ( .A1(n114), .A2(n113), .ZN(Y[21]) );
  AOI22_X1 U48 ( .A1(A4[21]), .A2(n74), .B1(A0[21]), .B2(n2), .ZN(n114) );
  AOI222_X1 U49 ( .A1(A2[21]), .A2(n83), .B1(A1[21]), .B2(n80), .C1(A3[21]), 
        .C2(n77), .ZN(n113) );
  NAND2_X1 U50 ( .A1(n112), .A2(n111), .ZN(Y[20]) );
  AOI22_X1 U51 ( .A1(A4[20]), .A2(n74), .B1(A0[20]), .B2(n2), .ZN(n112) );
  AOI222_X1 U52 ( .A1(A2[20]), .A2(n83), .B1(A1[20]), .B2(n80), .C1(A3[20]), 
        .C2(n77), .ZN(n111) );
  NAND2_X1 U53 ( .A1(n108), .A2(n107), .ZN(Y[19]) );
  AOI22_X1 U54 ( .A1(A4[19]), .A2(n73), .B1(A0[19]), .B2(n1), .ZN(n108) );
  AOI222_X1 U55 ( .A1(A2[19]), .A2(n82), .B1(A1[19]), .B2(n79), .C1(A3[19]), 
        .C2(n76), .ZN(n107) );
  NAND2_X1 U56 ( .A1(n106), .A2(n105), .ZN(Y[18]) );
  AOI22_X1 U57 ( .A1(A4[18]), .A2(n73), .B1(A0[18]), .B2(n1), .ZN(n106) );
  AOI222_X1 U58 ( .A1(A2[18]), .A2(n82), .B1(A1[18]), .B2(n79), .C1(A3[18]), 
        .C2(n76), .ZN(n105) );
  NAND2_X1 U59 ( .A1(n104), .A2(n103), .ZN(Y[17]) );
  AOI22_X1 U60 ( .A1(A4[17]), .A2(n73), .B1(A0[17]), .B2(n1), .ZN(n104) );
  AOI222_X1 U61 ( .A1(A2[17]), .A2(n82), .B1(A1[17]), .B2(n79), .C1(A3[17]), 
        .C2(n76), .ZN(n103) );
  NAND2_X1 U62 ( .A1(n102), .A2(n101), .ZN(Y[16]) );
  AOI22_X1 U63 ( .A1(A4[16]), .A2(n73), .B1(A0[16]), .B2(n1), .ZN(n102) );
  AOI222_X1 U64 ( .A1(A2[16]), .A2(n82), .B1(A1[16]), .B2(n79), .C1(A3[16]), 
        .C2(n76), .ZN(n101) );
  NAND2_X1 U65 ( .A1(n100), .A2(n99), .ZN(Y[15]) );
  AOI22_X1 U66 ( .A1(A4[15]), .A2(n73), .B1(A0[15]), .B2(n1), .ZN(n100) );
  AOI222_X1 U67 ( .A1(A2[15]), .A2(n82), .B1(A1[15]), .B2(n79), .C1(A3[15]), 
        .C2(n76), .ZN(n99) );
  NAND2_X1 U68 ( .A1(n98), .A2(n97), .ZN(Y[14]) );
  AOI22_X1 U69 ( .A1(A4[14]), .A2(n73), .B1(A0[14]), .B2(n1), .ZN(n98) );
  AOI222_X1 U70 ( .A1(A2[14]), .A2(n82), .B1(A1[14]), .B2(n79), .C1(A3[14]), 
        .C2(n76), .ZN(n97) );
  NAND2_X1 U71 ( .A1(n96), .A2(n95), .ZN(Y[13]) );
  AOI22_X1 U72 ( .A1(A4[13]), .A2(n73), .B1(A0[13]), .B2(n1), .ZN(n96) );
  AOI222_X1 U73 ( .A1(A2[13]), .A2(n82), .B1(A1[13]), .B2(n79), .C1(A3[13]), 
        .C2(n76), .ZN(n95) );
  NAND2_X1 U74 ( .A1(n94), .A2(n93), .ZN(Y[12]) );
  AOI22_X1 U75 ( .A1(A4[12]), .A2(n73), .B1(A0[12]), .B2(n1), .ZN(n94) );
  AOI222_X1 U76 ( .A1(A2[12]), .A2(n82), .B1(A1[12]), .B2(n79), .C1(A3[12]), 
        .C2(n76), .ZN(n93) );
  NAND2_X1 U77 ( .A1(n92), .A2(n91), .ZN(Y[11]) );
  AOI22_X1 U78 ( .A1(A4[11]), .A2(n73), .B1(A0[11]), .B2(n1), .ZN(n92) );
  AOI222_X1 U79 ( .A1(A2[11]), .A2(n82), .B1(A1[11]), .B2(n79), .C1(A3[11]), 
        .C2(n76), .ZN(n91) );
  NAND2_X1 U80 ( .A1(n155), .A2(n154), .ZN(Y[9]) );
  AOI22_X1 U81 ( .A1(A4[9]), .A2(n75), .B1(A0[9]), .B2(n72), .ZN(n155) );
  AOI222_X1 U82 ( .A1(A2[9]), .A2(n84), .B1(A1[9]), .B2(n81), .C1(A3[9]), .C2(
        n78), .ZN(n154) );
  NAND2_X1 U83 ( .A1(n148), .A2(n147), .ZN(Y[8]) );
  AOI22_X1 U84 ( .A1(A4[8]), .A2(n75), .B1(A0[8]), .B2(n72), .ZN(n148) );
  AOI222_X1 U85 ( .A1(A2[8]), .A2(n84), .B1(A1[8]), .B2(n81), .C1(A3[8]), .C2(
        n78), .ZN(n147) );
  NAND2_X1 U86 ( .A1(n90), .A2(n89), .ZN(Y[10]) );
  AOI22_X1 U87 ( .A1(A4[10]), .A2(n73), .B1(A0[10]), .B2(n1), .ZN(n90) );
  AOI222_X1 U88 ( .A1(A2[10]), .A2(n82), .B1(A1[10]), .B2(n79), .C1(A3[10]), 
        .C2(n76), .ZN(n89) );
  NAND2_X1 U89 ( .A1(n140), .A2(n139), .ZN(Y[4]) );
  AOI22_X1 U90 ( .A1(A4[4]), .A2(n75), .B1(A0[4]), .B2(n72), .ZN(n140) );
  AOI222_X1 U91 ( .A1(A2[4]), .A2(n84), .B1(A1[4]), .B2(n81), .C1(A3[4]), .C2(
        n78), .ZN(n139) );
  NOR3_X1 U92 ( .A1(SEL[0]), .A2(SEL[1]), .A3(n1), .ZN(n150) );
  NOR3_X1 U93 ( .A1(SEL[1]), .A2(SEL[2]), .A3(SEL[0]), .ZN(n149) );
  NOR3_X1 U94 ( .A1(SEL[0]), .A2(SEL[2]), .A3(n86), .ZN(n153) );
  NAND2_X1 U95 ( .A1(n144), .A2(n143), .ZN(Y[6]) );
  AOI222_X1 U96 ( .A1(A2[6]), .A2(n84), .B1(A1[6]), .B2(n81), .C1(A3[6]), .C2(
        n78), .ZN(n143) );
  AOI22_X1 U97 ( .A1(A4[6]), .A2(n75), .B1(A0[6]), .B2(n72), .ZN(n144) );
  NAND2_X1 U98 ( .A1(n142), .A2(n141), .ZN(Y[5]) );
  AOI222_X1 U99 ( .A1(A2[5]), .A2(n84), .B1(A1[5]), .B2(n81), .C1(A3[5]), .C2(
        n78), .ZN(n141) );
  AOI22_X1 U100 ( .A1(A4[5]), .A2(n75), .B1(A0[5]), .B2(n72), .ZN(n142) );
  AND3_X1 U101 ( .A1(SEL[0]), .A2(n85), .A3(SEL[1]), .ZN(n151) );
  AND3_X1 U102 ( .A1(n86), .A2(n85), .A3(SEL[0]), .ZN(n152) );
  INV_X1 U103 ( .A(SEL[1]), .ZN(n86) );
  NAND2_X1 U104 ( .A1(n146), .A2(n145), .ZN(Y[7]) );
  AOI22_X1 U105 ( .A1(A4[7]), .A2(n75), .B1(A0[7]), .B2(n72), .ZN(n146) );
  AOI222_X1 U106 ( .A1(A2[7]), .A2(n84), .B1(A1[7]), .B2(n81), .C1(A3[7]), 
        .C2(n78), .ZN(n145) );
  INV_X1 U107 ( .A(SEL[2]), .ZN(n85) );
  NAND2_X1 U108 ( .A1(n110), .A2(n109), .ZN(Y[1]) );
  AOI22_X1 U109 ( .A1(A4[1]), .A2(n73), .B1(A0[1]), .B2(n2), .ZN(n110) );
  AOI222_X1 U110 ( .A1(A2[1]), .A2(n83), .B1(A1[1]), .B2(n79), .C1(A3[1]), 
        .C2(n76), .ZN(n109) );
  NAND2_X1 U111 ( .A1(n138), .A2(n137), .ZN(Y[3]) );
  AOI22_X1 U112 ( .A1(A4[3]), .A2(n75), .B1(A0[3]), .B2(n72), .ZN(n138) );
  AOI222_X1 U113 ( .A1(A2[3]), .A2(n84), .B1(A1[3]), .B2(n81), .C1(A3[3]), 
        .C2(n78), .ZN(n137) );
  NAND2_X1 U114 ( .A1(n132), .A2(n131), .ZN(Y[2]) );
  AOI22_X1 U115 ( .A1(A4[2]), .A2(n74), .B1(A0[2]), .B2(n2), .ZN(n132) );
  AOI222_X1 U116 ( .A1(A2[2]), .A2(n84), .B1(A1[2]), .B2(n80), .C1(A3[2]), 
        .C2(n77), .ZN(n131) );
  NAND2_X1 U117 ( .A1(n88), .A2(n87), .ZN(Y[0]) );
  AOI22_X1 U118 ( .A1(A4[0]), .A2(n73), .B1(A0[0]), .B2(n1), .ZN(n88) );
  AOI222_X1 U119 ( .A1(A2[0]), .A2(n82), .B1(A1[0]), .B2(n79), .C1(A3[0]), 
        .C2(n76), .ZN(n87) );
endmodule


module my_xor_192 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_191 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_190 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_189 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_188 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_187 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_186 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_185 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_184 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_183 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_182 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_181 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_180 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_179 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_178 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_177 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_176 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_175 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_174 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_173 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_172 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_171 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_170 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_169 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_168 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_167 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_166 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_165 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_164 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_163 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_162 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_161 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_160 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_159 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_158 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_157 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_156 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_155 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_154 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_153 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_152 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_151 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_150 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_149 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_148 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_147 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_146 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_145 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_144 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_143 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_142 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_141 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_140 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_139 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_138 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_137 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_136 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_135 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_134 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_133 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_132 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_131 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_130 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_129 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module pg_net_189 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_188 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_187 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_186 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_185 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_184 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_183 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_182 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_181 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_180 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_179 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_178 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_177 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_176 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_175 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_174 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_173 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_172 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_171 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_170 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_169 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_168 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_167 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_166 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_165 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_164 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_163 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_162 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_161 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_160 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_159 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_158 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_157 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_156 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_155 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_154 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_153 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_152 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_151 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_150 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_149 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_148 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_147 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_146 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_145 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_144 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_143 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_142 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_141 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_140 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_139 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_138 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_137 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_136 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_135 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_134 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_133 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_132 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_131 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_130 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_129 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_128 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_127 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_BLOCK_189 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_188 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_187 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_186 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_185 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_184 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_183 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_182 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_181 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_180 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_179 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_178 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_177 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_176 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_175 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_174 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_173 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_172 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_171 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_170 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_169 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_168 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_167 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_166 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_165 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_164 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_163 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_162 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_161 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_160 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_159 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_51 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_158 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_157 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_156 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_155 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_154 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_153 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_152 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_151 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_150 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AOI21_X1 U1 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_149 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_148 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_147 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_146 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_145 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_144 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_50 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_143 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_142 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_141 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_140 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_139 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_138 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_137 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_49 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_136 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_135 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_134 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_133 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_132 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_131 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_48 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_47 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_130 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AND2_X1 U2 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_129 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_128 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_127 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_46 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_45 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_44 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_43 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_42 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_41 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_40 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_39 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_38 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_37 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_36 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_35 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module CARRY_GENERATOR_NBIT64_NBIT_PER_BLOCK4_0 ( A, B, Cin, Co );
  input [63:0] A;
  input [63:0] B;
  output [15:0] Co;
  input Cin;
  wire   \g_vector[5][63] , \g_vector[5][59] , \g_vector[5][55] ,
         \g_vector[5][51] , \g_vector[4][63] , \g_vector[4][59] ,
         \g_vector[4][47] , \g_vector[4][43] , \g_vector[4][31] ,
         \g_vector[4][27] , \g_vector[3][63] , \g_vector[3][55] ,
         \g_vector[3][47] , \g_vector[3][39] , \g_vector[3][31] ,
         \g_vector[3][23] , \g_vector[3][15] , \g_vector[2][63] ,
         \g_vector[2][59] , \g_vector[2][55] , \g_vector[2][51] ,
         \g_vector[2][47] , \g_vector[2][43] , \g_vector[2][39] ,
         \g_vector[2][35] , \g_vector[2][31] , \g_vector[2][27] ,
         \g_vector[2][23] , \g_vector[2][19] , \g_vector[2][15] ,
         \g_vector[2][11] , \g_vector[2][7] , \g_vector[1][63] ,
         \g_vector[1][61] , \g_vector[1][59] , \g_vector[1][57] ,
         \g_vector[1][55] , \g_vector[1][53] , \g_vector[1][51] ,
         \g_vector[1][49] , \g_vector[1][47] , \g_vector[1][45] ,
         \g_vector[1][43] , \g_vector[1][41] , \g_vector[1][39] ,
         \g_vector[1][37] , \g_vector[1][35] , \g_vector[1][33] ,
         \g_vector[1][31] , \g_vector[1][29] , \g_vector[1][27] ,
         \g_vector[1][25] , \g_vector[1][23] , \g_vector[1][21] ,
         \g_vector[1][19] , \g_vector[1][17] , \g_vector[1][15] ,
         \g_vector[1][13] , \g_vector[1][11] , \g_vector[1][9] ,
         \g_vector[1][7] , \g_vector[1][5] , \g_vector[1][3] ,
         \g_vector[1][1] , \g_vector[0][63] , \g_vector[0][62] ,
         \g_vector[0][61] , \g_vector[0][60] , \g_vector[0][59] ,
         \g_vector[0][58] , \g_vector[0][57] , \g_vector[0][56] ,
         \g_vector[0][55] , \g_vector[0][54] , \g_vector[0][53] ,
         \g_vector[0][52] , \g_vector[0][51] , \g_vector[0][50] ,
         \g_vector[0][49] , \g_vector[0][48] , \g_vector[0][47] ,
         \g_vector[0][46] , \g_vector[0][45] , \g_vector[0][44] ,
         \g_vector[0][43] , \g_vector[0][42] , \g_vector[0][41] ,
         \g_vector[0][40] , \g_vector[0][39] , \g_vector[0][38] ,
         \g_vector[0][37] , \g_vector[0][36] , \g_vector[0][35] ,
         \g_vector[0][34] , \g_vector[0][33] , \g_vector[0][32] ,
         \g_vector[0][31] , \g_vector[0][30] , \g_vector[0][29] ,
         \g_vector[0][28] , \g_vector[0][27] , \g_vector[0][26] ,
         \g_vector[0][25] , \g_vector[0][24] , \g_vector[0][23] ,
         \g_vector[0][22] , \g_vector[0][21] , \g_vector[0][20] ,
         \g_vector[0][19] , \g_vector[0][18] , \g_vector[0][17] ,
         \g_vector[0][16] , \g_vector[0][15] , \g_vector[0][14] ,
         \g_vector[0][13] , \g_vector[0][12] , \g_vector[0][11] ,
         \g_vector[0][10] , \g_vector[0][9] , \g_vector[0][8] ,
         \g_vector[0][7] , \g_vector[0][6] , \g_vector[0][5] ,
         \g_vector[0][4] , \g_vector[0][3] , \g_vector[0][2] ,
         \g_vector[0][1] , \g_vector[0][0] , \p_vector[5][63] ,
         \p_vector[5][59] , \p_vector[5][55] , \p_vector[5][51] ,
         \p_vector[4][63] , \p_vector[4][59] , \p_vector[4][47] ,
         \p_vector[4][43] , \p_vector[4][31] , \p_vector[4][27] ,
         \p_vector[3][63] , \p_vector[3][55] , \p_vector[3][47] ,
         \p_vector[3][39] , \p_vector[3][31] , \p_vector[3][23] ,
         \p_vector[3][15] , \p_vector[2][63] , \p_vector[2][59] ,
         \p_vector[2][55] , \p_vector[2][51] , \p_vector[2][47] ,
         \p_vector[2][43] , \p_vector[2][39] , \p_vector[2][35] ,
         \p_vector[2][31] , \p_vector[2][27] , \p_vector[2][23] ,
         \p_vector[2][19] , \p_vector[2][15] , \p_vector[2][11] ,
         \p_vector[2][7] , \p_vector[1][63] , \p_vector[1][61] ,
         \p_vector[1][59] , \p_vector[1][57] , \p_vector[1][55] ,
         \p_vector[1][53] , \p_vector[1][51] , \p_vector[1][49] ,
         \p_vector[1][47] , \p_vector[1][45] , \p_vector[1][43] ,
         \p_vector[1][41] , \p_vector[1][39] , \p_vector[1][37] ,
         \p_vector[1][35] , \p_vector[1][33] , \p_vector[1][31] ,
         \p_vector[1][29] , \p_vector[1][27] , \p_vector[1][25] ,
         \p_vector[1][23] , \p_vector[1][21] , \p_vector[1][19] ,
         \p_vector[1][17] , \p_vector[1][15] , \p_vector[1][13] ,
         \p_vector[1][11] , \p_vector[1][9] , \p_vector[1][7] ,
         \p_vector[1][5] , \p_vector[1][3] , \p_vector[0][63] ,
         \p_vector[0][62] , \p_vector[0][61] , \p_vector[0][60] ,
         \p_vector[0][59] , \p_vector[0][58] , \p_vector[0][57] ,
         \p_vector[0][56] , \p_vector[0][55] , \p_vector[0][54] ,
         \p_vector[0][53] , \p_vector[0][52] , \p_vector[0][51] ,
         \p_vector[0][50] , \p_vector[0][49] , \p_vector[0][48] ,
         \p_vector[0][47] , \p_vector[0][46] , \p_vector[0][45] ,
         \p_vector[0][44] , \p_vector[0][43] , \p_vector[0][42] ,
         \p_vector[0][41] , \p_vector[0][40] , \p_vector[0][39] ,
         \p_vector[0][38] , \p_vector[0][37] , \p_vector[0][36] ,
         \p_vector[0][35] , \p_vector[0][34] , \p_vector[0][33] ,
         \p_vector[0][32] , \p_vector[0][31] , \p_vector[0][30] ,
         \p_vector[0][29] , \p_vector[0][28] , \p_vector[0][27] ,
         \p_vector[0][26] , \p_vector[0][25] , \p_vector[0][24] ,
         \p_vector[0][23] , \p_vector[0][22] , \p_vector[0][21] ,
         \p_vector[0][20] , \p_vector[0][19] , \p_vector[0][18] ,
         \p_vector[0][17] , \p_vector[0][16] , \p_vector[0][15] ,
         \p_vector[0][14] , \p_vector[0][13] , \p_vector[0][12] ,
         \p_vector[0][11] , \p_vector[0][10] , \p_vector[0][9] ,
         \p_vector[0][8] , \p_vector[0][7] , \p_vector[0][6] ,
         \p_vector[0][5] , \p_vector[0][4] , \p_vector[0][3] ,
         \p_vector[0][2] , \p_vector[0][1] , n3, n1, n2;

  pg_net_189 pg_network_63 ( .a(A[63]), .b(B[63]), .p(\p_vector[0][63] ), .g(
        \g_vector[0][63] ) );
  pg_net_188 pg_network_62 ( .a(A[62]), .b(B[62]), .p(\p_vector[0][62] ), .g(
        \g_vector[0][62] ) );
  pg_net_187 pg_network_61 ( .a(A[61]), .b(B[61]), .p(\p_vector[0][61] ), .g(
        \g_vector[0][61] ) );
  pg_net_186 pg_network_60 ( .a(A[60]), .b(B[60]), .p(\p_vector[0][60] ), .g(
        \g_vector[0][60] ) );
  pg_net_185 pg_network_59 ( .a(A[59]), .b(B[59]), .p(\p_vector[0][59] ), .g(
        \g_vector[0][59] ) );
  pg_net_184 pg_network_58 ( .a(A[58]), .b(B[58]), .p(\p_vector[0][58] ), .g(
        \g_vector[0][58] ) );
  pg_net_183 pg_network_57 ( .a(A[57]), .b(B[57]), .p(\p_vector[0][57] ), .g(
        \g_vector[0][57] ) );
  pg_net_182 pg_network_56 ( .a(A[56]), .b(B[56]), .p(\p_vector[0][56] ), .g(
        \g_vector[0][56] ) );
  pg_net_181 pg_network_55 ( .a(A[55]), .b(B[55]), .p(\p_vector[0][55] ), .g(
        \g_vector[0][55] ) );
  pg_net_180 pg_network_54 ( .a(A[54]), .b(B[54]), .p(\p_vector[0][54] ), .g(
        \g_vector[0][54] ) );
  pg_net_179 pg_network_53 ( .a(A[53]), .b(B[53]), .p(\p_vector[0][53] ), .g(
        \g_vector[0][53] ) );
  pg_net_178 pg_network_52 ( .a(A[52]), .b(B[52]), .p(\p_vector[0][52] ), .g(
        \g_vector[0][52] ) );
  pg_net_177 pg_network_51 ( .a(A[51]), .b(B[51]), .p(\p_vector[0][51] ), .g(
        \g_vector[0][51] ) );
  pg_net_176 pg_network_50 ( .a(A[50]), .b(B[50]), .p(\p_vector[0][50] ), .g(
        \g_vector[0][50] ) );
  pg_net_175 pg_network_49 ( .a(A[49]), .b(B[49]), .p(\p_vector[0][49] ), .g(
        \g_vector[0][49] ) );
  pg_net_174 pg_network_48 ( .a(A[48]), .b(B[48]), .p(\p_vector[0][48] ), .g(
        \g_vector[0][48] ) );
  pg_net_173 pg_network_47 ( .a(A[47]), .b(B[47]), .p(\p_vector[0][47] ), .g(
        \g_vector[0][47] ) );
  pg_net_172 pg_network_46 ( .a(A[46]), .b(B[46]), .p(\p_vector[0][46] ), .g(
        \g_vector[0][46] ) );
  pg_net_171 pg_network_45 ( .a(A[45]), .b(B[45]), .p(\p_vector[0][45] ), .g(
        \g_vector[0][45] ) );
  pg_net_170 pg_network_44 ( .a(A[44]), .b(B[44]), .p(\p_vector[0][44] ), .g(
        \g_vector[0][44] ) );
  pg_net_169 pg_network_43 ( .a(A[43]), .b(B[43]), .p(\p_vector[0][43] ), .g(
        \g_vector[0][43] ) );
  pg_net_168 pg_network_42 ( .a(A[42]), .b(B[42]), .p(\p_vector[0][42] ), .g(
        \g_vector[0][42] ) );
  pg_net_167 pg_network_41 ( .a(A[41]), .b(B[41]), .p(\p_vector[0][41] ), .g(
        \g_vector[0][41] ) );
  pg_net_166 pg_network_40 ( .a(A[40]), .b(B[40]), .p(\p_vector[0][40] ), .g(
        \g_vector[0][40] ) );
  pg_net_165 pg_network_39 ( .a(A[39]), .b(B[39]), .p(\p_vector[0][39] ), .g(
        \g_vector[0][39] ) );
  pg_net_164 pg_network_38 ( .a(A[38]), .b(B[38]), .p(\p_vector[0][38] ), .g(
        \g_vector[0][38] ) );
  pg_net_163 pg_network_37 ( .a(A[37]), .b(B[37]), .p(\p_vector[0][37] ), .g(
        \g_vector[0][37] ) );
  pg_net_162 pg_network_36 ( .a(A[36]), .b(B[36]), .p(\p_vector[0][36] ), .g(
        \g_vector[0][36] ) );
  pg_net_161 pg_network_35 ( .a(A[35]), .b(B[35]), .p(\p_vector[0][35] ), .g(
        \g_vector[0][35] ) );
  pg_net_160 pg_network_34 ( .a(A[34]), .b(B[34]), .p(\p_vector[0][34] ), .g(
        \g_vector[0][34] ) );
  pg_net_159 pg_network_33 ( .a(A[33]), .b(B[33]), .p(\p_vector[0][33] ), .g(
        \g_vector[0][33] ) );
  pg_net_158 pg_network_32 ( .a(A[32]), .b(B[32]), .p(\p_vector[0][32] ), .g(
        \g_vector[0][32] ) );
  pg_net_157 pg_network_31 ( .a(A[31]), .b(B[31]), .p(\p_vector[0][31] ), .g(
        \g_vector[0][31] ) );
  pg_net_156 pg_network_30 ( .a(A[30]), .b(B[30]), .p(\p_vector[0][30] ), .g(
        \g_vector[0][30] ) );
  pg_net_155 pg_network_29 ( .a(A[29]), .b(B[29]), .p(\p_vector[0][29] ), .g(
        \g_vector[0][29] ) );
  pg_net_154 pg_network_28 ( .a(A[28]), .b(B[28]), .p(\p_vector[0][28] ), .g(
        \g_vector[0][28] ) );
  pg_net_153 pg_network_27 ( .a(A[27]), .b(B[27]), .p(\p_vector[0][27] ), .g(
        \g_vector[0][27] ) );
  pg_net_152 pg_network_26 ( .a(A[26]), .b(B[26]), .p(\p_vector[0][26] ), .g(
        \g_vector[0][26] ) );
  pg_net_151 pg_network_25 ( .a(A[25]), .b(B[25]), .p(\p_vector[0][25] ), .g(
        \g_vector[0][25] ) );
  pg_net_150 pg_network_24 ( .a(A[24]), .b(B[24]), .p(\p_vector[0][24] ), .g(
        \g_vector[0][24] ) );
  pg_net_149 pg_network_23 ( .a(A[23]), .b(B[23]), .p(\p_vector[0][23] ), .g(
        \g_vector[0][23] ) );
  pg_net_148 pg_network_22 ( .a(A[22]), .b(B[22]), .p(\p_vector[0][22] ), .g(
        \g_vector[0][22] ) );
  pg_net_147 pg_network_21 ( .a(A[21]), .b(B[21]), .p(\p_vector[0][21] ), .g(
        \g_vector[0][21] ) );
  pg_net_146 pg_network_20 ( .a(A[20]), .b(B[20]), .p(\p_vector[0][20] ), .g(
        \g_vector[0][20] ) );
  pg_net_145 pg_network_19 ( .a(A[19]), .b(B[19]), .p(\p_vector[0][19] ), .g(
        \g_vector[0][19] ) );
  pg_net_144 pg_network_18 ( .a(A[18]), .b(B[18]), .p(\p_vector[0][18] ), .g(
        \g_vector[0][18] ) );
  pg_net_143 pg_network_17 ( .a(A[17]), .b(B[17]), .p(\p_vector[0][17] ), .g(
        \g_vector[0][17] ) );
  pg_net_142 pg_network_16 ( .a(A[16]), .b(B[16]), .p(\p_vector[0][16] ), .g(
        \g_vector[0][16] ) );
  pg_net_141 pg_network_15 ( .a(A[15]), .b(B[15]), .p(\p_vector[0][15] ), .g(
        \g_vector[0][15] ) );
  pg_net_140 pg_network_14 ( .a(A[14]), .b(B[14]), .p(\p_vector[0][14] ), .g(
        \g_vector[0][14] ) );
  pg_net_139 pg_network_13 ( .a(A[13]), .b(B[13]), .p(\p_vector[0][13] ), .g(
        \g_vector[0][13] ) );
  pg_net_138 pg_network_12 ( .a(A[12]), .b(B[12]), .p(\p_vector[0][12] ), .g(
        \g_vector[0][12] ) );
  pg_net_137 pg_network_11 ( .a(A[11]), .b(B[11]), .p(\p_vector[0][11] ), .g(
        \g_vector[0][11] ) );
  pg_net_136 pg_network_10 ( .a(A[10]), .b(B[10]), .p(\p_vector[0][10] ), .g(
        \g_vector[0][10] ) );
  pg_net_135 pg_network_9 ( .a(A[9]), .b(B[9]), .p(\p_vector[0][9] ), .g(
        \g_vector[0][9] ) );
  pg_net_134 pg_network_8 ( .a(A[8]), .b(B[8]), .p(\p_vector[0][8] ), .g(
        \g_vector[0][8] ) );
  pg_net_133 pg_network_7 ( .a(A[7]), .b(B[7]), .p(\p_vector[0][7] ), .g(
        \g_vector[0][7] ) );
  pg_net_132 pg_network_6 ( .a(A[6]), .b(B[6]), .p(\p_vector[0][6] ), .g(
        \g_vector[0][6] ) );
  pg_net_131 pg_network_5 ( .a(A[5]), .b(B[5]), .p(\p_vector[0][5] ), .g(
        \g_vector[0][5] ) );
  pg_net_130 pg_network_4 ( .a(A[4]), .b(B[4]), .p(\p_vector[0][4] ), .g(
        \g_vector[0][4] ) );
  pg_net_129 pg_network_3 ( .a(A[3]), .b(B[3]), .p(\p_vector[0][3] ), .g(
        \g_vector[0][3] ) );
  pg_net_128 pg_network_2 ( .a(A[2]), .b(B[2]), .p(\p_vector[0][2] ), .g(
        \g_vector[0][2] ) );
  pg_net_127 pg_network_1 ( .a(A[1]), .b(B[1]), .p(\p_vector[0][1] ), .g(
        \g_vector[0][1] ) );
  PG_BLOCK_189 std_PG_1_63 ( .p2(\p_vector[0][63] ), .g2(\g_vector[0][63] ), 
        .p1(\p_vector[0][62] ), .g1(\g_vector[0][62] ), .PG_P(
        \p_vector[1][63] ), .PG_G(\g_vector[1][63] ) );
  PG_BLOCK_188 std_PG_1_61 ( .p2(\p_vector[0][61] ), .g2(\g_vector[0][61] ), 
        .p1(\p_vector[0][60] ), .g1(\g_vector[0][60] ), .PG_P(
        \p_vector[1][61] ), .PG_G(\g_vector[1][61] ) );
  PG_BLOCK_187 std_PG_1_59 ( .p2(\p_vector[0][59] ), .g2(\g_vector[0][59] ), 
        .p1(\p_vector[0][58] ), .g1(\g_vector[0][58] ), .PG_P(
        \p_vector[1][59] ), .PG_G(\g_vector[1][59] ) );
  PG_BLOCK_186 std_PG_1_57 ( .p2(\p_vector[0][57] ), .g2(\g_vector[0][57] ), 
        .p1(\p_vector[0][56] ), .g1(\g_vector[0][56] ), .PG_P(
        \p_vector[1][57] ), .PG_G(\g_vector[1][57] ) );
  PG_BLOCK_185 std_PG_1_55 ( .p2(\p_vector[0][55] ), .g2(\g_vector[0][55] ), 
        .p1(\p_vector[0][54] ), .g1(\g_vector[0][54] ), .PG_P(
        \p_vector[1][55] ), .PG_G(\g_vector[1][55] ) );
  PG_BLOCK_184 std_PG_1_53 ( .p2(\p_vector[0][53] ), .g2(\g_vector[0][53] ), 
        .p1(\p_vector[0][52] ), .g1(\g_vector[0][52] ), .PG_P(
        \p_vector[1][53] ), .PG_G(\g_vector[1][53] ) );
  PG_BLOCK_183 std_PG_1_51 ( .p2(\p_vector[0][51] ), .g2(\g_vector[0][51] ), 
        .p1(\p_vector[0][50] ), .g1(\g_vector[0][50] ), .PG_P(
        \p_vector[1][51] ), .PG_G(\g_vector[1][51] ) );
  PG_BLOCK_182 std_PG_1_49 ( .p2(\p_vector[0][49] ), .g2(\g_vector[0][49] ), 
        .p1(\p_vector[0][48] ), .g1(\g_vector[0][48] ), .PG_P(
        \p_vector[1][49] ), .PG_G(\g_vector[1][49] ) );
  PG_BLOCK_181 std_PG_1_47 ( .p2(\p_vector[0][47] ), .g2(\g_vector[0][47] ), 
        .p1(\p_vector[0][46] ), .g1(\g_vector[0][46] ), .PG_P(
        \p_vector[1][47] ), .PG_G(\g_vector[1][47] ) );
  PG_BLOCK_180 std_PG_1_45 ( .p2(\p_vector[0][45] ), .g2(\g_vector[0][45] ), 
        .p1(\p_vector[0][44] ), .g1(\g_vector[0][44] ), .PG_P(
        \p_vector[1][45] ), .PG_G(\g_vector[1][45] ) );
  PG_BLOCK_179 std_PG_1_43 ( .p2(\p_vector[0][43] ), .g2(\g_vector[0][43] ), 
        .p1(\p_vector[0][42] ), .g1(\g_vector[0][42] ), .PG_P(
        \p_vector[1][43] ), .PG_G(\g_vector[1][43] ) );
  PG_BLOCK_178 std_PG_1_41 ( .p2(\p_vector[0][41] ), .g2(\g_vector[0][41] ), 
        .p1(\p_vector[0][40] ), .g1(\g_vector[0][40] ), .PG_P(
        \p_vector[1][41] ), .PG_G(\g_vector[1][41] ) );
  PG_BLOCK_177 std_PG_1_39 ( .p2(\p_vector[0][39] ), .g2(\g_vector[0][39] ), 
        .p1(\p_vector[0][38] ), .g1(\g_vector[0][38] ), .PG_P(
        \p_vector[1][39] ), .PG_G(\g_vector[1][39] ) );
  PG_BLOCK_176 std_PG_1_37 ( .p2(\p_vector[0][37] ), .g2(\g_vector[0][37] ), 
        .p1(\p_vector[0][36] ), .g1(\g_vector[0][36] ), .PG_P(
        \p_vector[1][37] ), .PG_G(\g_vector[1][37] ) );
  PG_BLOCK_175 std_PG_1_35 ( .p2(\p_vector[0][35] ), .g2(\g_vector[0][35] ), 
        .p1(\p_vector[0][34] ), .g1(\g_vector[0][34] ), .PG_P(
        \p_vector[1][35] ), .PG_G(\g_vector[1][35] ) );
  PG_BLOCK_174 std_PG_1_33 ( .p2(\p_vector[0][33] ), .g2(\g_vector[0][33] ), 
        .p1(\p_vector[0][32] ), .g1(\g_vector[0][32] ), .PG_P(
        \p_vector[1][33] ), .PG_G(\g_vector[1][33] ) );
  PG_BLOCK_173 std_PG_1_31 ( .p2(\p_vector[0][31] ), .g2(\g_vector[0][31] ), 
        .p1(\p_vector[0][30] ), .g1(\g_vector[0][30] ), .PG_P(
        \p_vector[1][31] ), .PG_G(\g_vector[1][31] ) );
  PG_BLOCK_172 std_PG_1_29 ( .p2(\p_vector[0][29] ), .g2(\g_vector[0][29] ), 
        .p1(\p_vector[0][28] ), .g1(\g_vector[0][28] ), .PG_P(
        \p_vector[1][29] ), .PG_G(\g_vector[1][29] ) );
  PG_BLOCK_171 std_PG_1_27 ( .p2(\p_vector[0][27] ), .g2(\g_vector[0][27] ), 
        .p1(\p_vector[0][26] ), .g1(\g_vector[0][26] ), .PG_P(
        \p_vector[1][27] ), .PG_G(\g_vector[1][27] ) );
  PG_BLOCK_170 std_PG_1_25 ( .p2(\p_vector[0][25] ), .g2(\g_vector[0][25] ), 
        .p1(\p_vector[0][24] ), .g1(\g_vector[0][24] ), .PG_P(
        \p_vector[1][25] ), .PG_G(\g_vector[1][25] ) );
  PG_BLOCK_169 std_PG_1_23 ( .p2(\p_vector[0][23] ), .g2(\g_vector[0][23] ), 
        .p1(\p_vector[0][22] ), .g1(\g_vector[0][22] ), .PG_P(
        \p_vector[1][23] ), .PG_G(\g_vector[1][23] ) );
  PG_BLOCK_168 std_PG_1_21 ( .p2(\p_vector[0][21] ), .g2(\g_vector[0][21] ), 
        .p1(\p_vector[0][20] ), .g1(\g_vector[0][20] ), .PG_P(
        \p_vector[1][21] ), .PG_G(\g_vector[1][21] ) );
  PG_BLOCK_167 std_PG_1_19 ( .p2(\p_vector[0][19] ), .g2(\g_vector[0][19] ), 
        .p1(\p_vector[0][18] ), .g1(\g_vector[0][18] ), .PG_P(
        \p_vector[1][19] ), .PG_G(\g_vector[1][19] ) );
  PG_BLOCK_166 std_PG_1_17 ( .p2(\p_vector[0][17] ), .g2(\g_vector[0][17] ), 
        .p1(\p_vector[0][16] ), .g1(\g_vector[0][16] ), .PG_P(
        \p_vector[1][17] ), .PG_G(\g_vector[1][17] ) );
  PG_BLOCK_165 std_PG_1_15 ( .p2(\p_vector[0][15] ), .g2(\g_vector[0][15] ), 
        .p1(\p_vector[0][14] ), .g1(\g_vector[0][14] ), .PG_P(
        \p_vector[1][15] ), .PG_G(\g_vector[1][15] ) );
  PG_BLOCK_164 std_PG_1_13 ( .p2(\p_vector[0][13] ), .g2(\g_vector[0][13] ), 
        .p1(\p_vector[0][12] ), .g1(\g_vector[0][12] ), .PG_P(
        \p_vector[1][13] ), .PG_G(\g_vector[1][13] ) );
  PG_BLOCK_163 std_PG_1_11 ( .p2(\p_vector[0][11] ), .g2(\g_vector[0][11] ), 
        .p1(\p_vector[0][10] ), .g1(\g_vector[0][10] ), .PG_P(
        \p_vector[1][11] ), .PG_G(\g_vector[1][11] ) );
  PG_BLOCK_162 std_PG_1_9 ( .p2(\p_vector[0][9] ), .g2(\g_vector[0][9] ), .p1(
        \p_vector[0][8] ), .g1(\g_vector[0][8] ), .PG_P(\p_vector[1][9] ), 
        .PG_G(\g_vector[1][9] ) );
  PG_BLOCK_161 std_PG_1_7 ( .p2(\p_vector[0][7] ), .g2(\g_vector[0][7] ), .p1(
        \p_vector[0][6] ), .g1(\g_vector[0][6] ), .PG_P(\p_vector[1][7] ), 
        .PG_G(\g_vector[1][7] ) );
  PG_BLOCK_160 std_PG_1_5 ( .p2(\p_vector[0][5] ), .g2(\g_vector[0][5] ), .p1(
        \p_vector[0][4] ), .g1(\g_vector[0][4] ), .PG_P(\p_vector[1][5] ), 
        .PG_G(\g_vector[1][5] ) );
  PG_BLOCK_159 std_PG_1_3 ( .p2(\p_vector[0][3] ), .g2(\g_vector[0][3] ), .p1(
        \p_vector[0][2] ), .g1(\g_vector[0][2] ), .PG_P(\p_vector[1][3] ), 
        .PG_G(\g_vector[1][3] ) );
  G_BLOCK_51 std_G_1_1 ( .p2(\p_vector[0][1] ), .g2(\g_vector[0][1] ), .g1(
        \g_vector[0][0] ), .G(\g_vector[1][1] ) );
  PG_BLOCK_158 std_PG_2_63 ( .p2(\p_vector[1][63] ), .g2(\g_vector[1][63] ), 
        .p1(\p_vector[1][61] ), .g1(\g_vector[1][61] ), .PG_P(
        \p_vector[2][63] ), .PG_G(\g_vector[2][63] ) );
  PG_BLOCK_157 std_PG_2_59 ( .p2(\p_vector[1][59] ), .g2(\g_vector[1][59] ), 
        .p1(\p_vector[1][57] ), .g1(\g_vector[1][57] ), .PG_P(
        \p_vector[2][59] ), .PG_G(\g_vector[2][59] ) );
  PG_BLOCK_156 std_PG_2_55 ( .p2(\p_vector[1][55] ), .g2(\g_vector[1][55] ), 
        .p1(\p_vector[1][53] ), .g1(\g_vector[1][53] ), .PG_P(
        \p_vector[2][55] ), .PG_G(\g_vector[2][55] ) );
  PG_BLOCK_155 std_PG_2_51 ( .p2(\p_vector[1][51] ), .g2(\g_vector[1][51] ), 
        .p1(\p_vector[1][49] ), .g1(\g_vector[1][49] ), .PG_P(
        \p_vector[2][51] ), .PG_G(\g_vector[2][51] ) );
  PG_BLOCK_154 std_PG_2_47 ( .p2(\p_vector[1][47] ), .g2(\g_vector[1][47] ), 
        .p1(\p_vector[1][45] ), .g1(\g_vector[1][45] ), .PG_P(
        \p_vector[2][47] ), .PG_G(\g_vector[2][47] ) );
  PG_BLOCK_153 std_PG_2_43 ( .p2(\p_vector[1][43] ), .g2(\g_vector[1][43] ), 
        .p1(\p_vector[1][41] ), .g1(\g_vector[1][41] ), .PG_P(
        \p_vector[2][43] ), .PG_G(\g_vector[2][43] ) );
  PG_BLOCK_152 std_PG_2_39 ( .p2(\p_vector[1][39] ), .g2(\g_vector[1][39] ), 
        .p1(\p_vector[1][37] ), .g1(\g_vector[1][37] ), .PG_P(
        \p_vector[2][39] ), .PG_G(\g_vector[2][39] ) );
  PG_BLOCK_151 std_PG_2_35 ( .p2(\p_vector[1][35] ), .g2(\g_vector[1][35] ), 
        .p1(\p_vector[1][33] ), .g1(\g_vector[1][33] ), .PG_P(
        \p_vector[2][35] ), .PG_G(\g_vector[2][35] ) );
  PG_BLOCK_150 std_PG_2_31 ( .p2(\p_vector[1][31] ), .g2(\g_vector[1][31] ), 
        .p1(\p_vector[1][29] ), .g1(\g_vector[1][29] ), .PG_P(
        \p_vector[2][31] ), .PG_G(\g_vector[2][31] ) );
  PG_BLOCK_149 std_PG_2_27 ( .p2(\p_vector[1][27] ), .g2(\g_vector[1][27] ), 
        .p1(\p_vector[1][25] ), .g1(\g_vector[1][25] ), .PG_P(
        \p_vector[2][27] ), .PG_G(\g_vector[2][27] ) );
  PG_BLOCK_148 std_PG_2_23 ( .p2(\p_vector[1][23] ), .g2(\g_vector[1][23] ), 
        .p1(\p_vector[1][21] ), .g1(\g_vector[1][21] ), .PG_P(
        \p_vector[2][23] ), .PG_G(\g_vector[2][23] ) );
  PG_BLOCK_147 std_PG_2_19 ( .p2(\p_vector[1][19] ), .g2(\g_vector[1][19] ), 
        .p1(\p_vector[1][17] ), .g1(\g_vector[1][17] ), .PG_P(
        \p_vector[2][19] ), .PG_G(\g_vector[2][19] ) );
  PG_BLOCK_146 std_PG_2_15 ( .p2(\p_vector[1][15] ), .g2(\g_vector[1][15] ), 
        .p1(\p_vector[1][13] ), .g1(\g_vector[1][13] ), .PG_P(
        \p_vector[2][15] ), .PG_G(\g_vector[2][15] ) );
  PG_BLOCK_145 std_PG_2_11 ( .p2(\p_vector[1][11] ), .g2(\g_vector[1][11] ), 
        .p1(\p_vector[1][9] ), .g1(\g_vector[1][9] ), .PG_P(\p_vector[2][11] ), 
        .PG_G(\g_vector[2][11] ) );
  PG_BLOCK_144 std_PG_2_7 ( .p2(\p_vector[1][7] ), .g2(\g_vector[1][7] ), .p1(
        \p_vector[1][5] ), .g1(\g_vector[1][5] ), .PG_P(\p_vector[2][7] ), 
        .PG_G(\g_vector[2][7] ) );
  G_BLOCK_50 std_G_2_3 ( .p2(\p_vector[1][3] ), .g2(\g_vector[1][3] ), .g1(
        \g_vector[1][1] ), .G(Co[0]) );
  PG_BLOCK_143 std_PG_3_63 ( .p2(\p_vector[2][63] ), .g2(\g_vector[2][63] ), 
        .p1(\p_vector[2][59] ), .g1(\g_vector[2][59] ), .PG_P(
        \p_vector[3][63] ), .PG_G(\g_vector[3][63] ) );
  PG_BLOCK_142 std_PG_3_55 ( .p2(\p_vector[2][55] ), .g2(\g_vector[2][55] ), 
        .p1(\p_vector[2][51] ), .g1(\g_vector[2][51] ), .PG_P(
        \p_vector[3][55] ), .PG_G(\g_vector[3][55] ) );
  PG_BLOCK_141 std_PG_3_47 ( .p2(\p_vector[2][47] ), .g2(\g_vector[2][47] ), 
        .p1(\p_vector[2][43] ), .g1(\g_vector[2][43] ), .PG_P(
        \p_vector[3][47] ), .PG_G(\g_vector[3][47] ) );
  PG_BLOCK_140 std_PG_3_39 ( .p2(\p_vector[2][39] ), .g2(\g_vector[2][39] ), 
        .p1(\p_vector[2][35] ), .g1(\g_vector[2][35] ), .PG_P(
        \p_vector[3][39] ), .PG_G(\g_vector[3][39] ) );
  PG_BLOCK_139 std_PG_3_31 ( .p2(\p_vector[2][31] ), .g2(\g_vector[2][31] ), 
        .p1(\p_vector[2][27] ), .g1(\g_vector[2][27] ), .PG_P(
        \p_vector[3][31] ), .PG_G(\g_vector[3][31] ) );
  PG_BLOCK_138 std_PG_3_23 ( .p2(\p_vector[2][23] ), .g2(\g_vector[2][23] ), 
        .p1(\p_vector[2][19] ), .g1(\g_vector[2][19] ), .PG_P(
        \p_vector[3][23] ), .PG_G(\g_vector[3][23] ) );
  PG_BLOCK_137 std_PG_3_15 ( .p2(\p_vector[2][15] ), .g2(\g_vector[2][15] ), 
        .p1(\p_vector[2][11] ), .g1(\g_vector[2][11] ), .PG_P(
        \p_vector[3][15] ), .PG_G(\g_vector[3][15] ) );
  G_BLOCK_49 std_G_3_7 ( .p2(\p_vector[2][7] ), .g2(\g_vector[2][7] ), .g1(
        Co[0]), .G(Co[1]) );
  PG_BLOCK_136 std_PG_4_63 ( .p2(\p_vector[3][63] ), .g2(\g_vector[3][63] ), 
        .p1(\p_vector[3][55] ), .g1(\g_vector[3][55] ), .PG_P(
        \p_vector[4][63] ), .PG_G(\g_vector[4][63] ) );
  PG_BLOCK_135 add_PG_4_63_1 ( .p2(\p_vector[2][59] ), .g2(\g_vector[2][59] ), 
        .p1(\p_vector[3][55] ), .g1(\g_vector[3][55] ), .PG_P(
        \p_vector[4][59] ), .PG_G(\g_vector[4][59] ) );
  PG_BLOCK_134 std_PG_4_47 ( .p2(\p_vector[3][47] ), .g2(\g_vector[3][47] ), 
        .p1(\p_vector[3][39] ), .g1(\g_vector[3][39] ), .PG_P(
        \p_vector[4][47] ), .PG_G(\g_vector[4][47] ) );
  PG_BLOCK_133 add_PG_4_47_1 ( .p2(\p_vector[2][43] ), .g2(\g_vector[2][43] ), 
        .p1(\p_vector[3][39] ), .g1(\g_vector[3][39] ), .PG_P(
        \p_vector[4][43] ), .PG_G(\g_vector[4][43] ) );
  PG_BLOCK_132 std_PG_4_31 ( .p2(\p_vector[3][31] ), .g2(\g_vector[3][31] ), 
        .p1(\p_vector[3][23] ), .g1(\g_vector[3][23] ), .PG_P(
        \p_vector[4][31] ), .PG_G(\g_vector[4][31] ) );
  PG_BLOCK_131 add_PG_4_31_1 ( .p2(\p_vector[2][27] ), .g2(\g_vector[2][27] ), 
        .p1(\p_vector[3][23] ), .g1(\g_vector[3][23] ), .PG_P(
        \p_vector[4][27] ), .PG_G(\g_vector[4][27] ) );
  G_BLOCK_48 std_G_4_15 ( .p2(\p_vector[3][15] ), .g2(\g_vector[3][15] ), .g1(
        Co[1]), .G(Co[3]) );
  G_BLOCK_47 add_G_4_15_1 ( .p2(\p_vector[2][11] ), .g2(\g_vector[2][11] ), 
        .g1(Co[1]), .G(Co[2]) );
  PG_BLOCK_130 std_PG_5_63 ( .p2(\p_vector[4][63] ), .g2(\g_vector[4][63] ), 
        .p1(\p_vector[4][47] ), .g1(\g_vector[4][47] ), .PG_P(
        \p_vector[5][63] ), .PG_G(\g_vector[5][63] ) );
  PG_BLOCK_129 add_PG_5_63_1 ( .p2(\p_vector[4][59] ), .g2(\g_vector[4][59] ), 
        .p1(\p_vector[4][47] ), .g1(\g_vector[4][47] ), .PG_P(
        \p_vector[5][59] ), .PG_G(\g_vector[5][59] ) );
  PG_BLOCK_128 add_PG_5_63_2 ( .p2(\p_vector[3][55] ), .g2(\g_vector[3][55] ), 
        .p1(\p_vector[4][47] ), .g1(\g_vector[4][47] ), .PG_P(
        \p_vector[5][55] ), .PG_G(\g_vector[5][55] ) );
  PG_BLOCK_127 add_PG_5_63_3 ( .p2(\p_vector[2][51] ), .g2(\g_vector[2][51] ), 
        .p1(\p_vector[4][47] ), .g1(\g_vector[4][47] ), .PG_P(
        \p_vector[5][51] ), .PG_G(\g_vector[5][51] ) );
  G_BLOCK_46 std_G_5_31 ( .p2(\p_vector[4][31] ), .g2(\g_vector[4][31] ), .g1(
        Co[3]), .G(Co[7]) );
  G_BLOCK_45 add_G_5_31_1 ( .p2(\p_vector[4][27] ), .g2(\g_vector[4][27] ), 
        .g1(Co[3]), .G(Co[6]) );
  G_BLOCK_44 add_G_5_31_2 ( .p2(\p_vector[3][23] ), .g2(\g_vector[3][23] ), 
        .g1(Co[3]), .G(Co[5]) );
  G_BLOCK_43 add_G_5_31_3 ( .p2(\p_vector[2][19] ), .g2(\g_vector[2][19] ), 
        .g1(Co[3]), .G(Co[4]) );
  G_BLOCK_42 std_G_6_63 ( .p2(\p_vector[5][63] ), .g2(\g_vector[5][63] ), .g1(
        Co[7]), .G(Co[15]) );
  G_BLOCK_41 add_G_6_63_1 ( .p2(\p_vector[5][59] ), .g2(\g_vector[5][59] ), 
        .g1(Co[7]), .G(Co[14]) );
  G_BLOCK_40 add_G_6_63_2 ( .p2(\p_vector[5][55] ), .g2(\g_vector[5][55] ), 
        .g1(Co[7]), .G(Co[13]) );
  G_BLOCK_39 add_G_6_63_3 ( .p2(\p_vector[5][51] ), .g2(\g_vector[5][51] ), 
        .g1(Co[7]), .G(Co[12]) );
  G_BLOCK_38 add_G_6_63_4 ( .p2(\p_vector[4][47] ), .g2(\g_vector[4][47] ), 
        .g1(Co[7]), .G(Co[11]) );
  G_BLOCK_37 add_G_6_63_5 ( .p2(\p_vector[4][43] ), .g2(\g_vector[4][43] ), 
        .g1(Co[7]), .G(Co[10]) );
  G_BLOCK_36 add_G_6_63_6 ( .p2(\p_vector[3][39] ), .g2(\g_vector[3][39] ), 
        .g1(Co[7]), .G(Co[9]) );
  G_BLOCK_35 add_G_6_63_7 ( .p2(\p_vector[2][35] ), .g2(\g_vector[2][35] ), 
        .g1(Co[7]), .G(Co[8]) );
  OAI21_X1 U1 ( .B1(n2), .B2(n1), .A(n3), .ZN(\g_vector[0][0] ) );
  OAI21_X1 U2 ( .B1(A[0]), .B2(B[0]), .A(Cin), .ZN(n3) );
  INV_X1 U3 ( .A(A[0]), .ZN(n2) );
  INV_X1 U4 ( .A(B[0]), .ZN(n1) );
endmodule


module FA_384 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_383 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_382 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_381 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_96 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_384 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_383 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_382 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_381 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_380 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_379 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_378 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_377 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_95 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_380 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_379 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_378 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_377 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_192 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_191 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_190 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_189 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_GENERIC_NBIT4_48 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_192 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_191 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_190 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_189 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_48 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_96 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_95 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_48 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module FA_376 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_375 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_374 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_373 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_94 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_376 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_375 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_374 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_373 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_372 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_371 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_370 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_369 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_93 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_372 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_371 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_370 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_369 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_188 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_187 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_186 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_185 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_GENERIC_NBIT4_47 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_188 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_187 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_186 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_185 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_47 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_94 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_93 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_47 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module FA_368 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_367 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_366 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_365 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_92 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_368 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_367 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_366 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_365 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_364 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_363 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_362 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_361 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_91 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_364 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_363 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_362 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_361 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_184 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_183 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_182 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_181 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_GENERIC_NBIT4_46 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_184 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_183 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_182 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_181 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_46 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_92 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_91 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_46 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module FA_360 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_359 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_358 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_357 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_90 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_360 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_359 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_358 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_357 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_356 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_355 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_354 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_353 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_89 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_356 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_355 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_354 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_353 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_180 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_179 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_178 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_177 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_GENERIC_NBIT4_45 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_180 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_179 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_178 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_177 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_45 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_90 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_89 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_45 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module FA_352 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_351 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_350 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_349 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_88 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_352 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_351 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_350 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_349 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_348 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_347 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_346 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_345 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_87 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_348 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_347 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_346 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_345 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_176 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_175 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_174 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_173 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_GENERIC_NBIT4_44 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_176 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_175 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_174 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_173 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_44 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_88 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_87 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_44 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module FA_344 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_343 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_342 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_341 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_86 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_344 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_343 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_342 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_341 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_340 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_339 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_338 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_337 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_85 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_340 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_339 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_338 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_337 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_172 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_171 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_170 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_169 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_GENERIC_NBIT4_43 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_172 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_171 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_170 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_169 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_43 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_86 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_85 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_43 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module FA_336 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_335 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_334 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_333 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_84 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_336 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_335 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_334 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_333 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_332 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_331 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_330 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_329 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_83 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_332 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_331 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_330 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_329 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_168 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_167 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_166 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_165 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_GENERIC_NBIT4_42 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_168 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_167 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_166 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_165 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_42 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_84 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_83 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_42 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module FA_328 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_327 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_326 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_325 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_82 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_328 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_327 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_326 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_325 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_324 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_323 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_322 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_321 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_81 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_324 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_323 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_322 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_321 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_164 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_163 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_162 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_161 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_GENERIC_NBIT4_41 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_164 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_163 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_162 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_161 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_41 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_82 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_81 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_41 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module FA_320 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_319 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_318 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_317 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_80 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_320 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_319 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_318 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_317 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_316 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_315 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_314 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_313 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_79 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_316 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_315 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_314 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_313 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_160 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_159 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_158 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_157 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_GENERIC_NBIT4_40 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_160 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_159 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_158 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_157 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_40 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_80 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_79 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_40 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module FA_312 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_311 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_310 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_309 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_78 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_312 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_311 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_310 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_309 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_308 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_307 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_306 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_305 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_77 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_308 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_307 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_306 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_305 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_156 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_155 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_154 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_153 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_GENERIC_NBIT4_39 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_156 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_155 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_154 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_153 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_39 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_78 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_77 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_39 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module FA_304 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_303 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_302 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_301 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_76 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_304 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_303 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_302 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_301 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_300 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_299 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_298 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_297 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_75 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_300 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_299 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_298 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_297 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_152 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_151 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_150 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_149 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_GENERIC_NBIT4_38 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_152 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_151 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_150 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_149 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_38 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_76 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_75 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_38 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module FA_296 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_295 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_294 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_293 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_74 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_296 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_295 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_294 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_293 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_292 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_291 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_290 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_289 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_73 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_292 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_291 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_290 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_289 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_148 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_147 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_146 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_145 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_GENERIC_NBIT4_37 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_148 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_147 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_146 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_145 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_37 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_74 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_73 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_37 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module FA_288 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_287 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_286 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_285 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_72 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_288 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_287 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_286 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_285 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_284 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_283 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_282 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_281 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_71 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_284 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_283 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_282 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_281 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_144 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_143 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_142 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_141 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_GENERIC_NBIT4_36 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_144 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_143 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_142 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_141 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_36 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_72 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_71 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_36 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module FA_280 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_279 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_278 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_277 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_70 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_280 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_279 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_278 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_277 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_276 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_275 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_274 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_273 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_69 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_276 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_275 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_274 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_273 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_140 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_139 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_138 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_137 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_GENERIC_NBIT4_35 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_140 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_139 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_138 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_137 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_35 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_70 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_69 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_35 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module FA_272 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_271 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_270 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_269 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_68 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_272 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_271 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_270 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_269 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_268 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_267 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_266 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_265 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_67 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_268 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_267 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_266 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_265 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_136 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_135 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_134 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_133 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_GENERIC_NBIT4_34 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_136 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_135 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_134 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_133 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_34 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_68 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_67 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_34 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module FA_264 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_263 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_262 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_261 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_66 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_264 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_263 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_262 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_261 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_260 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_259 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_258 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_257 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_65 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_260 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_259 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_258 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_257 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_132 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_131 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_130 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_129 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_GENERIC_NBIT4_33 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_132 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_131 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_130 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_129 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_33 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_66 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_65 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_33 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module sum_generator_n_bit64_n_CSB16_0 ( A, B, C_in, S );
  input [63:0] A;
  input [63:0] B;
  input [15:0] C_in;
  output [63:0] S;


  carry_select_block_n4_48 csb_0 ( .A(A[3:0]), .B(B[3:0]), .C_sel(C_in[0]), 
        .S(S[3:0]) );
  carry_select_block_n4_47 csb_1 ( .A(A[7:4]), .B(B[7:4]), .C_sel(C_in[1]), 
        .S(S[7:4]) );
  carry_select_block_n4_46 csb_2 ( .A(A[11:8]), .B(B[11:8]), .C_sel(C_in[2]), 
        .S(S[11:8]) );
  carry_select_block_n4_45 csb_3 ( .A(A[15:12]), .B(B[15:12]), .C_sel(C_in[3]), 
        .S(S[15:12]) );
  carry_select_block_n4_44 csb_4 ( .A(A[19:16]), .B(B[19:16]), .C_sel(C_in[4]), 
        .S(S[19:16]) );
  carry_select_block_n4_43 csb_5 ( .A(A[23:20]), .B(B[23:20]), .C_sel(C_in[5]), 
        .S(S[23:20]) );
  carry_select_block_n4_42 csb_6 ( .A(A[27:24]), .B(B[27:24]), .C_sel(C_in[6]), 
        .S(S[27:24]) );
  carry_select_block_n4_41 csb_7 ( .A(A[31:28]), .B(B[31:28]), .C_sel(C_in[7]), 
        .S(S[31:28]) );
  carry_select_block_n4_40 csb_8 ( .A(A[35:32]), .B(B[35:32]), .C_sel(C_in[8]), 
        .S(S[35:32]) );
  carry_select_block_n4_39 csb_9 ( .A(A[39:36]), .B(B[39:36]), .C_sel(C_in[9]), 
        .S(S[39:36]) );
  carry_select_block_n4_38 csb_10 ( .A(A[43:40]), .B(B[43:40]), .C_sel(
        C_in[10]), .S(S[43:40]) );
  carry_select_block_n4_37 csb_11 ( .A(A[47:44]), .B(B[47:44]), .C_sel(
        C_in[11]), .S(S[47:44]) );
  carry_select_block_n4_36 csb_12 ( .A(A[51:48]), .B(B[51:48]), .C_sel(
        C_in[12]), .S(S[51:48]) );
  carry_select_block_n4_35 csb_13 ( .A(A[55:52]), .B(B[55:52]), .C_sel(
        C_in[13]), .S(S[55:52]) );
  carry_select_block_n4_34 csb_14 ( .A(A[59:56]), .B(B[59:56]), .C_sel(
        C_in[14]), .S(S[59:56]) );
  carry_select_block_n4_33 csb_15 ( .A(A[63:60]), .B(B[63:60]), .C_sel(
        C_in[15]), .S(S[63:60]) );
endmodule


module P4_ADDER_NBIT64_0 ( A, B, Cin, S, Cout, ovf );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Cin;
  output Cout, ovf;
  wire   n1, n2;
  wire   [63:0] xor_b;
  wire   [14:0] carry;

  XOR2_X1 U3 ( .A(xor_b[63]), .B(A[63]), .Z(n2) );
  my_xor_192 bc_xor_63 ( .A(B[63]), .B(Cin), .xor_out(xor_b[63]) );
  my_xor_191 bc_xor_62 ( .A(B[62]), .B(Cin), .xor_out(xor_b[62]) );
  my_xor_190 bc_xor_61 ( .A(B[61]), .B(Cin), .xor_out(xor_b[61]) );
  my_xor_189 bc_xor_60 ( .A(B[60]), .B(Cin), .xor_out(xor_b[60]) );
  my_xor_188 bc_xor_59 ( .A(B[59]), .B(Cin), .xor_out(xor_b[59]) );
  my_xor_187 bc_xor_58 ( .A(B[58]), .B(Cin), .xor_out(xor_b[58]) );
  my_xor_186 bc_xor_57 ( .A(B[57]), .B(Cin), .xor_out(xor_b[57]) );
  my_xor_185 bc_xor_56 ( .A(B[56]), .B(Cin), .xor_out(xor_b[56]) );
  my_xor_184 bc_xor_55 ( .A(B[55]), .B(Cin), .xor_out(xor_b[55]) );
  my_xor_183 bc_xor_54 ( .A(B[54]), .B(Cin), .xor_out(xor_b[54]) );
  my_xor_182 bc_xor_53 ( .A(B[53]), .B(Cin), .xor_out(xor_b[53]) );
  my_xor_181 bc_xor_52 ( .A(B[52]), .B(Cin), .xor_out(xor_b[52]) );
  my_xor_180 bc_xor_51 ( .A(B[51]), .B(Cin), .xor_out(xor_b[51]) );
  my_xor_179 bc_xor_50 ( .A(B[50]), .B(Cin), .xor_out(xor_b[50]) );
  my_xor_178 bc_xor_49 ( .A(B[49]), .B(Cin), .xor_out(xor_b[49]) );
  my_xor_177 bc_xor_48 ( .A(B[48]), .B(Cin), .xor_out(xor_b[48]) );
  my_xor_176 bc_xor_47 ( .A(B[47]), .B(Cin), .xor_out(xor_b[47]) );
  my_xor_175 bc_xor_46 ( .A(B[46]), .B(Cin), .xor_out(xor_b[46]) );
  my_xor_174 bc_xor_45 ( .A(B[45]), .B(Cin), .xor_out(xor_b[45]) );
  my_xor_173 bc_xor_44 ( .A(B[44]), .B(Cin), .xor_out(xor_b[44]) );
  my_xor_172 bc_xor_43 ( .A(B[43]), .B(Cin), .xor_out(xor_b[43]) );
  my_xor_171 bc_xor_42 ( .A(B[42]), .B(Cin), .xor_out(xor_b[42]) );
  my_xor_170 bc_xor_41 ( .A(B[41]), .B(Cin), .xor_out(xor_b[41]) );
  my_xor_169 bc_xor_40 ( .A(B[40]), .B(Cin), .xor_out(xor_b[40]) );
  my_xor_168 bc_xor_39 ( .A(B[39]), .B(Cin), .xor_out(xor_b[39]) );
  my_xor_167 bc_xor_38 ( .A(B[38]), .B(Cin), .xor_out(xor_b[38]) );
  my_xor_166 bc_xor_37 ( .A(B[37]), .B(Cin), .xor_out(xor_b[37]) );
  my_xor_165 bc_xor_36 ( .A(B[36]), .B(Cin), .xor_out(xor_b[36]) );
  my_xor_164 bc_xor_35 ( .A(B[35]), .B(Cin), .xor_out(xor_b[35]) );
  my_xor_163 bc_xor_34 ( .A(B[34]), .B(Cin), .xor_out(xor_b[34]) );
  my_xor_162 bc_xor_33 ( .A(B[33]), .B(Cin), .xor_out(xor_b[33]) );
  my_xor_161 bc_xor_32 ( .A(B[32]), .B(Cin), .xor_out(xor_b[32]) );
  my_xor_160 bc_xor_31 ( .A(B[31]), .B(Cin), .xor_out(xor_b[31]) );
  my_xor_159 bc_xor_30 ( .A(B[30]), .B(Cin), .xor_out(xor_b[30]) );
  my_xor_158 bc_xor_29 ( .A(B[29]), .B(Cin), .xor_out(xor_b[29]) );
  my_xor_157 bc_xor_28 ( .A(B[28]), .B(Cin), .xor_out(xor_b[28]) );
  my_xor_156 bc_xor_27 ( .A(B[27]), .B(Cin), .xor_out(xor_b[27]) );
  my_xor_155 bc_xor_26 ( .A(B[26]), .B(Cin), .xor_out(xor_b[26]) );
  my_xor_154 bc_xor_25 ( .A(B[25]), .B(Cin), .xor_out(xor_b[25]) );
  my_xor_153 bc_xor_24 ( .A(B[24]), .B(Cin), .xor_out(xor_b[24]) );
  my_xor_152 bc_xor_23 ( .A(B[23]), .B(Cin), .xor_out(xor_b[23]) );
  my_xor_151 bc_xor_22 ( .A(B[22]), .B(Cin), .xor_out(xor_b[22]) );
  my_xor_150 bc_xor_21 ( .A(B[21]), .B(Cin), .xor_out(xor_b[21]) );
  my_xor_149 bc_xor_20 ( .A(B[20]), .B(Cin), .xor_out(xor_b[20]) );
  my_xor_148 bc_xor_19 ( .A(B[19]), .B(Cin), .xor_out(xor_b[19]) );
  my_xor_147 bc_xor_18 ( .A(B[18]), .B(Cin), .xor_out(xor_b[18]) );
  my_xor_146 bc_xor_17 ( .A(B[17]), .B(Cin), .xor_out(xor_b[17]) );
  my_xor_145 bc_xor_16 ( .A(B[16]), .B(Cin), .xor_out(xor_b[16]) );
  my_xor_144 bc_xor_15 ( .A(B[15]), .B(Cin), .xor_out(xor_b[15]) );
  my_xor_143 bc_xor_14 ( .A(B[14]), .B(Cin), .xor_out(xor_b[14]) );
  my_xor_142 bc_xor_13 ( .A(B[13]), .B(Cin), .xor_out(xor_b[13]) );
  my_xor_141 bc_xor_12 ( .A(B[12]), .B(Cin), .xor_out(xor_b[12]) );
  my_xor_140 bc_xor_11 ( .A(B[11]), .B(Cin), .xor_out(xor_b[11]) );
  my_xor_139 bc_xor_10 ( .A(B[10]), .B(Cin), .xor_out(xor_b[10]) );
  my_xor_138 bc_xor_9 ( .A(B[9]), .B(Cin), .xor_out(xor_b[9]) );
  my_xor_137 bc_xor_8 ( .A(B[8]), .B(Cin), .xor_out(xor_b[8]) );
  my_xor_136 bc_xor_7 ( .A(B[7]), .B(Cin), .xor_out(xor_b[7]) );
  my_xor_135 bc_xor_6 ( .A(B[6]), .B(Cin), .xor_out(xor_b[6]) );
  my_xor_134 bc_xor_5 ( .A(B[5]), .B(Cin), .xor_out(xor_b[5]) );
  my_xor_133 bc_xor_4 ( .A(B[4]), .B(Cin), .xor_out(xor_b[4]) );
  my_xor_132 bc_xor_3 ( .A(B[3]), .B(Cin), .xor_out(xor_b[3]) );
  my_xor_131 bc_xor_2 ( .A(B[2]), .B(Cin), .xor_out(xor_b[2]) );
  my_xor_130 bc_xor_1 ( .A(B[1]), .B(Cin), .xor_out(xor_b[1]) );
  my_xor_129 bc_xor_0 ( .A(B[0]), .B(Cin), .xor_out(xor_b[0]) );
  CARRY_GENERATOR_NBIT64_NBIT_PER_BLOCK4_0 CG ( .A(A), .B(xor_b), .Cin(Cin), 
        .Co({Cout, carry}) );
  sum_generator_n_bit64_n_CSB16_0 SG ( .A(A), .B(xor_b), .C_in({carry, Cin}), 
        .S(S) );
  XNOR2_X1 U1 ( .A(A[63]), .B(S[63]), .ZN(n1) );
  NOR2_X1 U2 ( .A1(n1), .A2(n2), .ZN(ovf) );
endmodule


module shl1_NBIT32_1 ( A, Y );
  input [31:0] A;
  output [31:0] Y;
  wire   \A[30] , \A[29] , \A[28] , \A[27] , \A[26] , \A[25] , \A[24] ,
         \A[23] , \A[22] , \A[21] , \A[20] , \A[19] , \A[18] , \A[17] ,
         \A[16] , \A[15] , \A[14] , \A[13] , \A[12] , \A[11] , \A[10] , \A[9] ,
         \A[8] , \A[7] , \A[6] , \A[5] , \A[4] , \A[3] , \A[2] , \A[1] ,
         \A[0] ;
  assign Y[0] = 1'b0;
  assign Y[31] = \A[30] ;
  assign \A[30]  = A[30];
  assign Y[30] = \A[29] ;
  assign \A[29]  = A[29];
  assign Y[29] = \A[28] ;
  assign \A[28]  = A[28];
  assign Y[28] = \A[27] ;
  assign \A[27]  = A[27];
  assign Y[27] = \A[26] ;
  assign \A[26]  = A[26];
  assign Y[26] = \A[25] ;
  assign \A[25]  = A[25];
  assign Y[25] = \A[24] ;
  assign \A[24]  = A[24];
  assign Y[24] = \A[23] ;
  assign \A[23]  = A[23];
  assign Y[23] = \A[22] ;
  assign \A[22]  = A[22];
  assign Y[22] = \A[21] ;
  assign \A[21]  = A[21];
  assign Y[21] = \A[20] ;
  assign \A[20]  = A[20];
  assign Y[20] = \A[19] ;
  assign \A[19]  = A[19];
  assign Y[19] = \A[18] ;
  assign \A[18]  = A[18];
  assign Y[18] = \A[17] ;
  assign \A[17]  = A[17];
  assign Y[17] = \A[16] ;
  assign \A[16]  = A[16];
  assign Y[16] = \A[15] ;
  assign \A[15]  = A[15];
  assign Y[15] = \A[14] ;
  assign \A[14]  = A[14];
  assign Y[14] = \A[13] ;
  assign \A[13]  = A[13];
  assign Y[13] = \A[12] ;
  assign \A[12]  = A[12];
  assign Y[12] = \A[11] ;
  assign \A[11]  = A[11];
  assign Y[11] = \A[10] ;
  assign \A[10]  = A[10];
  assign Y[10] = \A[9] ;
  assign \A[9]  = A[9];
  assign Y[9] = \A[8] ;
  assign \A[8]  = A[8];
  assign Y[8] = \A[7] ;
  assign \A[7]  = A[7];
  assign Y[7] = \A[6] ;
  assign \A[6]  = A[6];
  assign Y[6] = \A[5] ;
  assign \A[5]  = A[5];
  assign Y[5] = \A[4] ;
  assign \A[4]  = A[4];
  assign Y[4] = \A[3] ;
  assign \A[3]  = A[3];
  assign Y[3] = \A[2] ;
  assign \A[2]  = A[2];
  assign Y[2] = \A[1] ;
  assign \A[1]  = A[1];
  assign Y[1] = \A[0] ;
  assign \A[0]  = A[0];

endmodule


module shl2_NBIT32_1 ( A, Y );
  input [31:0] A;
  output [31:0] Y;
  wire   \A[29] , \A[28] , \A[27] , \A[26] , \A[25] , \A[24] , \A[23] ,
         \A[22] , \A[21] , \A[20] , \A[19] , \A[18] , \A[17] , \A[16] ,
         \A[15] , \A[14] , \A[13] , \A[12] , \A[11] , \A[10] , \A[9] , \A[8] ,
         \A[7] , \A[6] , \A[5] , \A[4] , \A[3] , \A[2] , \A[1] , \A[0] ;
  assign Y[0] = 1'b0;
  assign Y[1] = 1'b0;
  assign Y[31] = \A[29] ;
  assign \A[29]  = A[29];
  assign Y[30] = \A[28] ;
  assign \A[28]  = A[28];
  assign Y[29] = \A[27] ;
  assign \A[27]  = A[27];
  assign Y[28] = \A[26] ;
  assign \A[26]  = A[26];
  assign Y[27] = \A[25] ;
  assign \A[25]  = A[25];
  assign Y[26] = \A[24] ;
  assign \A[24]  = A[24];
  assign Y[25] = \A[23] ;
  assign \A[23]  = A[23];
  assign Y[24] = \A[22] ;
  assign \A[22]  = A[22];
  assign Y[23] = \A[21] ;
  assign \A[21]  = A[21];
  assign Y[22] = \A[20] ;
  assign \A[20]  = A[20];
  assign Y[21] = \A[19] ;
  assign \A[19]  = A[19];
  assign Y[20] = \A[18] ;
  assign \A[18]  = A[18];
  assign Y[19] = \A[17] ;
  assign \A[17]  = A[17];
  assign Y[18] = \A[16] ;
  assign \A[16]  = A[16];
  assign Y[17] = \A[15] ;
  assign \A[15]  = A[15];
  assign Y[16] = \A[14] ;
  assign \A[14]  = A[14];
  assign Y[15] = \A[13] ;
  assign \A[13]  = A[13];
  assign Y[14] = \A[12] ;
  assign \A[12]  = A[12];
  assign Y[13] = \A[11] ;
  assign \A[11]  = A[11];
  assign Y[12] = \A[10] ;
  assign \A[10]  = A[10];
  assign Y[11] = \A[9] ;
  assign \A[9]  = A[9];
  assign Y[10] = \A[8] ;
  assign \A[8]  = A[8];
  assign Y[9] = \A[7] ;
  assign \A[7]  = A[7];
  assign Y[8] = \A[6] ;
  assign \A[6]  = A[6];
  assign Y[7] = \A[5] ;
  assign \A[5]  = A[5];
  assign Y[6] = \A[4] ;
  assign \A[4]  = A[4];
  assign Y[5] = \A[3] ;
  assign \A[3]  = A[3];
  assign Y[4] = \A[2] ;
  assign \A[2]  = A[2];
  assign Y[3] = \A[1] ;
  assign \A[1]  = A[1];
  assign Y[2] = \A[0] ;
  assign \A[0]  = A[0];

endmodule


module negate_NBIT32_2_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n56,
         n57, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U1 ( .A(n88), .B(n4), .Z(DIFF[5]) );
  XOR2_X1 U2 ( .A(n89), .B(n3), .Z(DIFF[4]) );
  AND2_X1 U3 ( .A1(n90), .A2(n56), .ZN(n3) );
  AND2_X1 U4 ( .A1(n89), .A2(n3), .ZN(n4) );
  AND2_X1 U5 ( .A1(n88), .A2(n4), .ZN(n5) );
  AND2_X1 U6 ( .A1(n87), .A2(n5), .ZN(n6) );
  AND2_X1 U7 ( .A1(n86), .A2(n6), .ZN(n7) );
  AND2_X1 U8 ( .A1(n85), .A2(n7), .ZN(n8) );
  AND2_X1 U9 ( .A1(n84), .A2(n8), .ZN(n9) );
  AND2_X1 U10 ( .A1(n83), .A2(n9), .ZN(n10) );
  AND2_X1 U11 ( .A1(n82), .A2(n10), .ZN(n11) );
  AND2_X1 U12 ( .A1(n81), .A2(n11), .ZN(n12) );
  AND2_X1 U13 ( .A1(n80), .A2(n12), .ZN(n13) );
  AND2_X1 U14 ( .A1(n79), .A2(n13), .ZN(n14) );
  AND2_X1 U15 ( .A1(n78), .A2(n14), .ZN(n15) );
  AND2_X1 U16 ( .A1(n77), .A2(n15), .ZN(n16) );
  AND2_X1 U17 ( .A1(n76), .A2(n16), .ZN(n17) );
  AND2_X1 U18 ( .A1(n75), .A2(n17), .ZN(n18) );
  AND2_X1 U19 ( .A1(n74), .A2(n18), .ZN(n19) );
  AND2_X1 U20 ( .A1(n73), .A2(n19), .ZN(n20) );
  AND2_X1 U21 ( .A1(n72), .A2(n20), .ZN(n21) );
  AND2_X1 U22 ( .A1(n71), .A2(n21), .ZN(n22) );
  AND2_X1 U23 ( .A1(n70), .A2(n22), .ZN(n23) );
  AND2_X1 U24 ( .A1(n69), .A2(n23), .ZN(n24) );
  AND2_X1 U25 ( .A1(n68), .A2(n24), .ZN(n25) );
  AND2_X1 U26 ( .A1(n67), .A2(n25), .ZN(n26) );
  AND2_X1 U27 ( .A1(n66), .A2(n26), .ZN(n27) );
  AND2_X1 U28 ( .A1(n65), .A2(n27), .ZN(n28) );
  AND2_X1 U29 ( .A1(n64), .A2(n28), .ZN(n29) );
  NAND2_X1 U30 ( .A1(n63), .A2(n29), .ZN(n61) );
  XOR2_X1 U31 ( .A(n63), .B(n29), .Z(DIFF[30]) );
  XOR2_X1 U32 ( .A(n64), .B(n28), .Z(DIFF[29]) );
  XOR2_X1 U33 ( .A(n65), .B(n27), .Z(DIFF[28]) );
  XOR2_X1 U34 ( .A(n66), .B(n26), .Z(DIFF[27]) );
  XOR2_X1 U35 ( .A(n67), .B(n25), .Z(DIFF[26]) );
  XOR2_X1 U36 ( .A(n68), .B(n24), .Z(DIFF[25]) );
  XOR2_X1 U37 ( .A(n69), .B(n23), .Z(DIFF[24]) );
  XOR2_X1 U38 ( .A(n70), .B(n22), .Z(DIFF[23]) );
  XOR2_X1 U39 ( .A(n71), .B(n21), .Z(DIFF[22]) );
  XOR2_X1 U40 ( .A(n72), .B(n20), .Z(DIFF[21]) );
  XOR2_X1 U41 ( .A(n73), .B(n19), .Z(DIFF[20]) );
  XOR2_X1 U42 ( .A(n74), .B(n18), .Z(DIFF[19]) );
  XOR2_X1 U43 ( .A(n75), .B(n17), .Z(DIFF[18]) );
  XOR2_X1 U44 ( .A(n76), .B(n16), .Z(DIFF[17]) );
  XOR2_X1 U45 ( .A(n77), .B(n15), .Z(DIFF[16]) );
  XOR2_X1 U46 ( .A(n78), .B(n14), .Z(DIFF[15]) );
  XOR2_X1 U47 ( .A(n79), .B(n13), .Z(DIFF[14]) );
  XOR2_X1 U48 ( .A(n80), .B(n12), .Z(DIFF[13]) );
  XOR2_X1 U49 ( .A(n81), .B(n11), .Z(DIFF[12]) );
  XOR2_X1 U50 ( .A(n82), .B(n10), .Z(DIFF[11]) );
  XOR2_X1 U51 ( .A(n83), .B(n9), .Z(DIFF[10]) );
  XOR2_X1 U52 ( .A(n84), .B(n8), .Z(DIFF[9]) );
  XOR2_X1 U53 ( .A(n85), .B(n7), .Z(DIFF[8]) );
  XOR2_X1 U54 ( .A(n86), .B(n6), .Z(DIFF[7]) );
  XOR2_X1 U55 ( .A(n87), .B(n5), .Z(DIFF[6]) );
  XOR2_X1 U56 ( .A(n90), .B(n56), .Z(DIFF[3]) );
  AND2_X1 U57 ( .A1(n91), .A2(n57), .ZN(n56) );
  AND2_X1 U58 ( .A1(n92), .A2(n62), .ZN(n57) );
  XOR2_X1 U59 ( .A(n91), .B(n57), .Z(DIFF[2]) );
  XOR2_X1 U60 ( .A(n92), .B(n62), .Z(DIFF[1]) );
  INV_X1 U61 ( .A(B[3]), .ZN(n90) );
  INV_X1 U62 ( .A(B[4]), .ZN(n89) );
  INV_X1 U63 ( .A(B[5]), .ZN(n88) );
  INV_X1 U64 ( .A(B[6]), .ZN(n87) );
  INV_X1 U65 ( .A(B[7]), .ZN(n86) );
  INV_X1 U66 ( .A(B[8]), .ZN(n85) );
  INV_X1 U67 ( .A(B[9]), .ZN(n84) );
  INV_X1 U68 ( .A(B[10]), .ZN(n83) );
  INV_X1 U69 ( .A(B[11]), .ZN(n82) );
  INV_X1 U70 ( .A(B[12]), .ZN(n81) );
  INV_X1 U71 ( .A(B[13]), .ZN(n80) );
  XOR2_X1 U72 ( .A(B[31]), .B(n61), .Z(DIFF[31]) );
  INV_X1 U73 ( .A(B[14]), .ZN(n79) );
  INV_X1 U74 ( .A(B[15]), .ZN(n78) );
  INV_X1 U75 ( .A(B[16]), .ZN(n77) );
  INV_X1 U76 ( .A(B[17]), .ZN(n76) );
  INV_X1 U77 ( .A(B[18]), .ZN(n75) );
  INV_X1 U78 ( .A(B[19]), .ZN(n74) );
  INV_X1 U79 ( .A(B[20]), .ZN(n73) );
  INV_X1 U80 ( .A(B[21]), .ZN(n72) );
  INV_X1 U81 ( .A(B[22]), .ZN(n71) );
  INV_X1 U82 ( .A(B[23]), .ZN(n70) );
  INV_X1 U83 ( .A(B[24]), .ZN(n69) );
  INV_X1 U84 ( .A(B[25]), .ZN(n68) );
  INV_X1 U85 ( .A(B[26]), .ZN(n67) );
  INV_X1 U86 ( .A(B[27]), .ZN(n66) );
  INV_X1 U87 ( .A(B[28]), .ZN(n65) );
  INV_X1 U88 ( .A(B[29]), .ZN(n64) );
  INV_X1 U89 ( .A(B[30]), .ZN(n63) );
  INV_X1 U90 ( .A(\B[0] ), .ZN(n62) );
  INV_X1 U91 ( .A(B[1]), .ZN(n92) );
  INV_X1 U92 ( .A(B[2]), .ZN(n91) );
endmodule


module negate_NBIT32_2 ( A, Y );
  input [31:0] A;
  output [31:0] Y;


  negate_NBIT32_2_DW01_sub_0 sub_add_14_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .B(A), .CI(1'b0), .DIFF(Y) );
endmodule


module negate_NBIT32_1_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  XOR2_X1 U1 ( .A(B[31]), .B(n61), .Z(DIFF[31]) );
  XOR2_X1 U2 ( .A(n64), .B(n55), .Z(DIFF[30]) );
  XOR2_X1 U3 ( .A(n65), .B(n54), .Z(DIFF[29]) );
  XOR2_X1 U4 ( .A(n66), .B(n53), .Z(DIFF[28]) );
  XOR2_X1 U5 ( .A(n67), .B(n52), .Z(DIFF[27]) );
  XOR2_X1 U6 ( .A(n68), .B(n51), .Z(DIFF[26]) );
  XOR2_X1 U7 ( .A(n69), .B(n50), .Z(DIFF[25]) );
  XOR2_X1 U8 ( .A(n70), .B(n49), .Z(DIFF[24]) );
  XOR2_X1 U9 ( .A(n71), .B(n48), .Z(DIFF[23]) );
  XOR2_X1 U10 ( .A(n72), .B(n47), .Z(DIFF[22]) );
  XOR2_X1 U11 ( .A(n73), .B(n46), .Z(DIFF[21]) );
  XOR2_X1 U12 ( .A(n74), .B(n45), .Z(DIFF[20]) );
  XOR2_X1 U13 ( .A(n75), .B(n44), .Z(DIFF[19]) );
  XOR2_X1 U14 ( .A(n76), .B(n43), .Z(DIFF[18]) );
  XOR2_X1 U15 ( .A(n77), .B(n42), .Z(DIFF[17]) );
  XOR2_X1 U16 ( .A(n78), .B(n41), .Z(DIFF[16]) );
  XOR2_X1 U17 ( .A(n79), .B(n40), .Z(DIFF[15]) );
  XOR2_X1 U18 ( .A(n80), .B(n39), .Z(DIFF[14]) );
  XOR2_X1 U19 ( .A(n81), .B(n38), .Z(DIFF[13]) );
  XOR2_X1 U20 ( .A(n82), .B(n37), .Z(DIFF[12]) );
  XOR2_X1 U21 ( .A(n83), .B(n36), .Z(DIFF[11]) );
  XOR2_X1 U22 ( .A(n84), .B(n35), .Z(DIFF[10]) );
  XOR2_X1 U23 ( .A(n85), .B(n34), .Z(DIFF[9]) );
  XOR2_X1 U24 ( .A(n86), .B(n33), .Z(DIFF[8]) );
  XOR2_X1 U25 ( .A(n87), .B(n32), .Z(DIFF[7]) );
  XOR2_X1 U26 ( .A(n88), .B(n31), .Z(DIFF[6]) );
  XOR2_X1 U27 ( .A(n91), .B(n59), .Z(DIFF[3]) );
  XOR2_X1 U28 ( .A(n92), .B(n60), .Z(DIFF[2]) );
  XOR2_X1 U29 ( .A(n63), .B(n62), .Z(DIFF[1]) );
  AND2_X1 U30 ( .A1(n90), .A2(n58), .ZN(n30) );
  AND2_X1 U31 ( .A1(n89), .A2(n30), .ZN(n31) );
  AND2_X1 U32 ( .A1(n88), .A2(n31), .ZN(n32) );
  AND2_X1 U33 ( .A1(n87), .A2(n32), .ZN(n33) );
  AND2_X1 U34 ( .A1(n86), .A2(n33), .ZN(n34) );
  AND2_X1 U35 ( .A1(n85), .A2(n34), .ZN(n35) );
  AND2_X1 U36 ( .A1(n84), .A2(n35), .ZN(n36) );
  AND2_X1 U37 ( .A1(n83), .A2(n36), .ZN(n37) );
  AND2_X1 U38 ( .A1(n82), .A2(n37), .ZN(n38) );
  AND2_X1 U39 ( .A1(n81), .A2(n38), .ZN(n39) );
  AND2_X1 U40 ( .A1(n80), .A2(n39), .ZN(n40) );
  AND2_X1 U41 ( .A1(n79), .A2(n40), .ZN(n41) );
  AND2_X1 U42 ( .A1(n78), .A2(n41), .ZN(n42) );
  AND2_X1 U43 ( .A1(n77), .A2(n42), .ZN(n43) );
  AND2_X1 U44 ( .A1(n76), .A2(n43), .ZN(n44) );
  AND2_X1 U45 ( .A1(n75), .A2(n44), .ZN(n45) );
  AND2_X1 U46 ( .A1(n74), .A2(n45), .ZN(n46) );
  AND2_X1 U47 ( .A1(n73), .A2(n46), .ZN(n47) );
  AND2_X1 U48 ( .A1(n72), .A2(n47), .ZN(n48) );
  AND2_X1 U49 ( .A1(n71), .A2(n48), .ZN(n49) );
  AND2_X1 U50 ( .A1(n70), .A2(n49), .ZN(n50) );
  AND2_X1 U51 ( .A1(n69), .A2(n50), .ZN(n51) );
  AND2_X1 U52 ( .A1(n68), .A2(n51), .ZN(n52) );
  AND2_X1 U53 ( .A1(n67), .A2(n52), .ZN(n53) );
  AND2_X1 U54 ( .A1(n66), .A2(n53), .ZN(n54) );
  AND2_X1 U55 ( .A1(n65), .A2(n54), .ZN(n55) );
  XOR2_X1 U56 ( .A(n89), .B(n30), .Z(DIFF[5]) );
  XOR2_X1 U57 ( .A(n90), .B(n58), .Z(DIFF[4]) );
  AND2_X1 U58 ( .A1(n91), .A2(n59), .ZN(n58) );
  AND2_X1 U59 ( .A1(n92), .A2(n60), .ZN(n59) );
  AND2_X1 U60 ( .A1(n63), .A2(n62), .ZN(n60) );
  NAND2_X1 U61 ( .A1(n64), .A2(n55), .ZN(n61) );
  INV_X1 U62 ( .A(B[4]), .ZN(n90) );
  INV_X1 U63 ( .A(B[5]), .ZN(n89) );
  INV_X1 U64 ( .A(B[6]), .ZN(n88) );
  INV_X1 U65 ( .A(B[7]), .ZN(n87) );
  INV_X1 U66 ( .A(B[8]), .ZN(n86) );
  INV_X1 U67 ( .A(B[9]), .ZN(n85) );
  INV_X1 U68 ( .A(B[10]), .ZN(n84) );
  INV_X1 U69 ( .A(B[11]), .ZN(n83) );
  INV_X1 U70 ( .A(B[12]), .ZN(n82) );
  INV_X1 U71 ( .A(B[13]), .ZN(n81) );
  INV_X1 U72 ( .A(B[14]), .ZN(n80) );
  INV_X1 U73 ( .A(B[15]), .ZN(n79) );
  INV_X1 U74 ( .A(B[16]), .ZN(n78) );
  INV_X1 U75 ( .A(B[17]), .ZN(n77) );
  INV_X1 U76 ( .A(B[18]), .ZN(n76) );
  INV_X1 U77 ( .A(B[19]), .ZN(n75) );
  INV_X1 U78 ( .A(B[20]), .ZN(n74) );
  INV_X1 U79 ( .A(B[21]), .ZN(n73) );
  INV_X1 U80 ( .A(B[22]), .ZN(n72) );
  INV_X1 U81 ( .A(B[23]), .ZN(n71) );
  INV_X1 U82 ( .A(B[24]), .ZN(n70) );
  INV_X1 U83 ( .A(B[25]), .ZN(n69) );
  INV_X1 U84 ( .A(B[26]), .ZN(n68) );
  INV_X1 U85 ( .A(B[27]), .ZN(n67) );
  INV_X1 U86 ( .A(B[28]), .ZN(n66) );
  INV_X1 U87 ( .A(B[29]), .ZN(n65) );
  INV_X1 U88 ( .A(B[30]), .ZN(n64) );
  INV_X1 U89 ( .A(\B[0] ), .ZN(n62) );
  INV_X1 U90 ( .A(B[1]), .ZN(n63) );
  INV_X1 U91 ( .A(B[2]), .ZN(n92) );
  INV_X1 U92 ( .A(B[3]), .ZN(n91) );
endmodule


module negate_NBIT32_1 ( A, Y );
  input [31:0] A;
  output [31:0] Y;


  negate_NBIT32_1_DW01_sub_0 sub_add_14_b0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .B(A), .CI(1'b0), .DIFF(Y) );
endmodule


module mux51_gen_NBIT32_1 ( A0, A1, A2, A3, A4, SEL, Y );
  input [31:0] A0;
  input [31:0] A1;
  input [31:0] A2;
  input [31:0] A3;
  input [31:0] A4;
  input [2:0] SEL;
  output [31:0] Y;
  wire   n1, n2, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155;

  BUF_X1 U2 ( .A(n150), .Z(n74) );
  BUF_X1 U3 ( .A(n150), .Z(n73) );
  BUF_X1 U4 ( .A(n149), .Z(n1) );
  BUF_X1 U5 ( .A(n153), .Z(n83) );
  BUF_X1 U6 ( .A(n153), .Z(n82) );
  BUF_X1 U7 ( .A(n153), .Z(n84) );
  BUF_X1 U8 ( .A(n152), .Z(n80) );
  BUF_X1 U9 ( .A(n152), .Z(n79) );
  BUF_X1 U10 ( .A(n151), .Z(n77) );
  BUF_X1 U11 ( .A(n151), .Z(n76) );
  BUF_X1 U12 ( .A(n150), .Z(n75) );
  BUF_X1 U13 ( .A(n152), .Z(n81) );
  BUF_X1 U14 ( .A(n151), .Z(n78) );
  BUF_X1 U15 ( .A(n149), .Z(n2) );
  BUF_X1 U16 ( .A(n149), .Z(n72) );
  NAND2_X1 U17 ( .A1(n134), .A2(n133), .ZN(Y[30]) );
  AOI22_X1 U18 ( .A1(A4[30]), .A2(n74), .B1(A0[30]), .B2(n72), .ZN(n134) );
  AOI222_X1 U19 ( .A1(A2[30]), .A2(n84), .B1(A1[30]), .B2(n80), .C1(A3[30]), 
        .C2(n77), .ZN(n133) );
  NAND2_X1 U20 ( .A1(n130), .A2(n129), .ZN(Y[29]) );
  AOI22_X1 U21 ( .A1(A4[29]), .A2(n74), .B1(A0[29]), .B2(n2), .ZN(n130) );
  AOI222_X1 U22 ( .A1(A2[29]), .A2(n83), .B1(A1[29]), .B2(n80), .C1(A3[29]), 
        .C2(n77), .ZN(n129) );
  NAND2_X1 U23 ( .A1(n128), .A2(n127), .ZN(Y[28]) );
  AOI22_X1 U24 ( .A1(A4[28]), .A2(n74), .B1(A0[28]), .B2(n2), .ZN(n128) );
  AOI222_X1 U25 ( .A1(A2[28]), .A2(n83), .B1(A1[28]), .B2(n80), .C1(A3[28]), 
        .C2(n77), .ZN(n127) );
  NAND2_X1 U26 ( .A1(n126), .A2(n125), .ZN(Y[27]) );
  AOI22_X1 U27 ( .A1(A4[27]), .A2(n74), .B1(A0[27]), .B2(n2), .ZN(n126) );
  AOI222_X1 U28 ( .A1(A2[27]), .A2(n83), .B1(A1[27]), .B2(n80), .C1(A3[27]), 
        .C2(n77), .ZN(n125) );
  NAND2_X1 U29 ( .A1(n124), .A2(n123), .ZN(Y[26]) );
  AOI22_X1 U30 ( .A1(A4[26]), .A2(n74), .B1(A0[26]), .B2(n2), .ZN(n124) );
  AOI222_X1 U31 ( .A1(A2[26]), .A2(n83), .B1(A1[26]), .B2(n80), .C1(A3[26]), 
        .C2(n77), .ZN(n123) );
  NAND2_X1 U32 ( .A1(n122), .A2(n121), .ZN(Y[25]) );
  AOI22_X1 U33 ( .A1(A4[25]), .A2(n74), .B1(A0[25]), .B2(n2), .ZN(n122) );
  AOI222_X1 U34 ( .A1(A2[25]), .A2(n83), .B1(A1[25]), .B2(n80), .C1(A3[25]), 
        .C2(n77), .ZN(n121) );
  NAND2_X1 U35 ( .A1(n120), .A2(n119), .ZN(Y[24]) );
  AOI22_X1 U36 ( .A1(A4[24]), .A2(n74), .B1(A0[24]), .B2(n2), .ZN(n120) );
  AOI222_X1 U37 ( .A1(A2[24]), .A2(n83), .B1(A1[24]), .B2(n80), .C1(A3[24]), 
        .C2(n77), .ZN(n119) );
  NAND2_X1 U38 ( .A1(n118), .A2(n117), .ZN(Y[23]) );
  AOI22_X1 U39 ( .A1(A4[23]), .A2(n74), .B1(A0[23]), .B2(n2), .ZN(n118) );
  AOI222_X1 U40 ( .A1(A2[23]), .A2(n83), .B1(A1[23]), .B2(n80), .C1(A3[23]), 
        .C2(n77), .ZN(n117) );
  NAND2_X1 U41 ( .A1(n116), .A2(n115), .ZN(Y[22]) );
  AOI22_X1 U42 ( .A1(A4[22]), .A2(n74), .B1(A0[22]), .B2(n2), .ZN(n116) );
  AOI222_X1 U43 ( .A1(A2[22]), .A2(n83), .B1(A1[22]), .B2(n80), .C1(A3[22]), 
        .C2(n77), .ZN(n115) );
  NAND2_X1 U44 ( .A1(n114), .A2(n113), .ZN(Y[21]) );
  AOI22_X1 U45 ( .A1(A4[21]), .A2(n74), .B1(A0[21]), .B2(n2), .ZN(n114) );
  AOI222_X1 U46 ( .A1(A2[21]), .A2(n83), .B1(A1[21]), .B2(n80), .C1(A3[21]), 
        .C2(n77), .ZN(n113) );
  NAND2_X1 U47 ( .A1(n136), .A2(n135), .ZN(Y[31]) );
  AOI22_X1 U48 ( .A1(A4[31]), .A2(n75), .B1(A0[31]), .B2(n72), .ZN(n136) );
  AOI222_X1 U49 ( .A1(A2[31]), .A2(n84), .B1(A1[31]), .B2(n81), .C1(A3[31]), 
        .C2(n78), .ZN(n135) );
  NAND2_X1 U50 ( .A1(n112), .A2(n111), .ZN(Y[20]) );
  AOI22_X1 U51 ( .A1(A4[20]), .A2(n74), .B1(A0[20]), .B2(n2), .ZN(n112) );
  AOI222_X1 U52 ( .A1(A2[20]), .A2(n83), .B1(A1[20]), .B2(n80), .C1(A3[20]), 
        .C2(n77), .ZN(n111) );
  NAND2_X1 U53 ( .A1(n108), .A2(n107), .ZN(Y[19]) );
  AOI22_X1 U54 ( .A1(A4[19]), .A2(n73), .B1(A0[19]), .B2(n1), .ZN(n108) );
  AOI222_X1 U55 ( .A1(A2[19]), .A2(n82), .B1(A1[19]), .B2(n79), .C1(A3[19]), 
        .C2(n76), .ZN(n107) );
  NAND2_X1 U56 ( .A1(n106), .A2(n105), .ZN(Y[18]) );
  AOI22_X1 U57 ( .A1(A4[18]), .A2(n73), .B1(A0[18]), .B2(n1), .ZN(n106) );
  AOI222_X1 U58 ( .A1(A2[18]), .A2(n82), .B1(A1[18]), .B2(n79), .C1(A3[18]), 
        .C2(n76), .ZN(n105) );
  NAND2_X1 U59 ( .A1(n104), .A2(n103), .ZN(Y[17]) );
  AOI22_X1 U60 ( .A1(A4[17]), .A2(n73), .B1(A0[17]), .B2(n1), .ZN(n104) );
  AOI222_X1 U61 ( .A1(A2[17]), .A2(n82), .B1(A1[17]), .B2(n79), .C1(A3[17]), 
        .C2(n76), .ZN(n103) );
  NAND2_X1 U62 ( .A1(n102), .A2(n101), .ZN(Y[16]) );
  AOI22_X1 U63 ( .A1(A4[16]), .A2(n73), .B1(A0[16]), .B2(n1), .ZN(n102) );
  AOI222_X1 U64 ( .A1(A2[16]), .A2(n82), .B1(A1[16]), .B2(n79), .C1(A3[16]), 
        .C2(n76), .ZN(n101) );
  NAND2_X1 U65 ( .A1(n100), .A2(n99), .ZN(Y[15]) );
  AOI22_X1 U66 ( .A1(A4[15]), .A2(n73), .B1(A0[15]), .B2(n1), .ZN(n100) );
  AOI222_X1 U67 ( .A1(A2[15]), .A2(n82), .B1(A1[15]), .B2(n79), .C1(A3[15]), 
        .C2(n76), .ZN(n99) );
  NAND2_X1 U68 ( .A1(n98), .A2(n97), .ZN(Y[14]) );
  AOI22_X1 U69 ( .A1(A4[14]), .A2(n73), .B1(A0[14]), .B2(n1), .ZN(n98) );
  AOI222_X1 U70 ( .A1(A2[14]), .A2(n82), .B1(A1[14]), .B2(n79), .C1(A3[14]), 
        .C2(n76), .ZN(n97) );
  NAND2_X1 U71 ( .A1(n96), .A2(n95), .ZN(Y[13]) );
  AOI22_X1 U72 ( .A1(A4[13]), .A2(n73), .B1(A0[13]), .B2(n1), .ZN(n96) );
  AOI222_X1 U73 ( .A1(A2[13]), .A2(n82), .B1(A1[13]), .B2(n79), .C1(A3[13]), 
        .C2(n76), .ZN(n95) );
  NAND2_X1 U74 ( .A1(n94), .A2(n93), .ZN(Y[12]) );
  AOI22_X1 U75 ( .A1(A4[12]), .A2(n73), .B1(A0[12]), .B2(n1), .ZN(n94) );
  AOI222_X1 U76 ( .A1(A2[12]), .A2(n82), .B1(A1[12]), .B2(n79), .C1(A3[12]), 
        .C2(n76), .ZN(n93) );
  NAND2_X1 U77 ( .A1(n92), .A2(n91), .ZN(Y[11]) );
  AOI22_X1 U78 ( .A1(A4[11]), .A2(n73), .B1(A0[11]), .B2(n1), .ZN(n92) );
  AOI222_X1 U79 ( .A1(A2[11]), .A2(n82), .B1(A1[11]), .B2(n79), .C1(A3[11]), 
        .C2(n76), .ZN(n91) );
  NAND2_X1 U80 ( .A1(n90), .A2(n89), .ZN(Y[10]) );
  AOI22_X1 U81 ( .A1(A4[10]), .A2(n73), .B1(A0[10]), .B2(n1), .ZN(n90) );
  AOI222_X1 U82 ( .A1(A2[10]), .A2(n82), .B1(A1[10]), .B2(n79), .C1(A3[10]), 
        .C2(n76), .ZN(n89) );
  NAND2_X1 U83 ( .A1(n155), .A2(n154), .ZN(Y[9]) );
  AOI22_X1 U84 ( .A1(A4[9]), .A2(n75), .B1(A0[9]), .B2(n72), .ZN(n155) );
  AOI222_X1 U85 ( .A1(A2[9]), .A2(n84), .B1(A1[9]), .B2(n81), .C1(A3[9]), .C2(
        n78), .ZN(n154) );
  NAND2_X1 U86 ( .A1(n148), .A2(n147), .ZN(Y[8]) );
  AOI22_X1 U87 ( .A1(A4[8]), .A2(n75), .B1(A0[8]), .B2(n72), .ZN(n148) );
  AOI222_X1 U88 ( .A1(A2[8]), .A2(n84), .B1(A1[8]), .B2(n81), .C1(A3[8]), .C2(
        n78), .ZN(n147) );
  NAND2_X1 U89 ( .A1(n146), .A2(n145), .ZN(Y[7]) );
  AOI22_X1 U90 ( .A1(A4[7]), .A2(n75), .B1(A0[7]), .B2(n72), .ZN(n146) );
  AOI222_X1 U91 ( .A1(A2[7]), .A2(n84), .B1(A1[7]), .B2(n81), .C1(A3[7]), .C2(
        n78), .ZN(n145) );
  NAND2_X1 U92 ( .A1(n138), .A2(n137), .ZN(Y[3]) );
  AOI22_X1 U93 ( .A1(A4[3]), .A2(n75), .B1(A0[3]), .B2(n72), .ZN(n138) );
  AOI222_X1 U94 ( .A1(A2[3]), .A2(n84), .B1(A1[3]), .B2(n81), .C1(A3[3]), .C2(
        n78), .ZN(n137) );
  NOR3_X1 U95 ( .A1(SEL[0]), .A2(SEL[1]), .A3(n1), .ZN(n150) );
  NOR3_X1 U96 ( .A1(SEL[1]), .A2(SEL[2]), .A3(SEL[0]), .ZN(n149) );
  NOR3_X1 U97 ( .A1(SEL[0]), .A2(SEL[2]), .A3(n86), .ZN(n153) );
  NAND2_X1 U98 ( .A1(n142), .A2(n141), .ZN(Y[5]) );
  AOI222_X1 U99 ( .A1(A2[5]), .A2(n84), .B1(A1[5]), .B2(n81), .C1(A3[5]), .C2(
        n78), .ZN(n141) );
  AOI22_X1 U100 ( .A1(A4[5]), .A2(n75), .B1(A0[5]), .B2(n72), .ZN(n142) );
  NAND2_X1 U101 ( .A1(n140), .A2(n139), .ZN(Y[4]) );
  AOI222_X1 U102 ( .A1(A2[4]), .A2(n84), .B1(A1[4]), .B2(n81), .C1(A3[4]), 
        .C2(n78), .ZN(n139) );
  AOI22_X1 U103 ( .A1(A4[4]), .A2(n75), .B1(A0[4]), .B2(n72), .ZN(n140) );
  AND3_X1 U104 ( .A1(SEL[0]), .A2(n85), .A3(SEL[1]), .ZN(n151) );
  AND3_X1 U105 ( .A1(n86), .A2(n85), .A3(SEL[0]), .ZN(n152) );
  INV_X1 U106 ( .A(SEL[1]), .ZN(n86) );
  NAND2_X1 U107 ( .A1(n144), .A2(n143), .ZN(Y[6]) );
  AOI22_X1 U108 ( .A1(A4[6]), .A2(n75), .B1(A0[6]), .B2(n72), .ZN(n144) );
  AOI222_X1 U109 ( .A1(A2[6]), .A2(n84), .B1(A1[6]), .B2(n81), .C1(A3[6]), 
        .C2(n78), .ZN(n143) );
  INV_X1 U110 ( .A(SEL[2]), .ZN(n85) );
  NAND2_X1 U111 ( .A1(n110), .A2(n109), .ZN(Y[1]) );
  AOI22_X1 U112 ( .A1(A4[1]), .A2(n73), .B1(A0[1]), .B2(n2), .ZN(n110) );
  AOI222_X1 U113 ( .A1(A2[1]), .A2(n83), .B1(A1[1]), .B2(n79), .C1(A3[1]), 
        .C2(n76), .ZN(n109) );
  NAND2_X1 U114 ( .A1(n132), .A2(n131), .ZN(Y[2]) );
  AOI22_X1 U115 ( .A1(A4[2]), .A2(n74), .B1(A0[2]), .B2(n2), .ZN(n132) );
  AOI222_X1 U116 ( .A1(A2[2]), .A2(n84), .B1(A1[2]), .B2(n80), .C1(A3[2]), 
        .C2(n77), .ZN(n131) );
  NAND2_X1 U117 ( .A1(n88), .A2(n87), .ZN(Y[0]) );
  AOI22_X1 U118 ( .A1(A4[0]), .A2(n73), .B1(A0[0]), .B2(n1), .ZN(n88) );
  AOI222_X1 U119 ( .A1(A2[0]), .A2(n82), .B1(A1[0]), .B2(n79), .C1(A3[0]), 
        .C2(n76), .ZN(n87) );
endmodule


module my_xor_128 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_127 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_126 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_125 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_124 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_123 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_122 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_121 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_120 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_119 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_118 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_117 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_116 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_115 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_114 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_113 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_112 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_111 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_110 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_109 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_108 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_107 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_106 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_105 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_104 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_103 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_102 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_101 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_100 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_99 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_98 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_97 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_96 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_95 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_94 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_93 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_92 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_91 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_90 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_89 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_88 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_87 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_86 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_85 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_84 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_83 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_82 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_81 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_80 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_79 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_78 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_77 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_76 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_75 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_74 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_73 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_72 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_71 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_70 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_69 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_68 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_67 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_66 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_65 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module pg_net_126 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_125 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_124 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_123 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_122 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_121 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_120 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_119 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_118 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_117 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_116 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_115 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_114 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_113 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_112 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_111 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_110 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_109 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_108 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_107 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_106 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_105 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_104 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_103 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_102 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_101 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_100 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_99 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_98 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_97 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_96 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_95 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_94 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_93 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_92 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_91 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_90 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_89 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_88 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_87 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_86 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_85 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_84 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_83 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_82 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_81 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_80 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_79 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_78 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_77 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_76 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_75 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_74 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_73 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_72 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_71 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_70 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_69 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_68 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_67 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_66 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_65 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_64 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_BLOCK_126 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_125 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_124 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_123 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_122 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_121 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_120 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_119 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_118 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_117 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_116 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_115 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_114 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_113 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_112 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_111 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_110 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_109 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_108 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_107 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_106 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_105 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_104 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_103 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_102 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_101 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_100 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_99 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_98 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_97 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_96 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_34 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_95 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_94 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_93 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_92 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_91 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_90 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_89 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_88 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_87 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AOI21_X1 U1 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_86 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_85 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_84 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_83 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_82 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_81 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_33 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_80 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_79 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_78 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_77 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_76 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_75 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_74 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_32 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_73 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_72 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_71 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_70 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_69 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_68 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_31 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_30 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_67 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AND2_X1 U2 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_66 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_65 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_64 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_29 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_28 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_27 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_26 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_25 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_24 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_23 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_22 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_21 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_20 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_19 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_18 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module CARRY_GENERATOR_NBIT64_NBIT_PER_BLOCK4_2 ( A, B, Cin, Co );
  input [63:0] A;
  input [63:0] B;
  output [15:0] Co;
  input Cin;
  wire   \g_vector[5][63] , \g_vector[5][59] , \g_vector[5][55] ,
         \g_vector[5][51] , \g_vector[4][63] , \g_vector[4][59] ,
         \g_vector[4][47] , \g_vector[4][43] , \g_vector[4][31] ,
         \g_vector[4][27] , \g_vector[3][63] , \g_vector[3][55] ,
         \g_vector[3][47] , \g_vector[3][39] , \g_vector[3][31] ,
         \g_vector[3][23] , \g_vector[3][15] , \g_vector[2][63] ,
         \g_vector[2][59] , \g_vector[2][55] , \g_vector[2][51] ,
         \g_vector[2][47] , \g_vector[2][43] , \g_vector[2][39] ,
         \g_vector[2][35] , \g_vector[2][31] , \g_vector[2][27] ,
         \g_vector[2][23] , \g_vector[2][19] , \g_vector[2][15] ,
         \g_vector[2][11] , \g_vector[2][7] , \g_vector[1][63] ,
         \g_vector[1][61] , \g_vector[1][59] , \g_vector[1][57] ,
         \g_vector[1][55] , \g_vector[1][53] , \g_vector[1][51] ,
         \g_vector[1][49] , \g_vector[1][47] , \g_vector[1][45] ,
         \g_vector[1][43] , \g_vector[1][41] , \g_vector[1][39] ,
         \g_vector[1][37] , \g_vector[1][35] , \g_vector[1][33] ,
         \g_vector[1][31] , \g_vector[1][29] , \g_vector[1][27] ,
         \g_vector[1][25] , \g_vector[1][23] , \g_vector[1][21] ,
         \g_vector[1][19] , \g_vector[1][17] , \g_vector[1][15] ,
         \g_vector[1][13] , \g_vector[1][11] , \g_vector[1][9] ,
         \g_vector[1][7] , \g_vector[1][5] , \g_vector[1][3] ,
         \g_vector[1][1] , \g_vector[0][63] , \g_vector[0][62] ,
         \g_vector[0][61] , \g_vector[0][60] , \g_vector[0][59] ,
         \g_vector[0][58] , \g_vector[0][57] , \g_vector[0][56] ,
         \g_vector[0][55] , \g_vector[0][54] , \g_vector[0][53] ,
         \g_vector[0][52] , \g_vector[0][51] , \g_vector[0][50] ,
         \g_vector[0][49] , \g_vector[0][48] , \g_vector[0][47] ,
         \g_vector[0][46] , \g_vector[0][45] , \g_vector[0][44] ,
         \g_vector[0][43] , \g_vector[0][42] , \g_vector[0][41] ,
         \g_vector[0][40] , \g_vector[0][39] , \g_vector[0][38] ,
         \g_vector[0][37] , \g_vector[0][36] , \g_vector[0][35] ,
         \g_vector[0][34] , \g_vector[0][33] , \g_vector[0][32] ,
         \g_vector[0][31] , \g_vector[0][30] , \g_vector[0][29] ,
         \g_vector[0][28] , \g_vector[0][27] , \g_vector[0][26] ,
         \g_vector[0][25] , \g_vector[0][24] , \g_vector[0][23] ,
         \g_vector[0][22] , \g_vector[0][21] , \g_vector[0][20] ,
         \g_vector[0][19] , \g_vector[0][18] , \g_vector[0][17] ,
         \g_vector[0][16] , \g_vector[0][15] , \g_vector[0][14] ,
         \g_vector[0][13] , \g_vector[0][12] , \g_vector[0][11] ,
         \g_vector[0][10] , \g_vector[0][9] , \g_vector[0][8] ,
         \g_vector[0][7] , \g_vector[0][6] , \g_vector[0][5] ,
         \g_vector[0][4] , \g_vector[0][3] , \g_vector[0][2] ,
         \g_vector[0][1] , \g_vector[0][0] , \p_vector[5][63] ,
         \p_vector[5][59] , \p_vector[5][55] , \p_vector[5][51] ,
         \p_vector[4][63] , \p_vector[4][59] , \p_vector[4][47] ,
         \p_vector[4][43] , \p_vector[4][31] , \p_vector[4][27] ,
         \p_vector[3][63] , \p_vector[3][55] , \p_vector[3][47] ,
         \p_vector[3][39] , \p_vector[3][31] , \p_vector[3][23] ,
         \p_vector[3][15] , \p_vector[2][63] , \p_vector[2][59] ,
         \p_vector[2][55] , \p_vector[2][51] , \p_vector[2][47] ,
         \p_vector[2][43] , \p_vector[2][39] , \p_vector[2][35] ,
         \p_vector[2][31] , \p_vector[2][27] , \p_vector[2][23] ,
         \p_vector[2][19] , \p_vector[2][15] , \p_vector[2][11] ,
         \p_vector[2][7] , \p_vector[1][63] , \p_vector[1][61] ,
         \p_vector[1][59] , \p_vector[1][57] , \p_vector[1][55] ,
         \p_vector[1][53] , \p_vector[1][51] , \p_vector[1][49] ,
         \p_vector[1][47] , \p_vector[1][45] , \p_vector[1][43] ,
         \p_vector[1][41] , \p_vector[1][39] , \p_vector[1][37] ,
         \p_vector[1][35] , \p_vector[1][33] , \p_vector[1][31] ,
         \p_vector[1][29] , \p_vector[1][27] , \p_vector[1][25] ,
         \p_vector[1][23] , \p_vector[1][21] , \p_vector[1][19] ,
         \p_vector[1][17] , \p_vector[1][15] , \p_vector[1][13] ,
         \p_vector[1][11] , \p_vector[1][9] , \p_vector[1][7] ,
         \p_vector[1][5] , \p_vector[1][3] , \p_vector[0][63] ,
         \p_vector[0][62] , \p_vector[0][61] , \p_vector[0][60] ,
         \p_vector[0][59] , \p_vector[0][58] , \p_vector[0][57] ,
         \p_vector[0][56] , \p_vector[0][55] , \p_vector[0][54] ,
         \p_vector[0][53] , \p_vector[0][52] , \p_vector[0][51] ,
         \p_vector[0][50] , \p_vector[0][49] , \p_vector[0][48] ,
         \p_vector[0][47] , \p_vector[0][46] , \p_vector[0][45] ,
         \p_vector[0][44] , \p_vector[0][43] , \p_vector[0][42] ,
         \p_vector[0][41] , \p_vector[0][40] , \p_vector[0][39] ,
         \p_vector[0][38] , \p_vector[0][37] , \p_vector[0][36] ,
         \p_vector[0][35] , \p_vector[0][34] , \p_vector[0][33] ,
         \p_vector[0][32] , \p_vector[0][31] , \p_vector[0][30] ,
         \p_vector[0][29] , \p_vector[0][28] , \p_vector[0][27] ,
         \p_vector[0][26] , \p_vector[0][25] , \p_vector[0][24] ,
         \p_vector[0][23] , \p_vector[0][22] , \p_vector[0][21] ,
         \p_vector[0][20] , \p_vector[0][19] , \p_vector[0][18] ,
         \p_vector[0][17] , \p_vector[0][16] , \p_vector[0][15] ,
         \p_vector[0][14] , \p_vector[0][13] , \p_vector[0][12] ,
         \p_vector[0][11] , \p_vector[0][10] , \p_vector[0][9] ,
         \p_vector[0][8] , \p_vector[0][7] , \p_vector[0][6] ,
         \p_vector[0][5] , \p_vector[0][4] , \p_vector[0][3] ,
         \p_vector[0][2] , \p_vector[0][1] , n1, n2, n4;

  pg_net_126 pg_network_63 ( .a(A[63]), .b(B[63]), .p(\p_vector[0][63] ), .g(
        \g_vector[0][63] ) );
  pg_net_125 pg_network_62 ( .a(A[62]), .b(B[62]), .p(\p_vector[0][62] ), .g(
        \g_vector[0][62] ) );
  pg_net_124 pg_network_61 ( .a(A[61]), .b(B[61]), .p(\p_vector[0][61] ), .g(
        \g_vector[0][61] ) );
  pg_net_123 pg_network_60 ( .a(A[60]), .b(B[60]), .p(\p_vector[0][60] ), .g(
        \g_vector[0][60] ) );
  pg_net_122 pg_network_59 ( .a(A[59]), .b(B[59]), .p(\p_vector[0][59] ), .g(
        \g_vector[0][59] ) );
  pg_net_121 pg_network_58 ( .a(A[58]), .b(B[58]), .p(\p_vector[0][58] ), .g(
        \g_vector[0][58] ) );
  pg_net_120 pg_network_57 ( .a(A[57]), .b(B[57]), .p(\p_vector[0][57] ), .g(
        \g_vector[0][57] ) );
  pg_net_119 pg_network_56 ( .a(A[56]), .b(B[56]), .p(\p_vector[0][56] ), .g(
        \g_vector[0][56] ) );
  pg_net_118 pg_network_55 ( .a(A[55]), .b(B[55]), .p(\p_vector[0][55] ), .g(
        \g_vector[0][55] ) );
  pg_net_117 pg_network_54 ( .a(A[54]), .b(B[54]), .p(\p_vector[0][54] ), .g(
        \g_vector[0][54] ) );
  pg_net_116 pg_network_53 ( .a(A[53]), .b(B[53]), .p(\p_vector[0][53] ), .g(
        \g_vector[0][53] ) );
  pg_net_115 pg_network_52 ( .a(A[52]), .b(B[52]), .p(\p_vector[0][52] ), .g(
        \g_vector[0][52] ) );
  pg_net_114 pg_network_51 ( .a(A[51]), .b(B[51]), .p(\p_vector[0][51] ), .g(
        \g_vector[0][51] ) );
  pg_net_113 pg_network_50 ( .a(A[50]), .b(B[50]), .p(\p_vector[0][50] ), .g(
        \g_vector[0][50] ) );
  pg_net_112 pg_network_49 ( .a(A[49]), .b(B[49]), .p(\p_vector[0][49] ), .g(
        \g_vector[0][49] ) );
  pg_net_111 pg_network_48 ( .a(A[48]), .b(B[48]), .p(\p_vector[0][48] ), .g(
        \g_vector[0][48] ) );
  pg_net_110 pg_network_47 ( .a(A[47]), .b(B[47]), .p(\p_vector[0][47] ), .g(
        \g_vector[0][47] ) );
  pg_net_109 pg_network_46 ( .a(A[46]), .b(B[46]), .p(\p_vector[0][46] ), .g(
        \g_vector[0][46] ) );
  pg_net_108 pg_network_45 ( .a(A[45]), .b(B[45]), .p(\p_vector[0][45] ), .g(
        \g_vector[0][45] ) );
  pg_net_107 pg_network_44 ( .a(A[44]), .b(B[44]), .p(\p_vector[0][44] ), .g(
        \g_vector[0][44] ) );
  pg_net_106 pg_network_43 ( .a(A[43]), .b(B[43]), .p(\p_vector[0][43] ), .g(
        \g_vector[0][43] ) );
  pg_net_105 pg_network_42 ( .a(A[42]), .b(B[42]), .p(\p_vector[0][42] ), .g(
        \g_vector[0][42] ) );
  pg_net_104 pg_network_41 ( .a(A[41]), .b(B[41]), .p(\p_vector[0][41] ), .g(
        \g_vector[0][41] ) );
  pg_net_103 pg_network_40 ( .a(A[40]), .b(B[40]), .p(\p_vector[0][40] ), .g(
        \g_vector[0][40] ) );
  pg_net_102 pg_network_39 ( .a(A[39]), .b(B[39]), .p(\p_vector[0][39] ), .g(
        \g_vector[0][39] ) );
  pg_net_101 pg_network_38 ( .a(A[38]), .b(B[38]), .p(\p_vector[0][38] ), .g(
        \g_vector[0][38] ) );
  pg_net_100 pg_network_37 ( .a(A[37]), .b(B[37]), .p(\p_vector[0][37] ), .g(
        \g_vector[0][37] ) );
  pg_net_99 pg_network_36 ( .a(A[36]), .b(B[36]), .p(\p_vector[0][36] ), .g(
        \g_vector[0][36] ) );
  pg_net_98 pg_network_35 ( .a(A[35]), .b(B[35]), .p(\p_vector[0][35] ), .g(
        \g_vector[0][35] ) );
  pg_net_97 pg_network_34 ( .a(A[34]), .b(B[34]), .p(\p_vector[0][34] ), .g(
        \g_vector[0][34] ) );
  pg_net_96 pg_network_33 ( .a(A[33]), .b(B[33]), .p(\p_vector[0][33] ), .g(
        \g_vector[0][33] ) );
  pg_net_95 pg_network_32 ( .a(A[32]), .b(B[32]), .p(\p_vector[0][32] ), .g(
        \g_vector[0][32] ) );
  pg_net_94 pg_network_31 ( .a(A[31]), .b(B[31]), .p(\p_vector[0][31] ), .g(
        \g_vector[0][31] ) );
  pg_net_93 pg_network_30 ( .a(A[30]), .b(B[30]), .p(\p_vector[0][30] ), .g(
        \g_vector[0][30] ) );
  pg_net_92 pg_network_29 ( .a(A[29]), .b(B[29]), .p(\p_vector[0][29] ), .g(
        \g_vector[0][29] ) );
  pg_net_91 pg_network_28 ( .a(A[28]), .b(B[28]), .p(\p_vector[0][28] ), .g(
        \g_vector[0][28] ) );
  pg_net_90 pg_network_27 ( .a(A[27]), .b(B[27]), .p(\p_vector[0][27] ), .g(
        \g_vector[0][27] ) );
  pg_net_89 pg_network_26 ( .a(A[26]), .b(B[26]), .p(\p_vector[0][26] ), .g(
        \g_vector[0][26] ) );
  pg_net_88 pg_network_25 ( .a(A[25]), .b(B[25]), .p(\p_vector[0][25] ), .g(
        \g_vector[0][25] ) );
  pg_net_87 pg_network_24 ( .a(A[24]), .b(B[24]), .p(\p_vector[0][24] ), .g(
        \g_vector[0][24] ) );
  pg_net_86 pg_network_23 ( .a(A[23]), .b(B[23]), .p(\p_vector[0][23] ), .g(
        \g_vector[0][23] ) );
  pg_net_85 pg_network_22 ( .a(A[22]), .b(B[22]), .p(\p_vector[0][22] ), .g(
        \g_vector[0][22] ) );
  pg_net_84 pg_network_21 ( .a(A[21]), .b(B[21]), .p(\p_vector[0][21] ), .g(
        \g_vector[0][21] ) );
  pg_net_83 pg_network_20 ( .a(A[20]), .b(B[20]), .p(\p_vector[0][20] ), .g(
        \g_vector[0][20] ) );
  pg_net_82 pg_network_19 ( .a(A[19]), .b(B[19]), .p(\p_vector[0][19] ), .g(
        \g_vector[0][19] ) );
  pg_net_81 pg_network_18 ( .a(A[18]), .b(B[18]), .p(\p_vector[0][18] ), .g(
        \g_vector[0][18] ) );
  pg_net_80 pg_network_17 ( .a(A[17]), .b(B[17]), .p(\p_vector[0][17] ), .g(
        \g_vector[0][17] ) );
  pg_net_79 pg_network_16 ( .a(A[16]), .b(B[16]), .p(\p_vector[0][16] ), .g(
        \g_vector[0][16] ) );
  pg_net_78 pg_network_15 ( .a(A[15]), .b(B[15]), .p(\p_vector[0][15] ), .g(
        \g_vector[0][15] ) );
  pg_net_77 pg_network_14 ( .a(A[14]), .b(B[14]), .p(\p_vector[0][14] ), .g(
        \g_vector[0][14] ) );
  pg_net_76 pg_network_13 ( .a(A[13]), .b(B[13]), .p(\p_vector[0][13] ), .g(
        \g_vector[0][13] ) );
  pg_net_75 pg_network_12 ( .a(A[12]), .b(B[12]), .p(\p_vector[0][12] ), .g(
        \g_vector[0][12] ) );
  pg_net_74 pg_network_11 ( .a(A[11]), .b(B[11]), .p(\p_vector[0][11] ), .g(
        \g_vector[0][11] ) );
  pg_net_73 pg_network_10 ( .a(A[10]), .b(B[10]), .p(\p_vector[0][10] ), .g(
        \g_vector[0][10] ) );
  pg_net_72 pg_network_9 ( .a(A[9]), .b(B[9]), .p(\p_vector[0][9] ), .g(
        \g_vector[0][9] ) );
  pg_net_71 pg_network_8 ( .a(A[8]), .b(B[8]), .p(\p_vector[0][8] ), .g(
        \g_vector[0][8] ) );
  pg_net_70 pg_network_7 ( .a(A[7]), .b(B[7]), .p(\p_vector[0][7] ), .g(
        \g_vector[0][7] ) );
  pg_net_69 pg_network_6 ( .a(A[6]), .b(B[6]), .p(\p_vector[0][6] ), .g(
        \g_vector[0][6] ) );
  pg_net_68 pg_network_5 ( .a(A[5]), .b(B[5]), .p(\p_vector[0][5] ), .g(
        \g_vector[0][5] ) );
  pg_net_67 pg_network_4 ( .a(A[4]), .b(B[4]), .p(\p_vector[0][4] ), .g(
        \g_vector[0][4] ) );
  pg_net_66 pg_network_3 ( .a(A[3]), .b(B[3]), .p(\p_vector[0][3] ), .g(
        \g_vector[0][3] ) );
  pg_net_65 pg_network_2 ( .a(A[2]), .b(B[2]), .p(\p_vector[0][2] ), .g(
        \g_vector[0][2] ) );
  pg_net_64 pg_network_1 ( .a(A[1]), .b(B[1]), .p(\p_vector[0][1] ), .g(
        \g_vector[0][1] ) );
  PG_BLOCK_126 std_PG_1_63 ( .p2(\p_vector[0][63] ), .g2(\g_vector[0][63] ), 
        .p1(\p_vector[0][62] ), .g1(\g_vector[0][62] ), .PG_P(
        \p_vector[1][63] ), .PG_G(\g_vector[1][63] ) );
  PG_BLOCK_125 std_PG_1_61 ( .p2(\p_vector[0][61] ), .g2(\g_vector[0][61] ), 
        .p1(\p_vector[0][60] ), .g1(\g_vector[0][60] ), .PG_P(
        \p_vector[1][61] ), .PG_G(\g_vector[1][61] ) );
  PG_BLOCK_124 std_PG_1_59 ( .p2(\p_vector[0][59] ), .g2(\g_vector[0][59] ), 
        .p1(\p_vector[0][58] ), .g1(\g_vector[0][58] ), .PG_P(
        \p_vector[1][59] ), .PG_G(\g_vector[1][59] ) );
  PG_BLOCK_123 std_PG_1_57 ( .p2(\p_vector[0][57] ), .g2(\g_vector[0][57] ), 
        .p1(\p_vector[0][56] ), .g1(\g_vector[0][56] ), .PG_P(
        \p_vector[1][57] ), .PG_G(\g_vector[1][57] ) );
  PG_BLOCK_122 std_PG_1_55 ( .p2(\p_vector[0][55] ), .g2(\g_vector[0][55] ), 
        .p1(\p_vector[0][54] ), .g1(\g_vector[0][54] ), .PG_P(
        \p_vector[1][55] ), .PG_G(\g_vector[1][55] ) );
  PG_BLOCK_121 std_PG_1_53 ( .p2(\p_vector[0][53] ), .g2(\g_vector[0][53] ), 
        .p1(\p_vector[0][52] ), .g1(\g_vector[0][52] ), .PG_P(
        \p_vector[1][53] ), .PG_G(\g_vector[1][53] ) );
  PG_BLOCK_120 std_PG_1_51 ( .p2(\p_vector[0][51] ), .g2(\g_vector[0][51] ), 
        .p1(\p_vector[0][50] ), .g1(\g_vector[0][50] ), .PG_P(
        \p_vector[1][51] ), .PG_G(\g_vector[1][51] ) );
  PG_BLOCK_119 std_PG_1_49 ( .p2(\p_vector[0][49] ), .g2(\g_vector[0][49] ), 
        .p1(\p_vector[0][48] ), .g1(\g_vector[0][48] ), .PG_P(
        \p_vector[1][49] ), .PG_G(\g_vector[1][49] ) );
  PG_BLOCK_118 std_PG_1_47 ( .p2(\p_vector[0][47] ), .g2(\g_vector[0][47] ), 
        .p1(\p_vector[0][46] ), .g1(\g_vector[0][46] ), .PG_P(
        \p_vector[1][47] ), .PG_G(\g_vector[1][47] ) );
  PG_BLOCK_117 std_PG_1_45 ( .p2(\p_vector[0][45] ), .g2(\g_vector[0][45] ), 
        .p1(\p_vector[0][44] ), .g1(\g_vector[0][44] ), .PG_P(
        \p_vector[1][45] ), .PG_G(\g_vector[1][45] ) );
  PG_BLOCK_116 std_PG_1_43 ( .p2(\p_vector[0][43] ), .g2(\g_vector[0][43] ), 
        .p1(\p_vector[0][42] ), .g1(\g_vector[0][42] ), .PG_P(
        \p_vector[1][43] ), .PG_G(\g_vector[1][43] ) );
  PG_BLOCK_115 std_PG_1_41 ( .p2(\p_vector[0][41] ), .g2(\g_vector[0][41] ), 
        .p1(\p_vector[0][40] ), .g1(\g_vector[0][40] ), .PG_P(
        \p_vector[1][41] ), .PG_G(\g_vector[1][41] ) );
  PG_BLOCK_114 std_PG_1_39 ( .p2(\p_vector[0][39] ), .g2(\g_vector[0][39] ), 
        .p1(\p_vector[0][38] ), .g1(\g_vector[0][38] ), .PG_P(
        \p_vector[1][39] ), .PG_G(\g_vector[1][39] ) );
  PG_BLOCK_113 std_PG_1_37 ( .p2(\p_vector[0][37] ), .g2(\g_vector[0][37] ), 
        .p1(\p_vector[0][36] ), .g1(\g_vector[0][36] ), .PG_P(
        \p_vector[1][37] ), .PG_G(\g_vector[1][37] ) );
  PG_BLOCK_112 std_PG_1_35 ( .p2(\p_vector[0][35] ), .g2(\g_vector[0][35] ), 
        .p1(\p_vector[0][34] ), .g1(\g_vector[0][34] ), .PG_P(
        \p_vector[1][35] ), .PG_G(\g_vector[1][35] ) );
  PG_BLOCK_111 std_PG_1_33 ( .p2(\p_vector[0][33] ), .g2(\g_vector[0][33] ), 
        .p1(\p_vector[0][32] ), .g1(\g_vector[0][32] ), .PG_P(
        \p_vector[1][33] ), .PG_G(\g_vector[1][33] ) );
  PG_BLOCK_110 std_PG_1_31 ( .p2(\p_vector[0][31] ), .g2(\g_vector[0][31] ), 
        .p1(\p_vector[0][30] ), .g1(\g_vector[0][30] ), .PG_P(
        \p_vector[1][31] ), .PG_G(\g_vector[1][31] ) );
  PG_BLOCK_109 std_PG_1_29 ( .p2(\p_vector[0][29] ), .g2(\g_vector[0][29] ), 
        .p1(\p_vector[0][28] ), .g1(\g_vector[0][28] ), .PG_P(
        \p_vector[1][29] ), .PG_G(\g_vector[1][29] ) );
  PG_BLOCK_108 std_PG_1_27 ( .p2(\p_vector[0][27] ), .g2(\g_vector[0][27] ), 
        .p1(\p_vector[0][26] ), .g1(\g_vector[0][26] ), .PG_P(
        \p_vector[1][27] ), .PG_G(\g_vector[1][27] ) );
  PG_BLOCK_107 std_PG_1_25 ( .p2(\p_vector[0][25] ), .g2(\g_vector[0][25] ), 
        .p1(\p_vector[0][24] ), .g1(\g_vector[0][24] ), .PG_P(
        \p_vector[1][25] ), .PG_G(\g_vector[1][25] ) );
  PG_BLOCK_106 std_PG_1_23 ( .p2(\p_vector[0][23] ), .g2(\g_vector[0][23] ), 
        .p1(\p_vector[0][22] ), .g1(\g_vector[0][22] ), .PG_P(
        \p_vector[1][23] ), .PG_G(\g_vector[1][23] ) );
  PG_BLOCK_105 std_PG_1_21 ( .p2(\p_vector[0][21] ), .g2(\g_vector[0][21] ), 
        .p1(\p_vector[0][20] ), .g1(\g_vector[0][20] ), .PG_P(
        \p_vector[1][21] ), .PG_G(\g_vector[1][21] ) );
  PG_BLOCK_104 std_PG_1_19 ( .p2(\p_vector[0][19] ), .g2(\g_vector[0][19] ), 
        .p1(\p_vector[0][18] ), .g1(\g_vector[0][18] ), .PG_P(
        \p_vector[1][19] ), .PG_G(\g_vector[1][19] ) );
  PG_BLOCK_103 std_PG_1_17 ( .p2(\p_vector[0][17] ), .g2(\g_vector[0][17] ), 
        .p1(\p_vector[0][16] ), .g1(\g_vector[0][16] ), .PG_P(
        \p_vector[1][17] ), .PG_G(\g_vector[1][17] ) );
  PG_BLOCK_102 std_PG_1_15 ( .p2(\p_vector[0][15] ), .g2(\g_vector[0][15] ), 
        .p1(\p_vector[0][14] ), .g1(\g_vector[0][14] ), .PG_P(
        \p_vector[1][15] ), .PG_G(\g_vector[1][15] ) );
  PG_BLOCK_101 std_PG_1_13 ( .p2(\p_vector[0][13] ), .g2(\g_vector[0][13] ), 
        .p1(\p_vector[0][12] ), .g1(\g_vector[0][12] ), .PG_P(
        \p_vector[1][13] ), .PG_G(\g_vector[1][13] ) );
  PG_BLOCK_100 std_PG_1_11 ( .p2(\p_vector[0][11] ), .g2(\g_vector[0][11] ), 
        .p1(\p_vector[0][10] ), .g1(\g_vector[0][10] ), .PG_P(
        \p_vector[1][11] ), .PG_G(\g_vector[1][11] ) );
  PG_BLOCK_99 std_PG_1_9 ( .p2(\p_vector[0][9] ), .g2(\g_vector[0][9] ), .p1(
        \p_vector[0][8] ), .g1(\g_vector[0][8] ), .PG_P(\p_vector[1][9] ), 
        .PG_G(\g_vector[1][9] ) );
  PG_BLOCK_98 std_PG_1_7 ( .p2(\p_vector[0][7] ), .g2(\g_vector[0][7] ), .p1(
        \p_vector[0][6] ), .g1(\g_vector[0][6] ), .PG_P(\p_vector[1][7] ), 
        .PG_G(\g_vector[1][7] ) );
  PG_BLOCK_97 std_PG_1_5 ( .p2(\p_vector[0][5] ), .g2(\g_vector[0][5] ), .p1(
        \p_vector[0][4] ), .g1(\g_vector[0][4] ), .PG_P(\p_vector[1][5] ), 
        .PG_G(\g_vector[1][5] ) );
  PG_BLOCK_96 std_PG_1_3 ( .p2(\p_vector[0][3] ), .g2(\g_vector[0][3] ), .p1(
        \p_vector[0][2] ), .g1(\g_vector[0][2] ), .PG_P(\p_vector[1][3] ), 
        .PG_G(\g_vector[1][3] ) );
  G_BLOCK_34 std_G_1_1 ( .p2(\p_vector[0][1] ), .g2(\g_vector[0][1] ), .g1(
        \g_vector[0][0] ), .G(\g_vector[1][1] ) );
  PG_BLOCK_95 std_PG_2_63 ( .p2(\p_vector[1][63] ), .g2(\g_vector[1][63] ), 
        .p1(\p_vector[1][61] ), .g1(\g_vector[1][61] ), .PG_P(
        \p_vector[2][63] ), .PG_G(\g_vector[2][63] ) );
  PG_BLOCK_94 std_PG_2_59 ( .p2(\p_vector[1][59] ), .g2(\g_vector[1][59] ), 
        .p1(\p_vector[1][57] ), .g1(\g_vector[1][57] ), .PG_P(
        \p_vector[2][59] ), .PG_G(\g_vector[2][59] ) );
  PG_BLOCK_93 std_PG_2_55 ( .p2(\p_vector[1][55] ), .g2(\g_vector[1][55] ), 
        .p1(\p_vector[1][53] ), .g1(\g_vector[1][53] ), .PG_P(
        \p_vector[2][55] ), .PG_G(\g_vector[2][55] ) );
  PG_BLOCK_92 std_PG_2_51 ( .p2(\p_vector[1][51] ), .g2(\g_vector[1][51] ), 
        .p1(\p_vector[1][49] ), .g1(\g_vector[1][49] ), .PG_P(
        \p_vector[2][51] ), .PG_G(\g_vector[2][51] ) );
  PG_BLOCK_91 std_PG_2_47 ( .p2(\p_vector[1][47] ), .g2(\g_vector[1][47] ), 
        .p1(\p_vector[1][45] ), .g1(\g_vector[1][45] ), .PG_P(
        \p_vector[2][47] ), .PG_G(\g_vector[2][47] ) );
  PG_BLOCK_90 std_PG_2_43 ( .p2(\p_vector[1][43] ), .g2(\g_vector[1][43] ), 
        .p1(\p_vector[1][41] ), .g1(\g_vector[1][41] ), .PG_P(
        \p_vector[2][43] ), .PG_G(\g_vector[2][43] ) );
  PG_BLOCK_89 std_PG_2_39 ( .p2(\p_vector[1][39] ), .g2(\g_vector[1][39] ), 
        .p1(\p_vector[1][37] ), .g1(\g_vector[1][37] ), .PG_P(
        \p_vector[2][39] ), .PG_G(\g_vector[2][39] ) );
  PG_BLOCK_88 std_PG_2_35 ( .p2(\p_vector[1][35] ), .g2(\g_vector[1][35] ), 
        .p1(\p_vector[1][33] ), .g1(\g_vector[1][33] ), .PG_P(
        \p_vector[2][35] ), .PG_G(\g_vector[2][35] ) );
  PG_BLOCK_87 std_PG_2_31 ( .p2(\p_vector[1][31] ), .g2(\g_vector[1][31] ), 
        .p1(\p_vector[1][29] ), .g1(\g_vector[1][29] ), .PG_P(
        \p_vector[2][31] ), .PG_G(\g_vector[2][31] ) );
  PG_BLOCK_86 std_PG_2_27 ( .p2(\p_vector[1][27] ), .g2(\g_vector[1][27] ), 
        .p1(\p_vector[1][25] ), .g1(\g_vector[1][25] ), .PG_P(
        \p_vector[2][27] ), .PG_G(\g_vector[2][27] ) );
  PG_BLOCK_85 std_PG_2_23 ( .p2(\p_vector[1][23] ), .g2(\g_vector[1][23] ), 
        .p1(\p_vector[1][21] ), .g1(\g_vector[1][21] ), .PG_P(
        \p_vector[2][23] ), .PG_G(\g_vector[2][23] ) );
  PG_BLOCK_84 std_PG_2_19 ( .p2(\p_vector[1][19] ), .g2(\g_vector[1][19] ), 
        .p1(\p_vector[1][17] ), .g1(\g_vector[1][17] ), .PG_P(
        \p_vector[2][19] ), .PG_G(\g_vector[2][19] ) );
  PG_BLOCK_83 std_PG_2_15 ( .p2(\p_vector[1][15] ), .g2(\g_vector[1][15] ), 
        .p1(\p_vector[1][13] ), .g1(\g_vector[1][13] ), .PG_P(
        \p_vector[2][15] ), .PG_G(\g_vector[2][15] ) );
  PG_BLOCK_82 std_PG_2_11 ( .p2(\p_vector[1][11] ), .g2(\g_vector[1][11] ), 
        .p1(\p_vector[1][9] ), .g1(\g_vector[1][9] ), .PG_P(\p_vector[2][11] ), 
        .PG_G(\g_vector[2][11] ) );
  PG_BLOCK_81 std_PG_2_7 ( .p2(\p_vector[1][7] ), .g2(\g_vector[1][7] ), .p1(
        \p_vector[1][5] ), .g1(\g_vector[1][5] ), .PG_P(\p_vector[2][7] ), 
        .PG_G(\g_vector[2][7] ) );
  G_BLOCK_33 std_G_2_3 ( .p2(\p_vector[1][3] ), .g2(\g_vector[1][3] ), .g1(
        \g_vector[1][1] ), .G(Co[0]) );
  PG_BLOCK_80 std_PG_3_63 ( .p2(\p_vector[2][63] ), .g2(\g_vector[2][63] ), 
        .p1(\p_vector[2][59] ), .g1(\g_vector[2][59] ), .PG_P(
        \p_vector[3][63] ), .PG_G(\g_vector[3][63] ) );
  PG_BLOCK_79 std_PG_3_55 ( .p2(\p_vector[2][55] ), .g2(\g_vector[2][55] ), 
        .p1(\p_vector[2][51] ), .g1(\g_vector[2][51] ), .PG_P(
        \p_vector[3][55] ), .PG_G(\g_vector[3][55] ) );
  PG_BLOCK_78 std_PG_3_47 ( .p2(\p_vector[2][47] ), .g2(\g_vector[2][47] ), 
        .p1(\p_vector[2][43] ), .g1(\g_vector[2][43] ), .PG_P(
        \p_vector[3][47] ), .PG_G(\g_vector[3][47] ) );
  PG_BLOCK_77 std_PG_3_39 ( .p2(\p_vector[2][39] ), .g2(\g_vector[2][39] ), 
        .p1(\p_vector[2][35] ), .g1(\g_vector[2][35] ), .PG_P(
        \p_vector[3][39] ), .PG_G(\g_vector[3][39] ) );
  PG_BLOCK_76 std_PG_3_31 ( .p2(\p_vector[2][31] ), .g2(\g_vector[2][31] ), 
        .p1(\p_vector[2][27] ), .g1(\g_vector[2][27] ), .PG_P(
        \p_vector[3][31] ), .PG_G(\g_vector[3][31] ) );
  PG_BLOCK_75 std_PG_3_23 ( .p2(\p_vector[2][23] ), .g2(\g_vector[2][23] ), 
        .p1(\p_vector[2][19] ), .g1(\g_vector[2][19] ), .PG_P(
        \p_vector[3][23] ), .PG_G(\g_vector[3][23] ) );
  PG_BLOCK_74 std_PG_3_15 ( .p2(\p_vector[2][15] ), .g2(\g_vector[2][15] ), 
        .p1(\p_vector[2][11] ), .g1(\g_vector[2][11] ), .PG_P(
        \p_vector[3][15] ), .PG_G(\g_vector[3][15] ) );
  G_BLOCK_32 std_G_3_7 ( .p2(\p_vector[2][7] ), .g2(\g_vector[2][7] ), .g1(
        Co[0]), .G(Co[1]) );
  PG_BLOCK_73 std_PG_4_63 ( .p2(\p_vector[3][63] ), .g2(\g_vector[3][63] ), 
        .p1(\p_vector[3][55] ), .g1(\g_vector[3][55] ), .PG_P(
        \p_vector[4][63] ), .PG_G(\g_vector[4][63] ) );
  PG_BLOCK_72 add_PG_4_63_1 ( .p2(\p_vector[2][59] ), .g2(\g_vector[2][59] ), 
        .p1(\p_vector[3][55] ), .g1(\g_vector[3][55] ), .PG_P(
        \p_vector[4][59] ), .PG_G(\g_vector[4][59] ) );
  PG_BLOCK_71 std_PG_4_47 ( .p2(\p_vector[3][47] ), .g2(\g_vector[3][47] ), 
        .p1(\p_vector[3][39] ), .g1(\g_vector[3][39] ), .PG_P(
        \p_vector[4][47] ), .PG_G(\g_vector[4][47] ) );
  PG_BLOCK_70 add_PG_4_47_1 ( .p2(\p_vector[2][43] ), .g2(\g_vector[2][43] ), 
        .p1(\p_vector[3][39] ), .g1(\g_vector[3][39] ), .PG_P(
        \p_vector[4][43] ), .PG_G(\g_vector[4][43] ) );
  PG_BLOCK_69 std_PG_4_31 ( .p2(\p_vector[3][31] ), .g2(\g_vector[3][31] ), 
        .p1(\p_vector[3][23] ), .g1(\g_vector[3][23] ), .PG_P(
        \p_vector[4][31] ), .PG_G(\g_vector[4][31] ) );
  PG_BLOCK_68 add_PG_4_31_1 ( .p2(\p_vector[2][27] ), .g2(\g_vector[2][27] ), 
        .p1(\p_vector[3][23] ), .g1(\g_vector[3][23] ), .PG_P(
        \p_vector[4][27] ), .PG_G(\g_vector[4][27] ) );
  G_BLOCK_31 std_G_4_15 ( .p2(\p_vector[3][15] ), .g2(\g_vector[3][15] ), .g1(
        Co[1]), .G(Co[3]) );
  G_BLOCK_30 add_G_4_15_1 ( .p2(\p_vector[2][11] ), .g2(\g_vector[2][11] ), 
        .g1(Co[1]), .G(Co[2]) );
  PG_BLOCK_67 std_PG_5_63 ( .p2(\p_vector[4][63] ), .g2(\g_vector[4][63] ), 
        .p1(\p_vector[4][47] ), .g1(\g_vector[4][47] ), .PG_P(
        \p_vector[5][63] ), .PG_G(\g_vector[5][63] ) );
  PG_BLOCK_66 add_PG_5_63_1 ( .p2(\p_vector[4][59] ), .g2(\g_vector[4][59] ), 
        .p1(\p_vector[4][47] ), .g1(\g_vector[4][47] ), .PG_P(
        \p_vector[5][59] ), .PG_G(\g_vector[5][59] ) );
  PG_BLOCK_65 add_PG_5_63_2 ( .p2(\p_vector[3][55] ), .g2(\g_vector[3][55] ), 
        .p1(\p_vector[4][47] ), .g1(\g_vector[4][47] ), .PG_P(
        \p_vector[5][55] ), .PG_G(\g_vector[5][55] ) );
  PG_BLOCK_64 add_PG_5_63_3 ( .p2(\p_vector[2][51] ), .g2(\g_vector[2][51] ), 
        .p1(\p_vector[4][47] ), .g1(\g_vector[4][47] ), .PG_P(
        \p_vector[5][51] ), .PG_G(\g_vector[5][51] ) );
  G_BLOCK_29 std_G_5_31 ( .p2(\p_vector[4][31] ), .g2(\g_vector[4][31] ), .g1(
        Co[3]), .G(Co[7]) );
  G_BLOCK_28 add_G_5_31_1 ( .p2(\p_vector[4][27] ), .g2(\g_vector[4][27] ), 
        .g1(Co[3]), .G(Co[6]) );
  G_BLOCK_27 add_G_5_31_2 ( .p2(\p_vector[3][23] ), .g2(\g_vector[3][23] ), 
        .g1(Co[3]), .G(Co[5]) );
  G_BLOCK_26 add_G_5_31_3 ( .p2(\p_vector[2][19] ), .g2(\g_vector[2][19] ), 
        .g1(Co[3]), .G(Co[4]) );
  G_BLOCK_25 std_G_6_63 ( .p2(\p_vector[5][63] ), .g2(\g_vector[5][63] ), .g1(
        Co[7]), .G(Co[15]) );
  G_BLOCK_24 add_G_6_63_1 ( .p2(\p_vector[5][59] ), .g2(\g_vector[5][59] ), 
        .g1(Co[7]), .G(Co[14]) );
  G_BLOCK_23 add_G_6_63_2 ( .p2(\p_vector[5][55] ), .g2(\g_vector[5][55] ), 
        .g1(Co[7]), .G(Co[13]) );
  G_BLOCK_22 add_G_6_63_3 ( .p2(\p_vector[5][51] ), .g2(\g_vector[5][51] ), 
        .g1(Co[7]), .G(Co[12]) );
  G_BLOCK_21 add_G_6_63_4 ( .p2(\p_vector[4][47] ), .g2(\g_vector[4][47] ), 
        .g1(Co[7]), .G(Co[11]) );
  G_BLOCK_20 add_G_6_63_5 ( .p2(\p_vector[4][43] ), .g2(\g_vector[4][43] ), 
        .g1(Co[7]), .G(Co[10]) );
  G_BLOCK_19 add_G_6_63_6 ( .p2(\p_vector[3][39] ), .g2(\g_vector[3][39] ), 
        .g1(Co[7]), .G(Co[9]) );
  G_BLOCK_18 add_G_6_63_7 ( .p2(\p_vector[2][35] ), .g2(\g_vector[2][35] ), 
        .g1(Co[7]), .G(Co[8]) );
  OAI21_X1 U1 ( .B1(n2), .B2(n1), .A(n4), .ZN(\g_vector[0][0] ) );
  OAI21_X1 U2 ( .B1(A[0]), .B2(B[0]), .A(Cin), .ZN(n4) );
  INV_X1 U3 ( .A(A[0]), .ZN(n2) );
  INV_X1 U4 ( .A(B[0]), .ZN(n1) );
endmodule


module FA_256 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_255 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_254 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_253 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_64 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_256 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_255 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_254 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_253 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_252 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_251 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_250 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_249 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_63 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_252 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_251 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_250 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_249 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_128 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_127 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_126 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_125 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_GENERIC_NBIT4_32 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_128 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_127 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_126 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_125 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_32 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_64 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_63 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_32 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module FA_248 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_247 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_246 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_245 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_62 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_248 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_247 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_246 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_245 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_244 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_243 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_242 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_241 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_61 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_244 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_243 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_242 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_241 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_124 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_123 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_122 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_121 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_GENERIC_NBIT4_31 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_124 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_123 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_122 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_121 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_31 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_62 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_61 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_31 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module FA_240 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_239 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_238 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_237 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_60 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_240 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_239 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_238 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_237 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_236 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_235 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_234 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_233 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_59 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_236 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_235 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_234 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_233 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_120 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_119 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_118 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_117 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_GENERIC_NBIT4_30 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_120 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_119 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_118 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_117 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_30 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_60 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_59 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_30 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module FA_232 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_231 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_230 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_229 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_58 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_232 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_231 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_230 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_229 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_228 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_227 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_226 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_225 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_57 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_228 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_227 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_226 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_225 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_116 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_115 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_114 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_113 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_GENERIC_NBIT4_29 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_116 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_115 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_114 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_113 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_29 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_58 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_57 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_29 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module FA_224 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_223 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_222 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_221 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_56 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_224 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_223 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_222 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_221 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_220 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_219 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_218 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_217 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_55 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_220 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_219 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_218 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_217 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_112 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_111 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_110 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_109 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_GENERIC_NBIT4_28 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_112 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_111 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_110 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_109 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_28 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_56 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_55 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_28 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module FA_216 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_215 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_214 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_213 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_54 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_216 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_215 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_214 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_213 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_212 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_211 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_210 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_209 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_53 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_212 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_211 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_210 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_209 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_108 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_107 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_106 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_105 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_GENERIC_NBIT4_27 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_108 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_107 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_106 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_105 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_27 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_54 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_53 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_27 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module FA_208 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_207 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_206 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_205 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_52 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_208 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_207 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_206 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_205 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_204 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_203 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_202 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_201 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_51 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_204 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_203 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_202 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_201 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_104 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_103 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_102 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_101 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_GENERIC_NBIT4_26 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_104 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_103 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_102 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_101 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_26 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_52 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_51 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_26 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module FA_200 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_199 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_198 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_197 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_50 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_200 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_199 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_198 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_197 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_196 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_195 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_194 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_193 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_49 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_196 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_195 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_194 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_193 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_100 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_99 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_98 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_97 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_GENERIC_NBIT4_25 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_100 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_99 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_98 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_97 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_25 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_50 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_49 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_25 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module FA_192 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_191 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_190 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_189 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_48 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_192 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_191 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_190 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_189 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_188 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_187 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_186 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_185 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_47 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_188 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_187 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_186 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_185 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_96 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_95 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_94 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_93 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_GENERIC_NBIT4_24 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_96 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_95 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_94 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_93 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_24 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_48 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_47 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_24 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module FA_184 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_183 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_182 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_181 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_46 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_184 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_183 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_182 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_181 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_180 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_179 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_178 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_177 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_45 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_180 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_179 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_178 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_177 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_92 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_91 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_90 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_89 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_GENERIC_NBIT4_23 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_92 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_91 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_90 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_89 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_23 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_46 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_45 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_23 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module FA_176 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_175 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_174 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_173 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_44 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_176 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_175 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_174 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_173 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_172 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_171 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_170 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_169 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_43 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_172 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_171 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_170 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_169 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_88 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_87 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_86 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_85 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_GENERIC_NBIT4_22 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_88 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_87 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_86 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_85 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_22 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_44 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_43 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_22 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module FA_168 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_167 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_166 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_165 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_42 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_168 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_167 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_166 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_165 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_164 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_163 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_162 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_161 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_41 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_164 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_163 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_162 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_161 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_84 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_83 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_82 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_81 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_GENERIC_NBIT4_21 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_84 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_83 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_82 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_81 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_21 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_42 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_41 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_21 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module FA_160 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_159 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_158 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_157 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_40 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_160 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_159 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_158 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_157 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_156 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_155 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_154 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_153 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_39 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_156 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_155 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_154 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_153 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_80 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_79 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_78 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_77 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_GENERIC_NBIT4_20 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_80 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_79 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_78 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_77 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_20 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_40 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_39 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_20 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module FA_152 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_151 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_150 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_149 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_38 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_152 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_151 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_150 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_149 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_148 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_147 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_146 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_145 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_37 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_148 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_147 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_146 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_145 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_76 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_75 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_74 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_73 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_GENERIC_NBIT4_19 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_76 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_75 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_74 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_73 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_19 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_38 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_37 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_19 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module FA_144 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_143 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_142 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_141 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_36 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_144 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_143 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_142 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_141 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_140 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_139 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_138 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_137 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_35 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_140 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_139 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_138 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_137 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_72 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_71 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_70 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_69 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_GENERIC_NBIT4_18 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_72 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_71 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_70 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_69 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_18 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_36 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_35 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_18 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module FA_136 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_135 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_134 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_133 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_34 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_136 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_135 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_134 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_133 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_132 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_131 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_130 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_129 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_33 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_132 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_131 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_130 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_129 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_68 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_67 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_66 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_65 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(S), .ZN(n2) );
  INV_X1 U2 ( .A(n4), .ZN(Y) );
  AOI22_X1 U3 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
endmodule


module MUX21_GENERIC_NBIT4_17 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_68 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_67 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_66 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_65 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_17 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_34 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_33 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_17 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module sum_generator_n_bit64_n_CSB16_2 ( A, B, C_in, S );
  input [63:0] A;
  input [63:0] B;
  input [15:0] C_in;
  output [63:0] S;


  carry_select_block_n4_32 csb_0 ( .A(A[3:0]), .B(B[3:0]), .C_sel(C_in[0]), 
        .S(S[3:0]) );
  carry_select_block_n4_31 csb_1 ( .A(A[7:4]), .B(B[7:4]), .C_sel(C_in[1]), 
        .S(S[7:4]) );
  carry_select_block_n4_30 csb_2 ( .A(A[11:8]), .B(B[11:8]), .C_sel(C_in[2]), 
        .S(S[11:8]) );
  carry_select_block_n4_29 csb_3 ( .A(A[15:12]), .B(B[15:12]), .C_sel(C_in[3]), 
        .S(S[15:12]) );
  carry_select_block_n4_28 csb_4 ( .A(A[19:16]), .B(B[19:16]), .C_sel(C_in[4]), 
        .S(S[19:16]) );
  carry_select_block_n4_27 csb_5 ( .A(A[23:20]), .B(B[23:20]), .C_sel(C_in[5]), 
        .S(S[23:20]) );
  carry_select_block_n4_26 csb_6 ( .A(A[27:24]), .B(B[27:24]), .C_sel(C_in[6]), 
        .S(S[27:24]) );
  carry_select_block_n4_25 csb_7 ( .A(A[31:28]), .B(B[31:28]), .C_sel(C_in[7]), 
        .S(S[31:28]) );
  carry_select_block_n4_24 csb_8 ( .A(A[35:32]), .B(B[35:32]), .C_sel(C_in[8]), 
        .S(S[35:32]) );
  carry_select_block_n4_23 csb_9 ( .A(A[39:36]), .B(B[39:36]), .C_sel(C_in[9]), 
        .S(S[39:36]) );
  carry_select_block_n4_22 csb_10 ( .A(A[43:40]), .B(B[43:40]), .C_sel(
        C_in[10]), .S(S[43:40]) );
  carry_select_block_n4_21 csb_11 ( .A(A[47:44]), .B(B[47:44]), .C_sel(
        C_in[11]), .S(S[47:44]) );
  carry_select_block_n4_20 csb_12 ( .A(A[51:48]), .B(B[51:48]), .C_sel(
        C_in[12]), .S(S[51:48]) );
  carry_select_block_n4_19 csb_13 ( .A(A[55:52]), .B(B[55:52]), .C_sel(
        C_in[13]), .S(S[55:52]) );
  carry_select_block_n4_18 csb_14 ( .A(A[59:56]), .B(B[59:56]), .C_sel(
        C_in[14]), .S(S[59:56]) );
  carry_select_block_n4_17 csb_15 ( .A(A[63:60]), .B(B[63:60]), .C_sel(
        C_in[15]), .S(S[63:60]) );
endmodule


module P4_ADDER_NBIT64_2 ( A, B, Cin, S, Cout, ovf );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Cin;
  output Cout, ovf;
  wire   n3, n4;
  wire   [63:0] xor_b;
  wire   [14:0] carry;

  XOR2_X1 U3 ( .A(xor_b[63]), .B(A[63]), .Z(n3) );
  my_xor_128 bc_xor_63 ( .A(B[63]), .B(Cin), .xor_out(xor_b[63]) );
  my_xor_127 bc_xor_62 ( .A(B[62]), .B(Cin), .xor_out(xor_b[62]) );
  my_xor_126 bc_xor_61 ( .A(B[61]), .B(Cin), .xor_out(xor_b[61]) );
  my_xor_125 bc_xor_60 ( .A(B[60]), .B(Cin), .xor_out(xor_b[60]) );
  my_xor_124 bc_xor_59 ( .A(B[59]), .B(Cin), .xor_out(xor_b[59]) );
  my_xor_123 bc_xor_58 ( .A(B[58]), .B(Cin), .xor_out(xor_b[58]) );
  my_xor_122 bc_xor_57 ( .A(B[57]), .B(Cin), .xor_out(xor_b[57]) );
  my_xor_121 bc_xor_56 ( .A(B[56]), .B(Cin), .xor_out(xor_b[56]) );
  my_xor_120 bc_xor_55 ( .A(B[55]), .B(Cin), .xor_out(xor_b[55]) );
  my_xor_119 bc_xor_54 ( .A(B[54]), .B(Cin), .xor_out(xor_b[54]) );
  my_xor_118 bc_xor_53 ( .A(B[53]), .B(Cin), .xor_out(xor_b[53]) );
  my_xor_117 bc_xor_52 ( .A(B[52]), .B(Cin), .xor_out(xor_b[52]) );
  my_xor_116 bc_xor_51 ( .A(B[51]), .B(Cin), .xor_out(xor_b[51]) );
  my_xor_115 bc_xor_50 ( .A(B[50]), .B(Cin), .xor_out(xor_b[50]) );
  my_xor_114 bc_xor_49 ( .A(B[49]), .B(Cin), .xor_out(xor_b[49]) );
  my_xor_113 bc_xor_48 ( .A(B[48]), .B(Cin), .xor_out(xor_b[48]) );
  my_xor_112 bc_xor_47 ( .A(B[47]), .B(Cin), .xor_out(xor_b[47]) );
  my_xor_111 bc_xor_46 ( .A(B[46]), .B(Cin), .xor_out(xor_b[46]) );
  my_xor_110 bc_xor_45 ( .A(B[45]), .B(Cin), .xor_out(xor_b[45]) );
  my_xor_109 bc_xor_44 ( .A(B[44]), .B(Cin), .xor_out(xor_b[44]) );
  my_xor_108 bc_xor_43 ( .A(B[43]), .B(Cin), .xor_out(xor_b[43]) );
  my_xor_107 bc_xor_42 ( .A(B[42]), .B(Cin), .xor_out(xor_b[42]) );
  my_xor_106 bc_xor_41 ( .A(B[41]), .B(Cin), .xor_out(xor_b[41]) );
  my_xor_105 bc_xor_40 ( .A(B[40]), .B(Cin), .xor_out(xor_b[40]) );
  my_xor_104 bc_xor_39 ( .A(B[39]), .B(Cin), .xor_out(xor_b[39]) );
  my_xor_103 bc_xor_38 ( .A(B[38]), .B(Cin), .xor_out(xor_b[38]) );
  my_xor_102 bc_xor_37 ( .A(B[37]), .B(Cin), .xor_out(xor_b[37]) );
  my_xor_101 bc_xor_36 ( .A(B[36]), .B(Cin), .xor_out(xor_b[36]) );
  my_xor_100 bc_xor_35 ( .A(B[35]), .B(Cin), .xor_out(xor_b[35]) );
  my_xor_99 bc_xor_34 ( .A(B[34]), .B(Cin), .xor_out(xor_b[34]) );
  my_xor_98 bc_xor_33 ( .A(B[33]), .B(Cin), .xor_out(xor_b[33]) );
  my_xor_97 bc_xor_32 ( .A(B[32]), .B(Cin), .xor_out(xor_b[32]) );
  my_xor_96 bc_xor_31 ( .A(B[31]), .B(Cin), .xor_out(xor_b[31]) );
  my_xor_95 bc_xor_30 ( .A(B[30]), .B(Cin), .xor_out(xor_b[30]) );
  my_xor_94 bc_xor_29 ( .A(B[29]), .B(Cin), .xor_out(xor_b[29]) );
  my_xor_93 bc_xor_28 ( .A(B[28]), .B(Cin), .xor_out(xor_b[28]) );
  my_xor_92 bc_xor_27 ( .A(B[27]), .B(Cin), .xor_out(xor_b[27]) );
  my_xor_91 bc_xor_26 ( .A(B[26]), .B(Cin), .xor_out(xor_b[26]) );
  my_xor_90 bc_xor_25 ( .A(B[25]), .B(Cin), .xor_out(xor_b[25]) );
  my_xor_89 bc_xor_24 ( .A(B[24]), .B(Cin), .xor_out(xor_b[24]) );
  my_xor_88 bc_xor_23 ( .A(B[23]), .B(Cin), .xor_out(xor_b[23]) );
  my_xor_87 bc_xor_22 ( .A(B[22]), .B(Cin), .xor_out(xor_b[22]) );
  my_xor_86 bc_xor_21 ( .A(B[21]), .B(Cin), .xor_out(xor_b[21]) );
  my_xor_85 bc_xor_20 ( .A(B[20]), .B(Cin), .xor_out(xor_b[20]) );
  my_xor_84 bc_xor_19 ( .A(B[19]), .B(Cin), .xor_out(xor_b[19]) );
  my_xor_83 bc_xor_18 ( .A(B[18]), .B(Cin), .xor_out(xor_b[18]) );
  my_xor_82 bc_xor_17 ( .A(B[17]), .B(Cin), .xor_out(xor_b[17]) );
  my_xor_81 bc_xor_16 ( .A(B[16]), .B(Cin), .xor_out(xor_b[16]) );
  my_xor_80 bc_xor_15 ( .A(B[15]), .B(Cin), .xor_out(xor_b[15]) );
  my_xor_79 bc_xor_14 ( .A(B[14]), .B(Cin), .xor_out(xor_b[14]) );
  my_xor_78 bc_xor_13 ( .A(B[13]), .B(Cin), .xor_out(xor_b[13]) );
  my_xor_77 bc_xor_12 ( .A(B[12]), .B(Cin), .xor_out(xor_b[12]) );
  my_xor_76 bc_xor_11 ( .A(B[11]), .B(Cin), .xor_out(xor_b[11]) );
  my_xor_75 bc_xor_10 ( .A(B[10]), .B(Cin), .xor_out(xor_b[10]) );
  my_xor_74 bc_xor_9 ( .A(B[9]), .B(Cin), .xor_out(xor_b[9]) );
  my_xor_73 bc_xor_8 ( .A(B[8]), .B(Cin), .xor_out(xor_b[8]) );
  my_xor_72 bc_xor_7 ( .A(B[7]), .B(Cin), .xor_out(xor_b[7]) );
  my_xor_71 bc_xor_6 ( .A(B[6]), .B(Cin), .xor_out(xor_b[6]) );
  my_xor_70 bc_xor_5 ( .A(B[5]), .B(Cin), .xor_out(xor_b[5]) );
  my_xor_69 bc_xor_4 ( .A(B[4]), .B(Cin), .xor_out(xor_b[4]) );
  my_xor_68 bc_xor_3 ( .A(B[3]), .B(Cin), .xor_out(xor_b[3]) );
  my_xor_67 bc_xor_2 ( .A(B[2]), .B(Cin), .xor_out(xor_b[2]) );
  my_xor_66 bc_xor_1 ( .A(B[1]), .B(Cin), .xor_out(xor_b[1]) );
  my_xor_65 bc_xor_0 ( .A(B[0]), .B(Cin), .xor_out(xor_b[0]) );
  CARRY_GENERATOR_NBIT64_NBIT_PER_BLOCK4_2 CG ( .A(A), .B(xor_b), .Cin(Cin), 
        .Co({Cout, carry}) );
  sum_generator_n_bit64_n_CSB16_2 SG ( .A(A), .B(xor_b), .C_in({carry, Cin}), 
        .S(S) );
  NOR2_X1 U1 ( .A1(n4), .A2(n3), .ZN(ovf) );
  XNOR2_X1 U2 ( .A(A[63]), .B(S[63]), .ZN(n4) );
endmodule


module my_xor_64 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_63 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_62 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_61 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_60 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_59 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_58 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_57 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_56 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_55 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_54 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_53 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_52 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_51 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_50 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_49 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_48 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_47 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_46 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_45 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_44 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_43 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_42 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_41 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_40 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_39 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_38 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_37 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_36 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_35 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_34 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_33 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_32 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_31 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_30 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_29 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_28 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_27 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_26 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_25 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_24 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_23 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_22 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_21 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_20 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_19 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_18 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_17 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_16 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_15 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_14 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_13 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_12 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_11 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_10 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_9 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_8 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_7 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_6 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_5 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_4 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_3 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_2 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module my_xor_1 ( A, B, xor_out );
  input A, B;
  output xor_out;


  XOR2_X1 U1 ( .A(B), .B(A), .Z(xor_out) );
endmodule


module pg_net_63 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_62 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_61 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_60 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_59 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_58 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_57 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_56 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_55 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_54 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_53 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_52 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_51 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_50 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_49 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_48 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_47 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_46 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_45 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_44 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_43 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_42 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_41 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_40 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_39 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_38 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_37 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_36 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_35 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_34 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_33 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_32 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_31 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_30 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_29 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_28 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_27 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_26 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_25 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_24 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_23 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_22 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_21 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_20 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_19 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_18 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_17 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_16 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_15 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_14 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_13 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_12 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_11 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_10 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_9 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_8 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_7 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_6 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_5 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_4 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_3 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_2 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module pg_net_1 ( a, b, p, g );
  input a, b;
  output p, g;


  XOR2_X1 U2 ( .A(b), .B(a), .Z(p) );
  AND2_X1 U1 ( .A1(b), .A2(a), .ZN(g) );
endmodule


module PG_BLOCK_63 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_62 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_61 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_60 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_59 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_58 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_57 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_56 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_55 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_54 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_53 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_52 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_51 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_50 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_49 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_48 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_47 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_46 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_45 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_44 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_43 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_42 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_41 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_40 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_39 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_38 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_37 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_36 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_35 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_34 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_33 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_17 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_32 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_31 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_30 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_29 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_28 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_27 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_26 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_25 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_24 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AOI21_X1 U1 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_23 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_22 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_21 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_20 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_19 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_18 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_16 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_17 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_16 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_15 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_14 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_13 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_12 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_11 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_15 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_10 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_9 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U2 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
  AND2_X1 U3 ( .A1(p2), .A2(p1), .ZN(PG_P) );
endmodule


module PG_BLOCK_8 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_7 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AND2_X1 U2 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_6 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AND2_X1 U2 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_5 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  AND2_X1 U1 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  INV_X1 U2 ( .A(n3), .ZN(PG_G) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_14 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_13 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_4 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AND2_X1 U2 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_3 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AND2_X1 U2 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_2 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AND2_X1 U2 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module PG_BLOCK_1 ( p2, g2, p1, g1, PG_P, PG_G );
  input p2, g2, p1, g1;
  output PG_P, PG_G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(PG_G) );
  AND2_X1 U2 ( .A1(p2), .A2(p1), .ZN(PG_P) );
  AOI21_X1 U3 ( .B1(g1), .B2(p2), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_12 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_11 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_10 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_9 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_8 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_7 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_6 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_5 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_4 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_3 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_2 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module G_BLOCK_1 ( p2, g2, g1, G );
  input p2, g2, g1;
  output G;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G) );
  AOI21_X1 U2 ( .B1(p2), .B2(g1), .A(g2), .ZN(n3) );
endmodule


module CARRY_GENERATOR_NBIT64_NBIT_PER_BLOCK4_1 ( A, B, Cin, Co );
  input [63:0] A;
  input [63:0] B;
  output [15:0] Co;
  input Cin;
  wire   \g_vector[5][63] , \g_vector[5][59] , \g_vector[5][55] ,
         \g_vector[5][51] , \g_vector[4][63] , \g_vector[4][59] ,
         \g_vector[4][47] , \g_vector[4][43] , \g_vector[4][31] ,
         \g_vector[4][27] , \g_vector[3][63] , \g_vector[3][55] ,
         \g_vector[3][47] , \g_vector[3][39] , \g_vector[3][31] ,
         \g_vector[3][23] , \g_vector[3][15] , \g_vector[2][63] ,
         \g_vector[2][59] , \g_vector[2][55] , \g_vector[2][51] ,
         \g_vector[2][47] , \g_vector[2][43] , \g_vector[2][39] ,
         \g_vector[2][35] , \g_vector[2][31] , \g_vector[2][27] ,
         \g_vector[2][23] , \g_vector[2][19] , \g_vector[2][15] ,
         \g_vector[2][11] , \g_vector[2][7] , \g_vector[1][63] ,
         \g_vector[1][61] , \g_vector[1][59] , \g_vector[1][57] ,
         \g_vector[1][55] , \g_vector[1][53] , \g_vector[1][51] ,
         \g_vector[1][49] , \g_vector[1][47] , \g_vector[1][45] ,
         \g_vector[1][43] , \g_vector[1][41] , \g_vector[1][39] ,
         \g_vector[1][37] , \g_vector[1][35] , \g_vector[1][33] ,
         \g_vector[1][31] , \g_vector[1][29] , \g_vector[1][27] ,
         \g_vector[1][25] , \g_vector[1][23] , \g_vector[1][21] ,
         \g_vector[1][19] , \g_vector[1][17] , \g_vector[1][15] ,
         \g_vector[1][13] , \g_vector[1][11] , \g_vector[1][9] ,
         \g_vector[1][7] , \g_vector[1][5] , \g_vector[1][3] ,
         \g_vector[1][1] , \g_vector[0][63] , \g_vector[0][62] ,
         \g_vector[0][61] , \g_vector[0][60] , \g_vector[0][59] ,
         \g_vector[0][58] , \g_vector[0][57] , \g_vector[0][56] ,
         \g_vector[0][55] , \g_vector[0][54] , \g_vector[0][53] ,
         \g_vector[0][52] , \g_vector[0][51] , \g_vector[0][50] ,
         \g_vector[0][49] , \g_vector[0][48] , \g_vector[0][47] ,
         \g_vector[0][46] , \g_vector[0][45] , \g_vector[0][44] ,
         \g_vector[0][43] , \g_vector[0][42] , \g_vector[0][41] ,
         \g_vector[0][40] , \g_vector[0][39] , \g_vector[0][38] ,
         \g_vector[0][37] , \g_vector[0][36] , \g_vector[0][35] ,
         \g_vector[0][34] , \g_vector[0][33] , \g_vector[0][32] ,
         \g_vector[0][31] , \g_vector[0][30] , \g_vector[0][29] ,
         \g_vector[0][28] , \g_vector[0][27] , \g_vector[0][26] ,
         \g_vector[0][25] , \g_vector[0][24] , \g_vector[0][23] ,
         \g_vector[0][22] , \g_vector[0][21] , \g_vector[0][20] ,
         \g_vector[0][19] , \g_vector[0][18] , \g_vector[0][17] ,
         \g_vector[0][16] , \g_vector[0][15] , \g_vector[0][14] ,
         \g_vector[0][13] , \g_vector[0][12] , \g_vector[0][11] ,
         \g_vector[0][10] , \g_vector[0][9] , \g_vector[0][8] ,
         \g_vector[0][7] , \g_vector[0][6] , \g_vector[0][5] ,
         \g_vector[0][4] , \g_vector[0][3] , \g_vector[0][2] ,
         \g_vector[0][1] , \g_vector[0][0] , \p_vector[5][63] ,
         \p_vector[5][59] , \p_vector[5][55] , \p_vector[5][51] ,
         \p_vector[4][63] , \p_vector[4][59] , \p_vector[4][47] ,
         \p_vector[4][43] , \p_vector[4][31] , \p_vector[4][27] ,
         \p_vector[3][63] , \p_vector[3][55] , \p_vector[3][47] ,
         \p_vector[3][39] , \p_vector[3][31] , \p_vector[3][23] ,
         \p_vector[3][15] , \p_vector[2][63] , \p_vector[2][59] ,
         \p_vector[2][55] , \p_vector[2][51] , \p_vector[2][47] ,
         \p_vector[2][43] , \p_vector[2][39] , \p_vector[2][35] ,
         \p_vector[2][31] , \p_vector[2][27] , \p_vector[2][23] ,
         \p_vector[2][19] , \p_vector[2][15] , \p_vector[2][11] ,
         \p_vector[2][7] , \p_vector[1][63] , \p_vector[1][61] ,
         \p_vector[1][59] , \p_vector[1][57] , \p_vector[1][55] ,
         \p_vector[1][53] , \p_vector[1][51] , \p_vector[1][49] ,
         \p_vector[1][47] , \p_vector[1][45] , \p_vector[1][43] ,
         \p_vector[1][41] , \p_vector[1][39] , \p_vector[1][37] ,
         \p_vector[1][35] , \p_vector[1][33] , \p_vector[1][31] ,
         \p_vector[1][29] , \p_vector[1][27] , \p_vector[1][25] ,
         \p_vector[1][23] , \p_vector[1][21] , \p_vector[1][19] ,
         \p_vector[1][17] , \p_vector[1][15] , \p_vector[1][13] ,
         \p_vector[1][11] , \p_vector[1][9] , \p_vector[1][7] ,
         \p_vector[1][5] , \p_vector[1][3] , \p_vector[0][63] ,
         \p_vector[0][62] , \p_vector[0][61] , \p_vector[0][60] ,
         \p_vector[0][59] , \p_vector[0][58] , \p_vector[0][57] ,
         \p_vector[0][56] , \p_vector[0][55] , \p_vector[0][54] ,
         \p_vector[0][53] , \p_vector[0][52] , \p_vector[0][51] ,
         \p_vector[0][50] , \p_vector[0][49] , \p_vector[0][48] ,
         \p_vector[0][47] , \p_vector[0][46] , \p_vector[0][45] ,
         \p_vector[0][44] , \p_vector[0][43] , \p_vector[0][42] ,
         \p_vector[0][41] , \p_vector[0][40] , \p_vector[0][39] ,
         \p_vector[0][38] , \p_vector[0][37] , \p_vector[0][36] ,
         \p_vector[0][35] , \p_vector[0][34] , \p_vector[0][33] ,
         \p_vector[0][32] , \p_vector[0][31] , \p_vector[0][30] ,
         \p_vector[0][29] , \p_vector[0][28] , \p_vector[0][27] ,
         \p_vector[0][26] , \p_vector[0][25] , \p_vector[0][24] ,
         \p_vector[0][23] , \p_vector[0][22] , \p_vector[0][21] ,
         \p_vector[0][20] , \p_vector[0][19] , \p_vector[0][18] ,
         \p_vector[0][17] , \p_vector[0][16] , \p_vector[0][15] ,
         \p_vector[0][14] , \p_vector[0][13] , \p_vector[0][12] ,
         \p_vector[0][11] , \p_vector[0][10] , \p_vector[0][9] ,
         \p_vector[0][8] , \p_vector[0][7] , \p_vector[0][6] ,
         \p_vector[0][5] , \p_vector[0][4] , \p_vector[0][3] ,
         \p_vector[0][2] , \p_vector[0][1] , n1, n2, n4;

  pg_net_63 pg_network_63 ( .a(A[63]), .b(B[63]), .p(\p_vector[0][63] ), .g(
        \g_vector[0][63] ) );
  pg_net_62 pg_network_62 ( .a(A[62]), .b(B[62]), .p(\p_vector[0][62] ), .g(
        \g_vector[0][62] ) );
  pg_net_61 pg_network_61 ( .a(A[61]), .b(B[61]), .p(\p_vector[0][61] ), .g(
        \g_vector[0][61] ) );
  pg_net_60 pg_network_60 ( .a(A[60]), .b(B[60]), .p(\p_vector[0][60] ), .g(
        \g_vector[0][60] ) );
  pg_net_59 pg_network_59 ( .a(A[59]), .b(B[59]), .p(\p_vector[0][59] ), .g(
        \g_vector[0][59] ) );
  pg_net_58 pg_network_58 ( .a(A[58]), .b(B[58]), .p(\p_vector[0][58] ), .g(
        \g_vector[0][58] ) );
  pg_net_57 pg_network_57 ( .a(A[57]), .b(B[57]), .p(\p_vector[0][57] ), .g(
        \g_vector[0][57] ) );
  pg_net_56 pg_network_56 ( .a(A[56]), .b(B[56]), .p(\p_vector[0][56] ), .g(
        \g_vector[0][56] ) );
  pg_net_55 pg_network_55 ( .a(A[55]), .b(B[55]), .p(\p_vector[0][55] ), .g(
        \g_vector[0][55] ) );
  pg_net_54 pg_network_54 ( .a(A[54]), .b(B[54]), .p(\p_vector[0][54] ), .g(
        \g_vector[0][54] ) );
  pg_net_53 pg_network_53 ( .a(A[53]), .b(B[53]), .p(\p_vector[0][53] ), .g(
        \g_vector[0][53] ) );
  pg_net_52 pg_network_52 ( .a(A[52]), .b(B[52]), .p(\p_vector[0][52] ), .g(
        \g_vector[0][52] ) );
  pg_net_51 pg_network_51 ( .a(A[51]), .b(B[51]), .p(\p_vector[0][51] ), .g(
        \g_vector[0][51] ) );
  pg_net_50 pg_network_50 ( .a(A[50]), .b(B[50]), .p(\p_vector[0][50] ), .g(
        \g_vector[0][50] ) );
  pg_net_49 pg_network_49 ( .a(A[49]), .b(B[49]), .p(\p_vector[0][49] ), .g(
        \g_vector[0][49] ) );
  pg_net_48 pg_network_48 ( .a(A[48]), .b(B[48]), .p(\p_vector[0][48] ), .g(
        \g_vector[0][48] ) );
  pg_net_47 pg_network_47 ( .a(A[47]), .b(B[47]), .p(\p_vector[0][47] ), .g(
        \g_vector[0][47] ) );
  pg_net_46 pg_network_46 ( .a(A[46]), .b(B[46]), .p(\p_vector[0][46] ), .g(
        \g_vector[0][46] ) );
  pg_net_45 pg_network_45 ( .a(A[45]), .b(B[45]), .p(\p_vector[0][45] ), .g(
        \g_vector[0][45] ) );
  pg_net_44 pg_network_44 ( .a(A[44]), .b(B[44]), .p(\p_vector[0][44] ), .g(
        \g_vector[0][44] ) );
  pg_net_43 pg_network_43 ( .a(A[43]), .b(B[43]), .p(\p_vector[0][43] ), .g(
        \g_vector[0][43] ) );
  pg_net_42 pg_network_42 ( .a(A[42]), .b(B[42]), .p(\p_vector[0][42] ), .g(
        \g_vector[0][42] ) );
  pg_net_41 pg_network_41 ( .a(A[41]), .b(B[41]), .p(\p_vector[0][41] ), .g(
        \g_vector[0][41] ) );
  pg_net_40 pg_network_40 ( .a(A[40]), .b(B[40]), .p(\p_vector[0][40] ), .g(
        \g_vector[0][40] ) );
  pg_net_39 pg_network_39 ( .a(A[39]), .b(B[39]), .p(\p_vector[0][39] ), .g(
        \g_vector[0][39] ) );
  pg_net_38 pg_network_38 ( .a(A[38]), .b(B[38]), .p(\p_vector[0][38] ), .g(
        \g_vector[0][38] ) );
  pg_net_37 pg_network_37 ( .a(A[37]), .b(B[37]), .p(\p_vector[0][37] ), .g(
        \g_vector[0][37] ) );
  pg_net_36 pg_network_36 ( .a(A[36]), .b(B[36]), .p(\p_vector[0][36] ), .g(
        \g_vector[0][36] ) );
  pg_net_35 pg_network_35 ( .a(A[35]), .b(B[35]), .p(\p_vector[0][35] ), .g(
        \g_vector[0][35] ) );
  pg_net_34 pg_network_34 ( .a(A[34]), .b(B[34]), .p(\p_vector[0][34] ), .g(
        \g_vector[0][34] ) );
  pg_net_33 pg_network_33 ( .a(A[33]), .b(B[33]), .p(\p_vector[0][33] ), .g(
        \g_vector[0][33] ) );
  pg_net_32 pg_network_32 ( .a(A[32]), .b(B[32]), .p(\p_vector[0][32] ), .g(
        \g_vector[0][32] ) );
  pg_net_31 pg_network_31 ( .a(A[31]), .b(B[31]), .p(\p_vector[0][31] ), .g(
        \g_vector[0][31] ) );
  pg_net_30 pg_network_30 ( .a(A[30]), .b(B[30]), .p(\p_vector[0][30] ), .g(
        \g_vector[0][30] ) );
  pg_net_29 pg_network_29 ( .a(A[29]), .b(B[29]), .p(\p_vector[0][29] ), .g(
        \g_vector[0][29] ) );
  pg_net_28 pg_network_28 ( .a(A[28]), .b(B[28]), .p(\p_vector[0][28] ), .g(
        \g_vector[0][28] ) );
  pg_net_27 pg_network_27 ( .a(A[27]), .b(B[27]), .p(\p_vector[0][27] ), .g(
        \g_vector[0][27] ) );
  pg_net_26 pg_network_26 ( .a(A[26]), .b(B[26]), .p(\p_vector[0][26] ), .g(
        \g_vector[0][26] ) );
  pg_net_25 pg_network_25 ( .a(A[25]), .b(B[25]), .p(\p_vector[0][25] ), .g(
        \g_vector[0][25] ) );
  pg_net_24 pg_network_24 ( .a(A[24]), .b(B[24]), .p(\p_vector[0][24] ), .g(
        \g_vector[0][24] ) );
  pg_net_23 pg_network_23 ( .a(A[23]), .b(B[23]), .p(\p_vector[0][23] ), .g(
        \g_vector[0][23] ) );
  pg_net_22 pg_network_22 ( .a(A[22]), .b(B[22]), .p(\p_vector[0][22] ), .g(
        \g_vector[0][22] ) );
  pg_net_21 pg_network_21 ( .a(A[21]), .b(B[21]), .p(\p_vector[0][21] ), .g(
        \g_vector[0][21] ) );
  pg_net_20 pg_network_20 ( .a(A[20]), .b(B[20]), .p(\p_vector[0][20] ), .g(
        \g_vector[0][20] ) );
  pg_net_19 pg_network_19 ( .a(A[19]), .b(B[19]), .p(\p_vector[0][19] ), .g(
        \g_vector[0][19] ) );
  pg_net_18 pg_network_18 ( .a(A[18]), .b(B[18]), .p(\p_vector[0][18] ), .g(
        \g_vector[0][18] ) );
  pg_net_17 pg_network_17 ( .a(A[17]), .b(B[17]), .p(\p_vector[0][17] ), .g(
        \g_vector[0][17] ) );
  pg_net_16 pg_network_16 ( .a(A[16]), .b(B[16]), .p(\p_vector[0][16] ), .g(
        \g_vector[0][16] ) );
  pg_net_15 pg_network_15 ( .a(A[15]), .b(B[15]), .p(\p_vector[0][15] ), .g(
        \g_vector[0][15] ) );
  pg_net_14 pg_network_14 ( .a(A[14]), .b(B[14]), .p(\p_vector[0][14] ), .g(
        \g_vector[0][14] ) );
  pg_net_13 pg_network_13 ( .a(A[13]), .b(B[13]), .p(\p_vector[0][13] ), .g(
        \g_vector[0][13] ) );
  pg_net_12 pg_network_12 ( .a(A[12]), .b(B[12]), .p(\p_vector[0][12] ), .g(
        \g_vector[0][12] ) );
  pg_net_11 pg_network_11 ( .a(A[11]), .b(B[11]), .p(\p_vector[0][11] ), .g(
        \g_vector[0][11] ) );
  pg_net_10 pg_network_10 ( .a(A[10]), .b(B[10]), .p(\p_vector[0][10] ), .g(
        \g_vector[0][10] ) );
  pg_net_9 pg_network_9 ( .a(A[9]), .b(B[9]), .p(\p_vector[0][9] ), .g(
        \g_vector[0][9] ) );
  pg_net_8 pg_network_8 ( .a(A[8]), .b(B[8]), .p(\p_vector[0][8] ), .g(
        \g_vector[0][8] ) );
  pg_net_7 pg_network_7 ( .a(A[7]), .b(B[7]), .p(\p_vector[0][7] ), .g(
        \g_vector[0][7] ) );
  pg_net_6 pg_network_6 ( .a(A[6]), .b(B[6]), .p(\p_vector[0][6] ), .g(
        \g_vector[0][6] ) );
  pg_net_5 pg_network_5 ( .a(A[5]), .b(B[5]), .p(\p_vector[0][5] ), .g(
        \g_vector[0][5] ) );
  pg_net_4 pg_network_4 ( .a(A[4]), .b(B[4]), .p(\p_vector[0][4] ), .g(
        \g_vector[0][4] ) );
  pg_net_3 pg_network_3 ( .a(A[3]), .b(B[3]), .p(\p_vector[0][3] ), .g(
        \g_vector[0][3] ) );
  pg_net_2 pg_network_2 ( .a(A[2]), .b(B[2]), .p(\p_vector[0][2] ), .g(
        \g_vector[0][2] ) );
  pg_net_1 pg_network_1 ( .a(A[1]), .b(B[1]), .p(\p_vector[0][1] ), .g(
        \g_vector[0][1] ) );
  PG_BLOCK_63 std_PG_1_63 ( .p2(\p_vector[0][63] ), .g2(\g_vector[0][63] ), 
        .p1(\p_vector[0][62] ), .g1(\g_vector[0][62] ), .PG_P(
        \p_vector[1][63] ), .PG_G(\g_vector[1][63] ) );
  PG_BLOCK_62 std_PG_1_61 ( .p2(\p_vector[0][61] ), .g2(\g_vector[0][61] ), 
        .p1(\p_vector[0][60] ), .g1(\g_vector[0][60] ), .PG_P(
        \p_vector[1][61] ), .PG_G(\g_vector[1][61] ) );
  PG_BLOCK_61 std_PG_1_59 ( .p2(\p_vector[0][59] ), .g2(\g_vector[0][59] ), 
        .p1(\p_vector[0][58] ), .g1(\g_vector[0][58] ), .PG_P(
        \p_vector[1][59] ), .PG_G(\g_vector[1][59] ) );
  PG_BLOCK_60 std_PG_1_57 ( .p2(\p_vector[0][57] ), .g2(\g_vector[0][57] ), 
        .p1(\p_vector[0][56] ), .g1(\g_vector[0][56] ), .PG_P(
        \p_vector[1][57] ), .PG_G(\g_vector[1][57] ) );
  PG_BLOCK_59 std_PG_1_55 ( .p2(\p_vector[0][55] ), .g2(\g_vector[0][55] ), 
        .p1(\p_vector[0][54] ), .g1(\g_vector[0][54] ), .PG_P(
        \p_vector[1][55] ), .PG_G(\g_vector[1][55] ) );
  PG_BLOCK_58 std_PG_1_53 ( .p2(\p_vector[0][53] ), .g2(\g_vector[0][53] ), 
        .p1(\p_vector[0][52] ), .g1(\g_vector[0][52] ), .PG_P(
        \p_vector[1][53] ), .PG_G(\g_vector[1][53] ) );
  PG_BLOCK_57 std_PG_1_51 ( .p2(\p_vector[0][51] ), .g2(\g_vector[0][51] ), 
        .p1(\p_vector[0][50] ), .g1(\g_vector[0][50] ), .PG_P(
        \p_vector[1][51] ), .PG_G(\g_vector[1][51] ) );
  PG_BLOCK_56 std_PG_1_49 ( .p2(\p_vector[0][49] ), .g2(\g_vector[0][49] ), 
        .p1(\p_vector[0][48] ), .g1(\g_vector[0][48] ), .PG_P(
        \p_vector[1][49] ), .PG_G(\g_vector[1][49] ) );
  PG_BLOCK_55 std_PG_1_47 ( .p2(\p_vector[0][47] ), .g2(\g_vector[0][47] ), 
        .p1(\p_vector[0][46] ), .g1(\g_vector[0][46] ), .PG_P(
        \p_vector[1][47] ), .PG_G(\g_vector[1][47] ) );
  PG_BLOCK_54 std_PG_1_45 ( .p2(\p_vector[0][45] ), .g2(\g_vector[0][45] ), 
        .p1(\p_vector[0][44] ), .g1(\g_vector[0][44] ), .PG_P(
        \p_vector[1][45] ), .PG_G(\g_vector[1][45] ) );
  PG_BLOCK_53 std_PG_1_43 ( .p2(\p_vector[0][43] ), .g2(\g_vector[0][43] ), 
        .p1(\p_vector[0][42] ), .g1(\g_vector[0][42] ), .PG_P(
        \p_vector[1][43] ), .PG_G(\g_vector[1][43] ) );
  PG_BLOCK_52 std_PG_1_41 ( .p2(\p_vector[0][41] ), .g2(\g_vector[0][41] ), 
        .p1(\p_vector[0][40] ), .g1(\g_vector[0][40] ), .PG_P(
        \p_vector[1][41] ), .PG_G(\g_vector[1][41] ) );
  PG_BLOCK_51 std_PG_1_39 ( .p2(\p_vector[0][39] ), .g2(\g_vector[0][39] ), 
        .p1(\p_vector[0][38] ), .g1(\g_vector[0][38] ), .PG_P(
        \p_vector[1][39] ), .PG_G(\g_vector[1][39] ) );
  PG_BLOCK_50 std_PG_1_37 ( .p2(\p_vector[0][37] ), .g2(\g_vector[0][37] ), 
        .p1(\p_vector[0][36] ), .g1(\g_vector[0][36] ), .PG_P(
        \p_vector[1][37] ), .PG_G(\g_vector[1][37] ) );
  PG_BLOCK_49 std_PG_1_35 ( .p2(\p_vector[0][35] ), .g2(\g_vector[0][35] ), 
        .p1(\p_vector[0][34] ), .g1(\g_vector[0][34] ), .PG_P(
        \p_vector[1][35] ), .PG_G(\g_vector[1][35] ) );
  PG_BLOCK_48 std_PG_1_33 ( .p2(\p_vector[0][33] ), .g2(\g_vector[0][33] ), 
        .p1(\p_vector[0][32] ), .g1(\g_vector[0][32] ), .PG_P(
        \p_vector[1][33] ), .PG_G(\g_vector[1][33] ) );
  PG_BLOCK_47 std_PG_1_31 ( .p2(\p_vector[0][31] ), .g2(\g_vector[0][31] ), 
        .p1(\p_vector[0][30] ), .g1(\g_vector[0][30] ), .PG_P(
        \p_vector[1][31] ), .PG_G(\g_vector[1][31] ) );
  PG_BLOCK_46 std_PG_1_29 ( .p2(\p_vector[0][29] ), .g2(\g_vector[0][29] ), 
        .p1(\p_vector[0][28] ), .g1(\g_vector[0][28] ), .PG_P(
        \p_vector[1][29] ), .PG_G(\g_vector[1][29] ) );
  PG_BLOCK_45 std_PG_1_27 ( .p2(\p_vector[0][27] ), .g2(\g_vector[0][27] ), 
        .p1(\p_vector[0][26] ), .g1(\g_vector[0][26] ), .PG_P(
        \p_vector[1][27] ), .PG_G(\g_vector[1][27] ) );
  PG_BLOCK_44 std_PG_1_25 ( .p2(\p_vector[0][25] ), .g2(\g_vector[0][25] ), 
        .p1(\p_vector[0][24] ), .g1(\g_vector[0][24] ), .PG_P(
        \p_vector[1][25] ), .PG_G(\g_vector[1][25] ) );
  PG_BLOCK_43 std_PG_1_23 ( .p2(\p_vector[0][23] ), .g2(\g_vector[0][23] ), 
        .p1(\p_vector[0][22] ), .g1(\g_vector[0][22] ), .PG_P(
        \p_vector[1][23] ), .PG_G(\g_vector[1][23] ) );
  PG_BLOCK_42 std_PG_1_21 ( .p2(\p_vector[0][21] ), .g2(\g_vector[0][21] ), 
        .p1(\p_vector[0][20] ), .g1(\g_vector[0][20] ), .PG_P(
        \p_vector[1][21] ), .PG_G(\g_vector[1][21] ) );
  PG_BLOCK_41 std_PG_1_19 ( .p2(\p_vector[0][19] ), .g2(\g_vector[0][19] ), 
        .p1(\p_vector[0][18] ), .g1(\g_vector[0][18] ), .PG_P(
        \p_vector[1][19] ), .PG_G(\g_vector[1][19] ) );
  PG_BLOCK_40 std_PG_1_17 ( .p2(\p_vector[0][17] ), .g2(\g_vector[0][17] ), 
        .p1(\p_vector[0][16] ), .g1(\g_vector[0][16] ), .PG_P(
        \p_vector[1][17] ), .PG_G(\g_vector[1][17] ) );
  PG_BLOCK_39 std_PG_1_15 ( .p2(\p_vector[0][15] ), .g2(\g_vector[0][15] ), 
        .p1(\p_vector[0][14] ), .g1(\g_vector[0][14] ), .PG_P(
        \p_vector[1][15] ), .PG_G(\g_vector[1][15] ) );
  PG_BLOCK_38 std_PG_1_13 ( .p2(\p_vector[0][13] ), .g2(\g_vector[0][13] ), 
        .p1(\p_vector[0][12] ), .g1(\g_vector[0][12] ), .PG_P(
        \p_vector[1][13] ), .PG_G(\g_vector[1][13] ) );
  PG_BLOCK_37 std_PG_1_11 ( .p2(\p_vector[0][11] ), .g2(\g_vector[0][11] ), 
        .p1(\p_vector[0][10] ), .g1(\g_vector[0][10] ), .PG_P(
        \p_vector[1][11] ), .PG_G(\g_vector[1][11] ) );
  PG_BLOCK_36 std_PG_1_9 ( .p2(\p_vector[0][9] ), .g2(\g_vector[0][9] ), .p1(
        \p_vector[0][8] ), .g1(\g_vector[0][8] ), .PG_P(\p_vector[1][9] ), 
        .PG_G(\g_vector[1][9] ) );
  PG_BLOCK_35 std_PG_1_7 ( .p2(\p_vector[0][7] ), .g2(\g_vector[0][7] ), .p1(
        \p_vector[0][6] ), .g1(\g_vector[0][6] ), .PG_P(\p_vector[1][7] ), 
        .PG_G(\g_vector[1][7] ) );
  PG_BLOCK_34 std_PG_1_5 ( .p2(\p_vector[0][5] ), .g2(\g_vector[0][5] ), .p1(
        \p_vector[0][4] ), .g1(\g_vector[0][4] ), .PG_P(\p_vector[1][5] ), 
        .PG_G(\g_vector[1][5] ) );
  PG_BLOCK_33 std_PG_1_3 ( .p2(\p_vector[0][3] ), .g2(\g_vector[0][3] ), .p1(
        \p_vector[0][2] ), .g1(\g_vector[0][2] ), .PG_P(\p_vector[1][3] ), 
        .PG_G(\g_vector[1][3] ) );
  G_BLOCK_17 std_G_1_1 ( .p2(\p_vector[0][1] ), .g2(\g_vector[0][1] ), .g1(
        \g_vector[0][0] ), .G(\g_vector[1][1] ) );
  PG_BLOCK_32 std_PG_2_63 ( .p2(\p_vector[1][63] ), .g2(\g_vector[1][63] ), 
        .p1(\p_vector[1][61] ), .g1(\g_vector[1][61] ), .PG_P(
        \p_vector[2][63] ), .PG_G(\g_vector[2][63] ) );
  PG_BLOCK_31 std_PG_2_59 ( .p2(\p_vector[1][59] ), .g2(\g_vector[1][59] ), 
        .p1(\p_vector[1][57] ), .g1(\g_vector[1][57] ), .PG_P(
        \p_vector[2][59] ), .PG_G(\g_vector[2][59] ) );
  PG_BLOCK_30 std_PG_2_55 ( .p2(\p_vector[1][55] ), .g2(\g_vector[1][55] ), 
        .p1(\p_vector[1][53] ), .g1(\g_vector[1][53] ), .PG_P(
        \p_vector[2][55] ), .PG_G(\g_vector[2][55] ) );
  PG_BLOCK_29 std_PG_2_51 ( .p2(\p_vector[1][51] ), .g2(\g_vector[1][51] ), 
        .p1(\p_vector[1][49] ), .g1(\g_vector[1][49] ), .PG_P(
        \p_vector[2][51] ), .PG_G(\g_vector[2][51] ) );
  PG_BLOCK_28 std_PG_2_47 ( .p2(\p_vector[1][47] ), .g2(\g_vector[1][47] ), 
        .p1(\p_vector[1][45] ), .g1(\g_vector[1][45] ), .PG_P(
        \p_vector[2][47] ), .PG_G(\g_vector[2][47] ) );
  PG_BLOCK_27 std_PG_2_43 ( .p2(\p_vector[1][43] ), .g2(\g_vector[1][43] ), 
        .p1(\p_vector[1][41] ), .g1(\g_vector[1][41] ), .PG_P(
        \p_vector[2][43] ), .PG_G(\g_vector[2][43] ) );
  PG_BLOCK_26 std_PG_2_39 ( .p2(\p_vector[1][39] ), .g2(\g_vector[1][39] ), 
        .p1(\p_vector[1][37] ), .g1(\g_vector[1][37] ), .PG_P(
        \p_vector[2][39] ), .PG_G(\g_vector[2][39] ) );
  PG_BLOCK_25 std_PG_2_35 ( .p2(\p_vector[1][35] ), .g2(\g_vector[1][35] ), 
        .p1(\p_vector[1][33] ), .g1(\g_vector[1][33] ), .PG_P(
        \p_vector[2][35] ), .PG_G(\g_vector[2][35] ) );
  PG_BLOCK_24 std_PG_2_31 ( .p2(\p_vector[1][31] ), .g2(\g_vector[1][31] ), 
        .p1(\p_vector[1][29] ), .g1(\g_vector[1][29] ), .PG_P(
        \p_vector[2][31] ), .PG_G(\g_vector[2][31] ) );
  PG_BLOCK_23 std_PG_2_27 ( .p2(\p_vector[1][27] ), .g2(\g_vector[1][27] ), 
        .p1(\p_vector[1][25] ), .g1(\g_vector[1][25] ), .PG_P(
        \p_vector[2][27] ), .PG_G(\g_vector[2][27] ) );
  PG_BLOCK_22 std_PG_2_23 ( .p2(\p_vector[1][23] ), .g2(\g_vector[1][23] ), 
        .p1(\p_vector[1][21] ), .g1(\g_vector[1][21] ), .PG_P(
        \p_vector[2][23] ), .PG_G(\g_vector[2][23] ) );
  PG_BLOCK_21 std_PG_2_19 ( .p2(\p_vector[1][19] ), .g2(\g_vector[1][19] ), 
        .p1(\p_vector[1][17] ), .g1(\g_vector[1][17] ), .PG_P(
        \p_vector[2][19] ), .PG_G(\g_vector[2][19] ) );
  PG_BLOCK_20 std_PG_2_15 ( .p2(\p_vector[1][15] ), .g2(\g_vector[1][15] ), 
        .p1(\p_vector[1][13] ), .g1(\g_vector[1][13] ), .PG_P(
        \p_vector[2][15] ), .PG_G(\g_vector[2][15] ) );
  PG_BLOCK_19 std_PG_2_11 ( .p2(\p_vector[1][11] ), .g2(\g_vector[1][11] ), 
        .p1(\p_vector[1][9] ), .g1(\g_vector[1][9] ), .PG_P(\p_vector[2][11] ), 
        .PG_G(\g_vector[2][11] ) );
  PG_BLOCK_18 std_PG_2_7 ( .p2(\p_vector[1][7] ), .g2(\g_vector[1][7] ), .p1(
        \p_vector[1][5] ), .g1(\g_vector[1][5] ), .PG_P(\p_vector[2][7] ), 
        .PG_G(\g_vector[2][7] ) );
  G_BLOCK_16 std_G_2_3 ( .p2(\p_vector[1][3] ), .g2(\g_vector[1][3] ), .g1(
        \g_vector[1][1] ), .G(Co[0]) );
  PG_BLOCK_17 std_PG_3_63 ( .p2(\p_vector[2][63] ), .g2(\g_vector[2][63] ), 
        .p1(\p_vector[2][59] ), .g1(\g_vector[2][59] ), .PG_P(
        \p_vector[3][63] ), .PG_G(\g_vector[3][63] ) );
  PG_BLOCK_16 std_PG_3_55 ( .p2(\p_vector[2][55] ), .g2(\g_vector[2][55] ), 
        .p1(\p_vector[2][51] ), .g1(\g_vector[2][51] ), .PG_P(
        \p_vector[3][55] ), .PG_G(\g_vector[3][55] ) );
  PG_BLOCK_15 std_PG_3_47 ( .p2(\p_vector[2][47] ), .g2(\g_vector[2][47] ), 
        .p1(\p_vector[2][43] ), .g1(\g_vector[2][43] ), .PG_P(
        \p_vector[3][47] ), .PG_G(\g_vector[3][47] ) );
  PG_BLOCK_14 std_PG_3_39 ( .p2(\p_vector[2][39] ), .g2(\g_vector[2][39] ), 
        .p1(\p_vector[2][35] ), .g1(\g_vector[2][35] ), .PG_P(
        \p_vector[3][39] ), .PG_G(\g_vector[3][39] ) );
  PG_BLOCK_13 std_PG_3_31 ( .p2(\p_vector[2][31] ), .g2(\g_vector[2][31] ), 
        .p1(\p_vector[2][27] ), .g1(\g_vector[2][27] ), .PG_P(
        \p_vector[3][31] ), .PG_G(\g_vector[3][31] ) );
  PG_BLOCK_12 std_PG_3_23 ( .p2(\p_vector[2][23] ), .g2(\g_vector[2][23] ), 
        .p1(\p_vector[2][19] ), .g1(\g_vector[2][19] ), .PG_P(
        \p_vector[3][23] ), .PG_G(\g_vector[3][23] ) );
  PG_BLOCK_11 std_PG_3_15 ( .p2(\p_vector[2][15] ), .g2(\g_vector[2][15] ), 
        .p1(\p_vector[2][11] ), .g1(\g_vector[2][11] ), .PG_P(
        \p_vector[3][15] ), .PG_G(\g_vector[3][15] ) );
  G_BLOCK_15 std_G_3_7 ( .p2(\p_vector[2][7] ), .g2(\g_vector[2][7] ), .g1(
        Co[0]), .G(Co[1]) );
  PG_BLOCK_10 std_PG_4_63 ( .p2(\p_vector[3][63] ), .g2(\g_vector[3][63] ), 
        .p1(\p_vector[3][55] ), .g1(\g_vector[3][55] ), .PG_P(
        \p_vector[4][63] ), .PG_G(\g_vector[4][63] ) );
  PG_BLOCK_9 add_PG_4_63_1 ( .p2(\p_vector[2][59] ), .g2(\g_vector[2][59] ), 
        .p1(\p_vector[3][55] ), .g1(\g_vector[3][55] ), .PG_P(
        \p_vector[4][59] ), .PG_G(\g_vector[4][59] ) );
  PG_BLOCK_8 std_PG_4_47 ( .p2(\p_vector[3][47] ), .g2(\g_vector[3][47] ), 
        .p1(\p_vector[3][39] ), .g1(\g_vector[3][39] ), .PG_P(
        \p_vector[4][47] ), .PG_G(\g_vector[4][47] ) );
  PG_BLOCK_7 add_PG_4_47_1 ( .p2(\p_vector[2][43] ), .g2(\g_vector[2][43] ), 
        .p1(\p_vector[3][39] ), .g1(\g_vector[3][39] ), .PG_P(
        \p_vector[4][43] ), .PG_G(\g_vector[4][43] ) );
  PG_BLOCK_6 std_PG_4_31 ( .p2(\p_vector[3][31] ), .g2(\g_vector[3][31] ), 
        .p1(\p_vector[3][23] ), .g1(\g_vector[3][23] ), .PG_P(
        \p_vector[4][31] ), .PG_G(\g_vector[4][31] ) );
  PG_BLOCK_5 add_PG_4_31_1 ( .p2(\p_vector[2][27] ), .g2(\g_vector[2][27] ), 
        .p1(\p_vector[3][23] ), .g1(\g_vector[3][23] ), .PG_P(
        \p_vector[4][27] ), .PG_G(\g_vector[4][27] ) );
  G_BLOCK_14 std_G_4_15 ( .p2(\p_vector[3][15] ), .g2(\g_vector[3][15] ), .g1(
        Co[1]), .G(Co[3]) );
  G_BLOCK_13 add_G_4_15_1 ( .p2(\p_vector[2][11] ), .g2(\g_vector[2][11] ), 
        .g1(Co[1]), .G(Co[2]) );
  PG_BLOCK_4 std_PG_5_63 ( .p2(\p_vector[4][63] ), .g2(\g_vector[4][63] ), 
        .p1(\p_vector[4][47] ), .g1(\g_vector[4][47] ), .PG_P(
        \p_vector[5][63] ), .PG_G(\g_vector[5][63] ) );
  PG_BLOCK_3 add_PG_5_63_1 ( .p2(\p_vector[4][59] ), .g2(\g_vector[4][59] ), 
        .p1(\p_vector[4][47] ), .g1(\g_vector[4][47] ), .PG_P(
        \p_vector[5][59] ), .PG_G(\g_vector[5][59] ) );
  PG_BLOCK_2 add_PG_5_63_2 ( .p2(\p_vector[3][55] ), .g2(\g_vector[3][55] ), 
        .p1(\p_vector[4][47] ), .g1(\g_vector[4][47] ), .PG_P(
        \p_vector[5][55] ), .PG_G(\g_vector[5][55] ) );
  PG_BLOCK_1 add_PG_5_63_3 ( .p2(\p_vector[2][51] ), .g2(\g_vector[2][51] ), 
        .p1(\p_vector[4][47] ), .g1(\g_vector[4][47] ), .PG_P(
        \p_vector[5][51] ), .PG_G(\g_vector[5][51] ) );
  G_BLOCK_12 std_G_5_31 ( .p2(\p_vector[4][31] ), .g2(\g_vector[4][31] ), .g1(
        Co[3]), .G(Co[7]) );
  G_BLOCK_11 add_G_5_31_1 ( .p2(\p_vector[4][27] ), .g2(\g_vector[4][27] ), 
        .g1(Co[3]), .G(Co[6]) );
  G_BLOCK_10 add_G_5_31_2 ( .p2(\p_vector[3][23] ), .g2(\g_vector[3][23] ), 
        .g1(Co[3]), .G(Co[5]) );
  G_BLOCK_9 add_G_5_31_3 ( .p2(\p_vector[2][19] ), .g2(\g_vector[2][19] ), 
        .g1(Co[3]), .G(Co[4]) );
  G_BLOCK_8 std_G_6_63 ( .p2(\p_vector[5][63] ), .g2(\g_vector[5][63] ), .g1(
        Co[7]), .G(Co[15]) );
  G_BLOCK_7 add_G_6_63_1 ( .p2(\p_vector[5][59] ), .g2(\g_vector[5][59] ), 
        .g1(Co[7]), .G(Co[14]) );
  G_BLOCK_6 add_G_6_63_2 ( .p2(\p_vector[5][55] ), .g2(\g_vector[5][55] ), 
        .g1(Co[7]), .G(Co[13]) );
  G_BLOCK_5 add_G_6_63_3 ( .p2(\p_vector[5][51] ), .g2(\g_vector[5][51] ), 
        .g1(Co[7]), .G(Co[12]) );
  G_BLOCK_4 add_G_6_63_4 ( .p2(\p_vector[4][47] ), .g2(\g_vector[4][47] ), 
        .g1(Co[7]), .G(Co[11]) );
  G_BLOCK_3 add_G_6_63_5 ( .p2(\p_vector[4][43] ), .g2(\g_vector[4][43] ), 
        .g1(Co[7]), .G(Co[10]) );
  G_BLOCK_2 add_G_6_63_6 ( .p2(\p_vector[3][39] ), .g2(\g_vector[3][39] ), 
        .g1(Co[7]), .G(Co[9]) );
  G_BLOCK_1 add_G_6_63_7 ( .p2(\p_vector[2][35] ), .g2(\g_vector[2][35] ), 
        .g1(Co[7]), .G(Co[8]) );
  OAI21_X1 U1 ( .B1(n2), .B2(n1), .A(n4), .ZN(\g_vector[0][0] ) );
  OAI21_X1 U2 ( .B1(A[0]), .B2(B[0]), .A(Cin), .ZN(n4) );
  INV_X1 U3 ( .A(A[0]), .ZN(n2) );
  INV_X1 U4 ( .A(B[0]), .ZN(n1) );
endmodule


module FA_128 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_127 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_126 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_125 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_32 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_128 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_127 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_126 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_125 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_124 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_123 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_122 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_121 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_31 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_124 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_123 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_122 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_121 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_64 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_63 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_62 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_61 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_GENERIC_NBIT4_16 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_64 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_63 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_62 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_61 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_16 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_32 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_31 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_16 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module FA_120 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_119 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_118 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_117 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_30 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_120 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_119 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_118 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_117 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_116 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_115 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_114 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_113 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_29 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_116 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_115 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_114 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_113 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_60 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_59 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_58 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_57 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_GENERIC_NBIT4_15 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_60 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_59 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_58 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_57 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_15 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_30 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_29 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_15 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module FA_112 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_111 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_110 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_109 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_28 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_112 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_111 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_110 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_109 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_108 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_107 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_106 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_105 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_27 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_108 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_107 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_106 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_105 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_56 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_55 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_54 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_53 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_GENERIC_NBIT4_14 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_56 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_55 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_54 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_53 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_14 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_28 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_27 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_14 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module FA_104 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_103 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_102 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_101 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_26 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_104 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_103 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_102 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_101 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_100 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_99 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_98 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_97 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_25 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_100 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_99 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_98 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_97 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_52 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_51 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_50 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_49 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_GENERIC_NBIT4_13 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_52 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_51 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_50 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_49 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_13 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_26 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_25 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_13 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module FA_96 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_95 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_94 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_93 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_24 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_96 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_95 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_94 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_93 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_92 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_91 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_90 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_89 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_23 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_92 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_91 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_90 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_89 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_48 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_47 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_46 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_45 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_GENERIC_NBIT4_12 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_48 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_47 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_46 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_45 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_12 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_24 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_23 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_12 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module FA_88 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_87 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_86 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_85 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_22 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_88 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_87 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_86 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_85 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_84 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_83 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_82 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_81 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_21 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_84 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_83 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_82 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_81 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_44 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_43 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_42 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_41 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_GENERIC_NBIT4_11 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_44 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_43 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_42 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_41 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_11 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_22 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_21 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_11 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module FA_80 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_79 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_78 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_77 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_20 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_80 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_79 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_78 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_77 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_76 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_75 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_74 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_73 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_19 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_76 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_75 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_74 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_73 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_40 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_39 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_38 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_37 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_GENERIC_NBIT4_10 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_40 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_39 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_38 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_37 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_10 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_20 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_19 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_10 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module FA_72 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_71 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_70 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_69 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_18 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_72 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_71 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_70 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_69 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_68 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_67 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_66 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_65 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_17 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_68 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_67 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_66 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_65 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_36 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_35 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_34 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_33 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_GENERIC_NBIT4_9 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_36 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_35 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_34 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_33 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_9 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_18 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_17 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_9 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module FA_64 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_63 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_62 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_61 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_16 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_64 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_63 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_62 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_61 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_60 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_59 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_58 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_57 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_15 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_60 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_59 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_58 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_57 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_32 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_31 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_30 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_29 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_GENERIC_NBIT4_8 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_32 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_31 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_30 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_29 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_8 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_16 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_15 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_8 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module FA_56 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_55 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_54 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_53 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_14 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_56 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_55 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_54 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_53 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_52 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_51 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_50 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_49 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_13 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_52 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_51 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_50 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_49 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_28 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_27 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_26 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_25 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_GENERIC_NBIT4_7 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_28 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_27 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_26 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_25 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_7 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_14 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_13 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_7 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module FA_48 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_47 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_46 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_45 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_12 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_48 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_47 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_46 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_45 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_44 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_43 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_42 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_41 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_11 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_44 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_43 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_42 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_41 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_24 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_23 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_22 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_21 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_GENERIC_NBIT4_6 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_24 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_23 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_22 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_21 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_6 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_12 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_11 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_6 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module FA_40 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_39 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_38 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_37 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_10 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_40 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_39 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_38 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_37 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_36 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_35 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_34 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_33 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_9 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_36 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_35 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_34 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_33 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_20 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_19 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_18 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_17 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_GENERIC_NBIT4_5 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_20 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_19 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_18 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_17 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_5 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_10 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_9 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_5 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module FA_32 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_31 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_30 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_29 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_8 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_32 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_31 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_30 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_29 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_28 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_27 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_26 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_25 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_7 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_28 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_27 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_26 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_25 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_16 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_15 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_14 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_13 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_GENERIC_NBIT4_4 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_16 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_15 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_14 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_13 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_4 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_8 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_7 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_4 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module FA_24 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_23 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_22 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_21 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_6 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_24 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_23 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_22 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_21 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_20 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_19 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_18 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_17 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_5 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_20 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_19 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_18 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_17 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_12 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_11 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_10 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_9 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_GENERIC_NBIT4_3 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_12 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_11 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_10 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_9 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_3 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_6 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_5 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_3 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module FA_16 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_15 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_14 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_13 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_4 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_16 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_15 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_14 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_13 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_12 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_11 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_10 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_9 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_3 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_12 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_11 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_10 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_9 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_8 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_7 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_6 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_5 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_GENERIC_NBIT4_2 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_8 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_7 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_6 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_5 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_2 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_4 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_3 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_2 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module FA_8 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_7 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_6 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_5 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_2 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_8 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_7 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_6 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_5 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module FA_4 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_3 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_2 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module RCA_GEN_NBIT4_1 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_4 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_3 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_2 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module MUX21_4 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_3 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_2 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_1 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n2, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n2), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n2) );
endmodule


module MUX21_GENERIC_NBIT4_1 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_4 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_3 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_2 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_1 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module carry_select_block_n4_1 ( A, B, C_sel, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input C_sel;

  wire   [3:0] sum0;
  wire   [3:0] sum1;

  RCA_GEN_NBIT4_2 RCA0 ( .A(A), .B(B), .Ci(1'b0), .S(sum0) );
  RCA_GEN_NBIT4_1 RCA1 ( .A(A), .B(B), .Ci(1'b1), .S(sum1) );
  MUX21_GENERIC_NBIT4_1 mux ( .A(sum0), .B(sum1), .SEL(C_sel), .Y(S) );
endmodule


module sum_generator_n_bit64_n_CSB16_1 ( A, B, C_in, S );
  input [63:0] A;
  input [63:0] B;
  input [15:0] C_in;
  output [63:0] S;


  carry_select_block_n4_16 csb_0 ( .A(A[3:0]), .B(B[3:0]), .C_sel(C_in[0]), 
        .S(S[3:0]) );
  carry_select_block_n4_15 csb_1 ( .A(A[7:4]), .B(B[7:4]), .C_sel(C_in[1]), 
        .S(S[7:4]) );
  carry_select_block_n4_14 csb_2 ( .A(A[11:8]), .B(B[11:8]), .C_sel(C_in[2]), 
        .S(S[11:8]) );
  carry_select_block_n4_13 csb_3 ( .A(A[15:12]), .B(B[15:12]), .C_sel(C_in[3]), 
        .S(S[15:12]) );
  carry_select_block_n4_12 csb_4 ( .A(A[19:16]), .B(B[19:16]), .C_sel(C_in[4]), 
        .S(S[19:16]) );
  carry_select_block_n4_11 csb_5 ( .A(A[23:20]), .B(B[23:20]), .C_sel(C_in[5]), 
        .S(S[23:20]) );
  carry_select_block_n4_10 csb_6 ( .A(A[27:24]), .B(B[27:24]), .C_sel(C_in[6]), 
        .S(S[27:24]) );
  carry_select_block_n4_9 csb_7 ( .A(A[31:28]), .B(B[31:28]), .C_sel(C_in[7]), 
        .S(S[31:28]) );
  carry_select_block_n4_8 csb_8 ( .A(A[35:32]), .B(B[35:32]), .C_sel(C_in[8]), 
        .S(S[35:32]) );
  carry_select_block_n4_7 csb_9 ( .A(A[39:36]), .B(B[39:36]), .C_sel(C_in[9]), 
        .S(S[39:36]) );
  carry_select_block_n4_6 csb_10 ( .A(A[43:40]), .B(B[43:40]), .C_sel(C_in[10]), .S(S[43:40]) );
  carry_select_block_n4_5 csb_11 ( .A(A[47:44]), .B(B[47:44]), .C_sel(C_in[11]), .S(S[47:44]) );
  carry_select_block_n4_4 csb_12 ( .A(A[51:48]), .B(B[51:48]), .C_sel(C_in[12]), .S(S[51:48]) );
  carry_select_block_n4_3 csb_13 ( .A(A[55:52]), .B(B[55:52]), .C_sel(C_in[13]), .S(S[55:52]) );
  carry_select_block_n4_2 csb_14 ( .A(A[59:56]), .B(B[59:56]), .C_sel(C_in[14]), .S(S[59:56]) );
  carry_select_block_n4_1 csb_15 ( .A(A[63:60]), .B(B[63:60]), .C_sel(C_in[15]), .S(S[63:60]) );
endmodule


module P4_ADDER_NBIT64_1 ( A, B, Cin, S, Cout, ovf );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Cin;
  output Cout, ovf;
  wire   n3, n4;
  wire   [63:0] xor_b;
  wire   [14:0] carry;

  XOR2_X1 U3 ( .A(xor_b[63]), .B(A[63]), .Z(n3) );
  my_xor_64 bc_xor_63 ( .A(B[63]), .B(Cin), .xor_out(xor_b[63]) );
  my_xor_63 bc_xor_62 ( .A(B[62]), .B(Cin), .xor_out(xor_b[62]) );
  my_xor_62 bc_xor_61 ( .A(B[61]), .B(Cin), .xor_out(xor_b[61]) );
  my_xor_61 bc_xor_60 ( .A(B[60]), .B(Cin), .xor_out(xor_b[60]) );
  my_xor_60 bc_xor_59 ( .A(B[59]), .B(Cin), .xor_out(xor_b[59]) );
  my_xor_59 bc_xor_58 ( .A(B[58]), .B(Cin), .xor_out(xor_b[58]) );
  my_xor_58 bc_xor_57 ( .A(B[57]), .B(Cin), .xor_out(xor_b[57]) );
  my_xor_57 bc_xor_56 ( .A(B[56]), .B(Cin), .xor_out(xor_b[56]) );
  my_xor_56 bc_xor_55 ( .A(B[55]), .B(Cin), .xor_out(xor_b[55]) );
  my_xor_55 bc_xor_54 ( .A(B[54]), .B(Cin), .xor_out(xor_b[54]) );
  my_xor_54 bc_xor_53 ( .A(B[53]), .B(Cin), .xor_out(xor_b[53]) );
  my_xor_53 bc_xor_52 ( .A(B[52]), .B(Cin), .xor_out(xor_b[52]) );
  my_xor_52 bc_xor_51 ( .A(B[51]), .B(Cin), .xor_out(xor_b[51]) );
  my_xor_51 bc_xor_50 ( .A(B[50]), .B(Cin), .xor_out(xor_b[50]) );
  my_xor_50 bc_xor_49 ( .A(B[49]), .B(Cin), .xor_out(xor_b[49]) );
  my_xor_49 bc_xor_48 ( .A(B[48]), .B(Cin), .xor_out(xor_b[48]) );
  my_xor_48 bc_xor_47 ( .A(B[47]), .B(Cin), .xor_out(xor_b[47]) );
  my_xor_47 bc_xor_46 ( .A(B[46]), .B(Cin), .xor_out(xor_b[46]) );
  my_xor_46 bc_xor_45 ( .A(B[45]), .B(Cin), .xor_out(xor_b[45]) );
  my_xor_45 bc_xor_44 ( .A(B[44]), .B(Cin), .xor_out(xor_b[44]) );
  my_xor_44 bc_xor_43 ( .A(B[43]), .B(Cin), .xor_out(xor_b[43]) );
  my_xor_43 bc_xor_42 ( .A(B[42]), .B(Cin), .xor_out(xor_b[42]) );
  my_xor_42 bc_xor_41 ( .A(B[41]), .B(Cin), .xor_out(xor_b[41]) );
  my_xor_41 bc_xor_40 ( .A(B[40]), .B(Cin), .xor_out(xor_b[40]) );
  my_xor_40 bc_xor_39 ( .A(B[39]), .B(Cin), .xor_out(xor_b[39]) );
  my_xor_39 bc_xor_38 ( .A(B[38]), .B(Cin), .xor_out(xor_b[38]) );
  my_xor_38 bc_xor_37 ( .A(B[37]), .B(Cin), .xor_out(xor_b[37]) );
  my_xor_37 bc_xor_36 ( .A(B[36]), .B(Cin), .xor_out(xor_b[36]) );
  my_xor_36 bc_xor_35 ( .A(B[35]), .B(Cin), .xor_out(xor_b[35]) );
  my_xor_35 bc_xor_34 ( .A(B[34]), .B(Cin), .xor_out(xor_b[34]) );
  my_xor_34 bc_xor_33 ( .A(B[33]), .B(Cin), .xor_out(xor_b[33]) );
  my_xor_33 bc_xor_32 ( .A(B[32]), .B(Cin), .xor_out(xor_b[32]) );
  my_xor_32 bc_xor_31 ( .A(B[31]), .B(Cin), .xor_out(xor_b[31]) );
  my_xor_31 bc_xor_30 ( .A(B[30]), .B(Cin), .xor_out(xor_b[30]) );
  my_xor_30 bc_xor_29 ( .A(B[29]), .B(Cin), .xor_out(xor_b[29]) );
  my_xor_29 bc_xor_28 ( .A(B[28]), .B(Cin), .xor_out(xor_b[28]) );
  my_xor_28 bc_xor_27 ( .A(B[27]), .B(Cin), .xor_out(xor_b[27]) );
  my_xor_27 bc_xor_26 ( .A(B[26]), .B(Cin), .xor_out(xor_b[26]) );
  my_xor_26 bc_xor_25 ( .A(B[25]), .B(Cin), .xor_out(xor_b[25]) );
  my_xor_25 bc_xor_24 ( .A(B[24]), .B(Cin), .xor_out(xor_b[24]) );
  my_xor_24 bc_xor_23 ( .A(B[23]), .B(Cin), .xor_out(xor_b[23]) );
  my_xor_23 bc_xor_22 ( .A(B[22]), .B(Cin), .xor_out(xor_b[22]) );
  my_xor_22 bc_xor_21 ( .A(B[21]), .B(Cin), .xor_out(xor_b[21]) );
  my_xor_21 bc_xor_20 ( .A(B[20]), .B(Cin), .xor_out(xor_b[20]) );
  my_xor_20 bc_xor_19 ( .A(B[19]), .B(Cin), .xor_out(xor_b[19]) );
  my_xor_19 bc_xor_18 ( .A(B[18]), .B(Cin), .xor_out(xor_b[18]) );
  my_xor_18 bc_xor_17 ( .A(B[17]), .B(Cin), .xor_out(xor_b[17]) );
  my_xor_17 bc_xor_16 ( .A(B[16]), .B(Cin), .xor_out(xor_b[16]) );
  my_xor_16 bc_xor_15 ( .A(B[15]), .B(Cin), .xor_out(xor_b[15]) );
  my_xor_15 bc_xor_14 ( .A(B[14]), .B(Cin), .xor_out(xor_b[14]) );
  my_xor_14 bc_xor_13 ( .A(B[13]), .B(Cin), .xor_out(xor_b[13]) );
  my_xor_13 bc_xor_12 ( .A(B[12]), .B(Cin), .xor_out(xor_b[12]) );
  my_xor_12 bc_xor_11 ( .A(B[11]), .B(Cin), .xor_out(xor_b[11]) );
  my_xor_11 bc_xor_10 ( .A(B[10]), .B(Cin), .xor_out(xor_b[10]) );
  my_xor_10 bc_xor_9 ( .A(B[9]), .B(Cin), .xor_out(xor_b[9]) );
  my_xor_9 bc_xor_8 ( .A(B[8]), .B(Cin), .xor_out(xor_b[8]) );
  my_xor_8 bc_xor_7 ( .A(B[7]), .B(Cin), .xor_out(xor_b[7]) );
  my_xor_7 bc_xor_6 ( .A(B[6]), .B(Cin), .xor_out(xor_b[6]) );
  my_xor_6 bc_xor_5 ( .A(B[5]), .B(Cin), .xor_out(xor_b[5]) );
  my_xor_5 bc_xor_4 ( .A(B[4]), .B(Cin), .xor_out(xor_b[4]) );
  my_xor_4 bc_xor_3 ( .A(B[3]), .B(Cin), .xor_out(xor_b[3]) );
  my_xor_3 bc_xor_2 ( .A(B[2]), .B(Cin), .xor_out(xor_b[2]) );
  my_xor_2 bc_xor_1 ( .A(B[1]), .B(Cin), .xor_out(xor_b[1]) );
  my_xor_1 bc_xor_0 ( .A(B[0]), .B(Cin), .xor_out(xor_b[0]) );
  CARRY_GENERATOR_NBIT64_NBIT_PER_BLOCK4_1 CG ( .A(A), .B(xor_b), .Cin(Cin), 
        .Co({Cout, carry}) );
  sum_generator_n_bit64_n_CSB16_1 SG ( .A(A), .B(xor_b), .C_in({carry, Cin}), 
        .S(S) );
  NOR2_X1 U1 ( .A1(n4), .A2(n3), .ZN(ovf) );
  XNOR2_X1 U2 ( .A(A[63]), .B(S[63]), .ZN(n4) );
endmodule


module boothmul_NBIT_in32 ( A, B, mulin_flag, CLK, RST, MULready, P );
  input [31:0] A;
  input [31:0] B;
  output [63:0] P;
  input mulin_flag, CLK, RST;
  output MULready;
  wire   flag_reg1, flag_reg2, \s_sel[3][2] , \s_sel[3][1] , \s_sel[3][0] ,
         \s_sel[2][2] , \s_sel[2][1] , \s_sel[2][0] , \s_sel[1][2] ,
         \s_sel[1][1] , \s_sel[1][0] , \s_sel[0][2] , \s_sel[0][1] ,
         \s_sel[0][0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60;
  wire   [31:0] mux1_reg1;
  wire   [31:0] mux2_reg1;
  wire   [31:0] A4_reg1;
  wire   [31:0] mux_reg2;
  wire   [63:0] sum_reg2;
  wire   [31:0] A4_reg2;
  wire   [31:0] mux_reg3;
  wire   [63:0] sum_reg3;
  wire   [2:0] enc_reg21;
  wire   [2:0] enc_reg31;
  wire   [2:0] enc_reg32;
  wire   [31:0] mux1_out;
  wire   [31:0] mux2_out;
  wire   [31:0] s_8A_1;
  wire   [31:0] mux_2_out;
  wire   [63:0] sum_2_out;
  wire   [31:0] s_2A_2;
  wire   [31:0] mux_3_out;
  wire   [63:0] sum_3_out;
  wire   [31:0] s_2A_1;
  wire   [31:0] s_4A_1;
  wire   [31:0] s_A_neg;
  wire   [31:0] s_2A_1_neg;
  wire   [31:0] s_4A_1_neg;
  wire   [31:0] s_8A_1_neg;
  wire   [31:0] s_A_2;
  wire   [31:0] s_A_2_neg;
  wire   [31:0] s_2A_2_neg;
  wire   [31:0] s_A_3;
  wire   [31:0] s_2A_3;
  wire   [31:0] s_A_3_neg;
  wire   [31:0] s_2A_3_neg;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11;

  DFFR_X1 flag_reg1_reg ( .D(mulin_flag), .CK(CLK), .RN(n60), .Q(flag_reg1) );
  DFFR_X1 \mux1_reg1_reg[31]  ( .D(mux1_out[31]), .CK(CLK), .RN(n60), .Q(
        mux1_reg1[31]) );
  DFFR_X1 \mux1_reg1_reg[30]  ( .D(mux1_out[30]), .CK(CLK), .RN(n59), .Q(
        mux1_reg1[30]) );
  DFFR_X1 \mux1_reg1_reg[29]  ( .D(mux1_out[29]), .CK(CLK), .RN(n59), .Q(
        mux1_reg1[29]) );
  DFFR_X1 \mux1_reg1_reg[28]  ( .D(mux1_out[28]), .CK(CLK), .RN(n59), .Q(
        mux1_reg1[28]) );
  DFFR_X1 \mux1_reg1_reg[27]  ( .D(mux1_out[27]), .CK(CLK), .RN(n59), .Q(
        mux1_reg1[27]) );
  DFFR_X1 \mux1_reg1_reg[26]  ( .D(mux1_out[26]), .CK(CLK), .RN(n59), .Q(
        mux1_reg1[26]) );
  DFFR_X1 \mux1_reg1_reg[25]  ( .D(mux1_out[25]), .CK(CLK), .RN(n59), .Q(
        mux1_reg1[25]) );
  DFFR_X1 \mux1_reg1_reg[24]  ( .D(mux1_out[24]), .CK(CLK), .RN(n59), .Q(
        mux1_reg1[24]) );
  DFFR_X1 \mux1_reg1_reg[23]  ( .D(mux1_out[23]), .CK(CLK), .RN(n59), .Q(
        mux1_reg1[23]) );
  DFFR_X1 \mux1_reg1_reg[22]  ( .D(mux1_out[22]), .CK(CLK), .RN(n59), .Q(
        mux1_reg1[22]) );
  DFFR_X1 \mux1_reg1_reg[21]  ( .D(mux1_out[21]), .CK(CLK), .RN(n59), .Q(
        mux1_reg1[21]) );
  DFFR_X1 \mux1_reg1_reg[20]  ( .D(mux1_out[20]), .CK(CLK), .RN(n59), .Q(
        mux1_reg1[20]) );
  DFFR_X1 \mux1_reg1_reg[19]  ( .D(mux1_out[19]), .CK(CLK), .RN(n58), .Q(
        mux1_reg1[19]) );
  DFFR_X1 \mux1_reg1_reg[18]  ( .D(mux1_out[18]), .CK(CLK), .RN(n58), .Q(
        mux1_reg1[18]) );
  DFFR_X1 \mux1_reg1_reg[17]  ( .D(mux1_out[17]), .CK(CLK), .RN(n58), .Q(
        mux1_reg1[17]) );
  DFFR_X1 \mux1_reg1_reg[16]  ( .D(mux1_out[16]), .CK(CLK), .RN(n58), .Q(
        mux1_reg1[16]) );
  DFFR_X1 \mux1_reg1_reg[15]  ( .D(mux1_out[15]), .CK(CLK), .RN(n58), .Q(
        mux1_reg1[15]) );
  DFFR_X1 \mux1_reg1_reg[14]  ( .D(mux1_out[14]), .CK(CLK), .RN(n58), .Q(
        mux1_reg1[14]) );
  DFFR_X1 \mux1_reg1_reg[13]  ( .D(mux1_out[13]), .CK(CLK), .RN(n58), .Q(
        mux1_reg1[13]) );
  DFFR_X1 \mux1_reg1_reg[12]  ( .D(mux1_out[12]), .CK(CLK), .RN(n58), .Q(
        mux1_reg1[12]) );
  DFFR_X1 \mux1_reg1_reg[11]  ( .D(mux1_out[11]), .CK(CLK), .RN(n58), .Q(
        mux1_reg1[11]) );
  DFFR_X1 \mux1_reg1_reg[10]  ( .D(mux1_out[10]), .CK(CLK), .RN(n58), .Q(
        mux1_reg1[10]) );
  DFFR_X1 \mux1_reg1_reg[9]  ( .D(mux1_out[9]), .CK(CLK), .RN(n58), .Q(
        mux1_reg1[9]) );
  DFFR_X1 \mux1_reg1_reg[8]  ( .D(mux1_out[8]), .CK(CLK), .RN(n57), .Q(
        mux1_reg1[8]) );
  DFFR_X1 \mux1_reg1_reg[7]  ( .D(mux1_out[7]), .CK(CLK), .RN(n57), .Q(
        mux1_reg1[7]) );
  DFFR_X1 \mux1_reg1_reg[6]  ( .D(mux1_out[6]), .CK(CLK), .RN(n57), .Q(
        mux1_reg1[6]) );
  DFFR_X1 \mux1_reg1_reg[5]  ( .D(mux1_out[5]), .CK(CLK), .RN(n57), .Q(
        mux1_reg1[5]) );
  DFFR_X1 \mux1_reg1_reg[4]  ( .D(mux1_out[4]), .CK(CLK), .RN(n57), .Q(
        mux1_reg1[4]) );
  DFFR_X1 \mux1_reg1_reg[3]  ( .D(mux1_out[3]), .CK(CLK), .RN(n57), .Q(
        mux1_reg1[3]) );
  DFFR_X1 \mux1_reg1_reg[2]  ( .D(mux1_out[2]), .CK(CLK), .RN(n57), .Q(
        mux1_reg1[2]) );
  DFFR_X1 \mux1_reg1_reg[1]  ( .D(mux1_out[1]), .CK(CLK), .RN(n57), .Q(
        mux1_reg1[1]) );
  DFFR_X1 \mux1_reg1_reg[0]  ( .D(mux1_out[0]), .CK(CLK), .RN(n57), .Q(
        mux1_reg1[0]) );
  DFFR_X1 \mux2_reg1_reg[31]  ( .D(mux2_out[31]), .CK(CLK), .RN(n57), .Q(
        mux2_reg1[31]) );
  DFFR_X1 \mux2_reg1_reg[30]  ( .D(mux2_out[30]), .CK(CLK), .RN(n57), .Q(
        mux2_reg1[30]) );
  DFFR_X1 \mux2_reg1_reg[29]  ( .D(mux2_out[29]), .CK(CLK), .RN(n56), .Q(
        mux2_reg1[29]) );
  DFFR_X1 \mux2_reg1_reg[28]  ( .D(mux2_out[28]), .CK(CLK), .RN(n56), .Q(
        mux2_reg1[28]) );
  DFFR_X1 \mux2_reg1_reg[27]  ( .D(mux2_out[27]), .CK(CLK), .RN(n56), .Q(
        mux2_reg1[27]) );
  DFFR_X1 \mux2_reg1_reg[26]  ( .D(mux2_out[26]), .CK(CLK), .RN(n56), .Q(
        mux2_reg1[26]) );
  DFFR_X1 \mux2_reg1_reg[25]  ( .D(mux2_out[25]), .CK(CLK), .RN(n56), .Q(
        mux2_reg1[25]) );
  DFFR_X1 \mux2_reg1_reg[24]  ( .D(mux2_out[24]), .CK(CLK), .RN(n56), .Q(
        mux2_reg1[24]) );
  DFFR_X1 \mux2_reg1_reg[23]  ( .D(mux2_out[23]), .CK(CLK), .RN(n56), .Q(
        mux2_reg1[23]) );
  DFFR_X1 \mux2_reg1_reg[22]  ( .D(mux2_out[22]), .CK(CLK), .RN(n56), .Q(
        mux2_reg1[22]) );
  DFFR_X1 \mux2_reg1_reg[21]  ( .D(mux2_out[21]), .CK(CLK), .RN(n56), .Q(
        mux2_reg1[21]) );
  DFFR_X1 \mux2_reg1_reg[20]  ( .D(mux2_out[20]), .CK(CLK), .RN(n56), .Q(
        mux2_reg1[20]) );
  DFFR_X1 \mux2_reg1_reg[19]  ( .D(mux2_out[19]), .CK(CLK), .RN(n56), .Q(
        mux2_reg1[19]) );
  DFFR_X1 \mux2_reg1_reg[18]  ( .D(mux2_out[18]), .CK(CLK), .RN(n55), .Q(
        mux2_reg1[18]) );
  DFFR_X1 \mux2_reg1_reg[17]  ( .D(mux2_out[17]), .CK(CLK), .RN(n55), .Q(
        mux2_reg1[17]) );
  DFFR_X1 \mux2_reg1_reg[16]  ( .D(mux2_out[16]), .CK(CLK), .RN(n55), .Q(
        mux2_reg1[16]) );
  DFFR_X1 \mux2_reg1_reg[15]  ( .D(mux2_out[15]), .CK(CLK), .RN(n55), .Q(
        mux2_reg1[15]) );
  DFFR_X1 \mux2_reg1_reg[14]  ( .D(mux2_out[14]), .CK(CLK), .RN(n55), .Q(
        mux2_reg1[14]) );
  DFFR_X1 \mux2_reg1_reg[13]  ( .D(mux2_out[13]), .CK(CLK), .RN(n55), .Q(
        mux2_reg1[13]) );
  DFFR_X1 \mux2_reg1_reg[12]  ( .D(mux2_out[12]), .CK(CLK), .RN(n55), .Q(
        mux2_reg1[12]) );
  DFFR_X1 \mux2_reg1_reg[11]  ( .D(mux2_out[11]), .CK(CLK), .RN(n55), .Q(
        mux2_reg1[11]) );
  DFFR_X1 \mux2_reg1_reg[10]  ( .D(mux2_out[10]), .CK(CLK), .RN(n55), .Q(
        mux2_reg1[10]) );
  DFFR_X1 \mux2_reg1_reg[9]  ( .D(mux2_out[9]), .CK(CLK), .RN(n55), .Q(
        mux2_reg1[9]) );
  DFFR_X1 \mux2_reg1_reg[8]  ( .D(mux2_out[8]), .CK(CLK), .RN(n55), .Q(
        mux2_reg1[8]) );
  DFFR_X1 \mux2_reg1_reg[7]  ( .D(mux2_out[7]), .CK(CLK), .RN(n54), .Q(
        mux2_reg1[7]) );
  DFFR_X1 \mux2_reg1_reg[6]  ( .D(mux2_out[6]), .CK(CLK), .RN(n54), .Q(
        mux2_reg1[6]) );
  DFFR_X1 \mux2_reg1_reg[5]  ( .D(mux2_out[5]), .CK(CLK), .RN(n54), .Q(
        mux2_reg1[5]) );
  DFFR_X1 \mux2_reg1_reg[4]  ( .D(mux2_out[4]), .CK(CLK), .RN(n54), .Q(
        mux2_reg1[4]) );
  DFFR_X1 \mux2_reg1_reg[3]  ( .D(mux2_out[3]), .CK(CLK), .RN(n54), .Q(
        mux2_reg1[3]) );
  DFFR_X1 \mux2_reg1_reg[2]  ( .D(mux2_out[2]), .CK(CLK), .RN(n54), .Q(
        mux2_reg1[2]) );
  DFFR_X1 \mux2_reg1_reg[1]  ( .D(mux2_out[1]), .CK(CLK), .RN(n54), .Q(
        mux2_reg1[1]) );
  DFFR_X1 \mux2_reg1_reg[0]  ( .D(mux2_out[0]), .CK(CLK), .RN(n54), .Q(
        mux2_reg1[0]) );
  DFFR_X1 \A4_reg1_reg[31]  ( .D(s_8A_1[31]), .CK(CLK), .RN(n54), .Q(
        A4_reg1[31]) );
  DFFR_X1 \A4_reg1_reg[30]  ( .D(s_8A_1[30]), .CK(CLK), .RN(n54), .Q(
        A4_reg1[30]) );
  DFFR_X1 \A4_reg1_reg[29]  ( .D(s_8A_1[29]), .CK(CLK), .RN(n54), .Q(
        A4_reg1[29]) );
  DFFR_X1 \A4_reg1_reg[28]  ( .D(s_8A_1[28]), .CK(CLK), .RN(n53), .Q(
        A4_reg1[28]) );
  DFFR_X1 \A4_reg1_reg[27]  ( .D(s_8A_1[27]), .CK(CLK), .RN(n53), .Q(
        A4_reg1[27]) );
  DFFR_X1 \A4_reg1_reg[26]  ( .D(s_8A_1[26]), .CK(CLK), .RN(n53), .Q(
        A4_reg1[26]) );
  DFFR_X1 \A4_reg1_reg[25]  ( .D(s_8A_1[25]), .CK(CLK), .RN(n53), .Q(
        A4_reg1[25]) );
  DFFR_X1 \A4_reg1_reg[24]  ( .D(s_8A_1[24]), .CK(CLK), .RN(n53), .Q(
        A4_reg1[24]) );
  DFFR_X1 \A4_reg1_reg[23]  ( .D(s_8A_1[23]), .CK(CLK), .RN(n53), .Q(
        A4_reg1[23]) );
  DFFR_X1 \A4_reg1_reg[22]  ( .D(s_8A_1[22]), .CK(CLK), .RN(n53), .Q(
        A4_reg1[22]) );
  DFFR_X1 \A4_reg1_reg[21]  ( .D(s_8A_1[21]), .CK(CLK), .RN(n53), .Q(
        A4_reg1[21]) );
  DFFR_X1 \A4_reg1_reg[20]  ( .D(s_8A_1[20]), .CK(CLK), .RN(n53), .Q(
        A4_reg1[20]) );
  DFFR_X1 \A4_reg1_reg[19]  ( .D(s_8A_1[19]), .CK(CLK), .RN(n53), .Q(
        A4_reg1[19]) );
  DFFR_X1 \A4_reg1_reg[18]  ( .D(s_8A_1[18]), .CK(CLK), .RN(n53), .Q(
        A4_reg1[18]) );
  DFFR_X1 \A4_reg1_reg[17]  ( .D(s_8A_1[17]), .CK(CLK), .RN(n52), .Q(
        A4_reg1[17]) );
  DFFR_X1 \A4_reg1_reg[16]  ( .D(s_8A_1[16]), .CK(CLK), .RN(n52), .Q(
        A4_reg1[16]) );
  DFFR_X1 \A4_reg1_reg[15]  ( .D(s_8A_1[15]), .CK(CLK), .RN(n52), .Q(
        A4_reg1[15]) );
  DFFR_X1 \A4_reg1_reg[14]  ( .D(s_8A_1[14]), .CK(CLK), .RN(n52), .Q(
        A4_reg1[14]) );
  DFFR_X1 \A4_reg1_reg[13]  ( .D(s_8A_1[13]), .CK(CLK), .RN(n52), .Q(
        A4_reg1[13]) );
  DFFR_X1 \A4_reg1_reg[12]  ( .D(s_8A_1[12]), .CK(CLK), .RN(n52), .Q(
        A4_reg1[12]) );
  DFFR_X1 \A4_reg1_reg[11]  ( .D(s_8A_1[11]), .CK(CLK), .RN(n52), .Q(
        A4_reg1[11]) );
  DFFR_X1 \A4_reg1_reg[10]  ( .D(s_8A_1[10]), .CK(CLK), .RN(n52), .Q(
        A4_reg1[10]) );
  DFFR_X1 \A4_reg1_reg[9]  ( .D(s_8A_1[9]), .CK(CLK), .RN(n52), .Q(A4_reg1[9])
         );
  DFFR_X1 \A4_reg1_reg[8]  ( .D(s_8A_1[8]), .CK(CLK), .RN(n52), .Q(A4_reg1[8])
         );
  DFFR_X1 \A4_reg1_reg[7]  ( .D(s_8A_1[7]), .CK(CLK), .RN(n52), .Q(A4_reg1[7])
         );
  DFFR_X1 \A4_reg1_reg[6]  ( .D(s_8A_1[6]), .CK(CLK), .RN(n51), .Q(A4_reg1[6])
         );
  DFFR_X1 \A4_reg1_reg[5]  ( .D(s_8A_1[5]), .CK(CLK), .RN(n51), .Q(A4_reg1[5])
         );
  DFFR_X1 \A4_reg1_reg[4]  ( .D(s_8A_1[4]), .CK(CLK), .RN(n51), .Q(A4_reg1[4])
         );
  DFFR_X1 \A4_reg1_reg[3]  ( .D(s_8A_1[3]), .CK(CLK), .RN(n51), .Q(A4_reg1[3])
         );
  DFFR_X1 flag_reg2_reg ( .D(flag_reg1), .CK(CLK), .RN(n51), .Q(flag_reg2) );
  DFFR_X1 \sum_reg2_reg[63]  ( .D(sum_2_out[63]), .CK(CLK), .RN(n51), .Q(
        sum_reg2[63]) );
  DFFR_X1 \sum_reg2_reg[62]  ( .D(sum_2_out[62]), .CK(CLK), .RN(n51), .Q(
        sum_reg2[62]) );
  DFFR_X1 \sum_reg2_reg[61]  ( .D(sum_2_out[61]), .CK(CLK), .RN(n51), .Q(
        sum_reg2[61]) );
  DFFR_X1 \sum_reg2_reg[60]  ( .D(sum_2_out[60]), .CK(CLK), .RN(n50), .Q(
        sum_reg2[60]) );
  DFFR_X1 \sum_reg2_reg[59]  ( .D(sum_2_out[59]), .CK(CLK), .RN(n50), .Q(
        sum_reg2[59]) );
  DFFR_X1 \sum_reg2_reg[58]  ( .D(sum_2_out[58]), .CK(CLK), .RN(n50), .Q(
        sum_reg2[58]) );
  DFFR_X1 \sum_reg2_reg[57]  ( .D(sum_2_out[57]), .CK(CLK), .RN(n50), .Q(
        sum_reg2[57]) );
  DFFR_X1 \sum_reg2_reg[56]  ( .D(sum_2_out[56]), .CK(CLK), .RN(n50), .Q(
        sum_reg2[56]) );
  DFFR_X1 \sum_reg2_reg[55]  ( .D(sum_2_out[55]), .CK(CLK), .RN(n50), .Q(
        sum_reg2[55]) );
  DFFR_X1 \sum_reg2_reg[54]  ( .D(sum_2_out[54]), .CK(CLK), .RN(n50), .Q(
        sum_reg2[54]) );
  DFFR_X1 \sum_reg2_reg[53]  ( .D(sum_2_out[53]), .CK(CLK), .RN(n50), .Q(
        sum_reg2[53]) );
  DFFR_X1 \sum_reg2_reg[52]  ( .D(sum_2_out[52]), .CK(CLK), .RN(n50), .Q(
        sum_reg2[52]) );
  DFFR_X1 \sum_reg2_reg[51]  ( .D(sum_2_out[51]), .CK(CLK), .RN(n50), .Q(
        sum_reg2[51]) );
  DFFR_X1 \sum_reg2_reg[50]  ( .D(sum_2_out[50]), .CK(CLK), .RN(n50), .Q(
        sum_reg2[50]) );
  DFFR_X1 \sum_reg2_reg[49]  ( .D(sum_2_out[49]), .CK(CLK), .RN(n49), .Q(
        sum_reg2[49]) );
  DFFR_X1 \sum_reg2_reg[48]  ( .D(sum_2_out[48]), .CK(CLK), .RN(n49), .Q(
        sum_reg2[48]) );
  DFFR_X1 \sum_reg2_reg[47]  ( .D(sum_2_out[47]), .CK(CLK), .RN(n49), .Q(
        sum_reg2[47]) );
  DFFR_X1 \sum_reg2_reg[46]  ( .D(sum_2_out[46]), .CK(CLK), .RN(n49), .Q(
        sum_reg2[46]) );
  DFFR_X1 \sum_reg2_reg[45]  ( .D(sum_2_out[45]), .CK(CLK), .RN(n49), .Q(
        sum_reg2[45]) );
  DFFR_X1 \sum_reg2_reg[44]  ( .D(sum_2_out[44]), .CK(CLK), .RN(n49), .Q(
        sum_reg2[44]) );
  DFFR_X1 \sum_reg2_reg[43]  ( .D(sum_2_out[43]), .CK(CLK), .RN(n49), .Q(
        sum_reg2[43]) );
  DFFR_X1 \sum_reg2_reg[42]  ( .D(sum_2_out[42]), .CK(CLK), .RN(n49), .Q(
        sum_reg2[42]) );
  DFFR_X1 \sum_reg2_reg[41]  ( .D(sum_2_out[41]), .CK(CLK), .RN(n49), .Q(
        sum_reg2[41]) );
  DFFR_X1 \sum_reg2_reg[40]  ( .D(sum_2_out[40]), .CK(CLK), .RN(n49), .Q(
        sum_reg2[40]) );
  DFFR_X1 \sum_reg2_reg[39]  ( .D(sum_2_out[39]), .CK(CLK), .RN(n49), .Q(
        sum_reg2[39]) );
  DFFR_X1 \sum_reg2_reg[38]  ( .D(sum_2_out[38]), .CK(CLK), .RN(n48), .Q(
        sum_reg2[38]) );
  DFFR_X1 \sum_reg2_reg[37]  ( .D(sum_2_out[37]), .CK(CLK), .RN(n48), .Q(
        sum_reg2[37]) );
  DFFR_X1 \sum_reg2_reg[36]  ( .D(sum_2_out[36]), .CK(CLK), .RN(n48), .Q(
        sum_reg2[36]) );
  DFFR_X1 \sum_reg2_reg[35]  ( .D(sum_2_out[35]), .CK(CLK), .RN(n48), .Q(
        sum_reg2[35]) );
  DFFR_X1 \sum_reg2_reg[34]  ( .D(sum_2_out[34]), .CK(CLK), .RN(n48), .Q(
        sum_reg2[34]) );
  DFFR_X1 \sum_reg2_reg[33]  ( .D(sum_2_out[33]), .CK(CLK), .RN(n48), .Q(
        sum_reg2[33]) );
  DFFR_X1 \sum_reg2_reg[32]  ( .D(sum_2_out[32]), .CK(CLK), .RN(n48), .Q(
        sum_reg2[32]) );
  DFFR_X1 \sum_reg2_reg[31]  ( .D(sum_2_out[31]), .CK(CLK), .RN(n48), .Q(
        sum_reg2[31]) );
  DFFR_X1 \sum_reg2_reg[30]  ( .D(sum_2_out[30]), .CK(CLK), .RN(n48), .Q(
        sum_reg2[30]) );
  DFFR_X1 \sum_reg2_reg[29]  ( .D(sum_2_out[29]), .CK(CLK), .RN(n48), .Q(
        sum_reg2[29]) );
  DFFR_X1 \sum_reg2_reg[28]  ( .D(sum_2_out[28]), .CK(CLK), .RN(n48), .Q(
        sum_reg2[28]) );
  DFFR_X1 \sum_reg2_reg[27]  ( .D(sum_2_out[27]), .CK(CLK), .RN(n47), .Q(
        sum_reg2[27]) );
  DFFR_X1 \sum_reg2_reg[26]  ( .D(sum_2_out[26]), .CK(CLK), .RN(n47), .Q(
        sum_reg2[26]) );
  DFFR_X1 \sum_reg2_reg[25]  ( .D(sum_2_out[25]), .CK(CLK), .RN(n47), .Q(
        sum_reg2[25]) );
  DFFR_X1 \sum_reg2_reg[24]  ( .D(sum_2_out[24]), .CK(CLK), .RN(n47), .Q(
        sum_reg2[24]) );
  DFFR_X1 \sum_reg2_reg[23]  ( .D(sum_2_out[23]), .CK(CLK), .RN(n47), .Q(
        sum_reg2[23]) );
  DFFR_X1 \sum_reg2_reg[22]  ( .D(sum_2_out[22]), .CK(CLK), .RN(n47), .Q(
        sum_reg2[22]) );
  DFFR_X1 \sum_reg2_reg[21]  ( .D(sum_2_out[21]), .CK(CLK), .RN(n47), .Q(
        sum_reg2[21]) );
  DFFR_X1 \sum_reg2_reg[20]  ( .D(sum_2_out[20]), .CK(CLK), .RN(n47), .Q(
        sum_reg2[20]) );
  DFFR_X1 \sum_reg2_reg[19]  ( .D(sum_2_out[19]), .CK(CLK), .RN(n47), .Q(
        sum_reg2[19]) );
  DFFR_X1 \sum_reg2_reg[18]  ( .D(sum_2_out[18]), .CK(CLK), .RN(n47), .Q(
        sum_reg2[18]) );
  DFFR_X1 \sum_reg2_reg[17]  ( .D(sum_2_out[17]), .CK(CLK), .RN(n47), .Q(
        sum_reg2[17]) );
  DFFR_X1 \sum_reg2_reg[16]  ( .D(sum_2_out[16]), .CK(CLK), .RN(n46), .Q(
        sum_reg2[16]) );
  DFFR_X1 \sum_reg2_reg[15]  ( .D(sum_2_out[15]), .CK(CLK), .RN(n46), .Q(
        sum_reg2[15]) );
  DFFR_X1 \sum_reg2_reg[14]  ( .D(sum_2_out[14]), .CK(CLK), .RN(n46), .Q(
        sum_reg2[14]) );
  DFFR_X1 \sum_reg2_reg[13]  ( .D(sum_2_out[13]), .CK(CLK), .RN(n46), .Q(
        sum_reg2[13]) );
  DFFR_X1 \sum_reg2_reg[12]  ( .D(sum_2_out[12]), .CK(CLK), .RN(n46), .Q(
        sum_reg2[12]) );
  DFFR_X1 \sum_reg2_reg[11]  ( .D(sum_2_out[11]), .CK(CLK), .RN(n46), .Q(
        sum_reg2[11]) );
  DFFR_X1 \sum_reg2_reg[10]  ( .D(sum_2_out[10]), .CK(CLK), .RN(n46), .Q(
        sum_reg2[10]) );
  DFFR_X1 \sum_reg2_reg[9]  ( .D(sum_2_out[9]), .CK(CLK), .RN(n46), .Q(
        sum_reg2[9]) );
  DFFR_X1 \sum_reg2_reg[8]  ( .D(sum_2_out[8]), .CK(CLK), .RN(n46), .Q(
        sum_reg2[8]) );
  DFFR_X1 \sum_reg2_reg[7]  ( .D(sum_2_out[7]), .CK(CLK), .RN(n46), .Q(
        sum_reg2[7]) );
  DFFR_X1 \sum_reg2_reg[6]  ( .D(sum_2_out[6]), .CK(CLK), .RN(n46), .Q(
        sum_reg2[6]) );
  DFFR_X1 \sum_reg2_reg[5]  ( .D(sum_2_out[5]), .CK(CLK), .RN(n45), .Q(
        sum_reg2[5]) );
  DFFR_X1 \sum_reg2_reg[4]  ( .D(sum_2_out[4]), .CK(CLK), .RN(n45), .Q(
        sum_reg2[4]) );
  DFFR_X1 \sum_reg2_reg[3]  ( .D(sum_2_out[3]), .CK(CLK), .RN(n45), .Q(
        sum_reg2[3]) );
  DFFR_X1 \sum_reg2_reg[2]  ( .D(sum_2_out[2]), .CK(CLK), .RN(n45), .Q(
        sum_reg2[2]) );
  DFFR_X1 \sum_reg2_reg[1]  ( .D(sum_2_out[1]), .CK(CLK), .RN(n45), .Q(
        sum_reg2[1]) );
  DFFR_X1 \sum_reg2_reg[0]  ( .D(sum_2_out[0]), .CK(CLK), .RN(n45), .Q(
        sum_reg2[0]) );
  DFFR_X1 \A4_reg2_reg[31]  ( .D(s_2A_2[31]), .CK(CLK), .RN(n45), .Q(
        A4_reg2[31]) );
  DFFR_X1 \A4_reg2_reg[30]  ( .D(s_2A_2[30]), .CK(CLK), .RN(n45), .Q(
        A4_reg2[30]) );
  DFFR_X1 \A4_reg2_reg[29]  ( .D(s_2A_2[29]), .CK(CLK), .RN(n45), .Q(
        A4_reg2[29]) );
  DFFR_X1 \A4_reg2_reg[28]  ( .D(s_2A_2[28]), .CK(CLK), .RN(n45), .Q(
        A4_reg2[28]) );
  DFFR_X1 \A4_reg2_reg[27]  ( .D(s_2A_2[27]), .CK(CLK), .RN(n45), .Q(
        A4_reg2[27]) );
  DFFR_X1 \A4_reg2_reg[26]  ( .D(s_2A_2[26]), .CK(CLK), .RN(n44), .Q(
        A4_reg2[26]) );
  DFFR_X1 \A4_reg2_reg[25]  ( .D(s_2A_2[25]), .CK(CLK), .RN(n44), .Q(
        A4_reg2[25]) );
  DFFR_X1 \A4_reg2_reg[24]  ( .D(s_2A_2[24]), .CK(CLK), .RN(n44), .Q(
        A4_reg2[24]) );
  DFFR_X1 \A4_reg2_reg[23]  ( .D(s_2A_2[23]), .CK(CLK), .RN(n44), .Q(
        A4_reg2[23]) );
  DFFR_X1 \A4_reg2_reg[22]  ( .D(s_2A_2[22]), .CK(CLK), .RN(n44), .Q(
        A4_reg2[22]) );
  DFFR_X1 \A4_reg2_reg[21]  ( .D(s_2A_2[21]), .CK(CLK), .RN(n44), .Q(
        A4_reg2[21]) );
  DFFR_X1 \A4_reg2_reg[20]  ( .D(s_2A_2[20]), .CK(CLK), .RN(n44), .Q(
        A4_reg2[20]) );
  DFFR_X1 \A4_reg2_reg[19]  ( .D(s_2A_2[19]), .CK(CLK), .RN(n44), .Q(
        A4_reg2[19]) );
  DFFR_X1 \A4_reg2_reg[18]  ( .D(s_2A_2[18]), .CK(CLK), .RN(n44), .Q(
        A4_reg2[18]) );
  DFFR_X1 \A4_reg2_reg[17]  ( .D(s_2A_2[17]), .CK(CLK), .RN(n44), .Q(
        A4_reg2[17]) );
  DFFR_X1 \A4_reg2_reg[16]  ( .D(s_2A_2[16]), .CK(CLK), .RN(n44), .Q(
        A4_reg2[16]) );
  DFFR_X1 \A4_reg2_reg[15]  ( .D(s_2A_2[15]), .CK(CLK), .RN(n43), .Q(
        A4_reg2[15]) );
  DFFR_X1 \A4_reg2_reg[14]  ( .D(s_2A_2[14]), .CK(CLK), .RN(n43), .Q(
        A4_reg2[14]) );
  DFFR_X1 \A4_reg2_reg[13]  ( .D(s_2A_2[13]), .CK(CLK), .RN(n43), .Q(
        A4_reg2[13]) );
  DFFR_X1 \A4_reg2_reg[12]  ( .D(s_2A_2[12]), .CK(CLK), .RN(n43), .Q(
        A4_reg2[12]) );
  DFFR_X1 \A4_reg2_reg[11]  ( .D(s_2A_2[11]), .CK(CLK), .RN(n43), .Q(
        A4_reg2[11]) );
  DFFR_X1 \A4_reg2_reg[10]  ( .D(s_2A_2[10]), .CK(CLK), .RN(n43), .Q(
        A4_reg2[10]) );
  DFFR_X1 \A4_reg2_reg[9]  ( .D(s_2A_2[9]), .CK(CLK), .RN(n43), .Q(A4_reg2[9])
         );
  DFFR_X1 \A4_reg2_reg[8]  ( .D(s_2A_2[8]), .CK(CLK), .RN(n43), .Q(A4_reg2[8])
         );
  DFFR_X1 \A4_reg2_reg[7]  ( .D(s_2A_2[7]), .CK(CLK), .RN(n43), .Q(A4_reg2[7])
         );
  DFFR_X1 \A4_reg2_reg[6]  ( .D(s_2A_2[6]), .CK(CLK), .RN(n43), .Q(A4_reg2[6])
         );
  DFFR_X1 \A4_reg2_reg[5]  ( .D(s_2A_2[5]), .CK(CLK), .RN(n43), .Q(A4_reg2[5])
         );
  DFFR_X1 \A4_reg2_reg[4]  ( .D(s_2A_2[4]), .CK(CLK), .RN(n42), .Q(A4_reg2[4])
         );
  DFFR_X1 \A4_reg2_reg[3]  ( .D(s_2A_2[3]), .CK(CLK), .RN(n42), .Q(A4_reg2[3])
         );
  DFFR_X1 \A4_reg2_reg[2]  ( .D(s_2A_2[2]), .CK(CLK), .RN(n42), .Q(A4_reg2[2])
         );
  DFFR_X1 flag_reg3_reg ( .D(flag_reg2), .CK(CLK), .RN(n42), .Q(MULready) );
  DFFR_X1 \enc_reg21_reg[2]  ( .D(\s_sel[2][2] ), .CK(CLK), .RN(n42), .Q(
        enc_reg21[2]) );
  DFFR_X1 \enc_reg21_reg[1]  ( .D(\s_sel[2][1] ), .CK(CLK), .RN(n42), .Q(
        enc_reg21[1]) );
  DFFR_X1 \enc_reg21_reg[0]  ( .D(\s_sel[2][0] ), .CK(CLK), .RN(n42), .Q(
        enc_reg21[0]) );
  DFFR_X1 \mux_reg2_reg[0]  ( .D(mux_2_out[0]), .CK(CLK), .RN(n42), .Q(
        mux_reg2[0]) );
  DFFR_X1 \mux_reg2_reg[1]  ( .D(mux_2_out[1]), .CK(CLK), .RN(n42), .Q(
        mux_reg2[1]) );
  DFFR_X1 \mux_reg2_reg[2]  ( .D(mux_2_out[2]), .CK(CLK), .RN(n41), .Q(
        mux_reg2[2]) );
  DFFR_X1 \mux_reg2_reg[3]  ( .D(mux_2_out[3]), .CK(CLK), .RN(n41), .Q(
        mux_reg2[3]) );
  DFFR_X1 \mux_reg2_reg[4]  ( .D(mux_2_out[4]), .CK(CLK), .RN(n41), .Q(
        mux_reg2[4]) );
  DFFR_X1 \mux_reg2_reg[5]  ( .D(mux_2_out[5]), .CK(CLK), .RN(n41), .Q(
        mux_reg2[5]) );
  DFFR_X1 \mux_reg2_reg[6]  ( .D(mux_2_out[6]), .CK(CLK), .RN(n41), .Q(
        mux_reg2[6]) );
  DFFR_X1 \mux_reg2_reg[7]  ( .D(mux_2_out[7]), .CK(CLK), .RN(n41), .Q(
        mux_reg2[7]) );
  DFFR_X1 \mux_reg2_reg[8]  ( .D(mux_2_out[8]), .CK(CLK), .RN(n41), .Q(
        mux_reg2[8]) );
  DFFR_X1 \mux_reg2_reg[9]  ( .D(mux_2_out[9]), .CK(CLK), .RN(n41), .Q(
        mux_reg2[9]) );
  DFFR_X1 \mux_reg2_reg[10]  ( .D(mux_2_out[10]), .CK(CLK), .RN(n41), .Q(
        mux_reg2[10]) );
  DFFR_X1 \mux_reg2_reg[11]  ( .D(mux_2_out[11]), .CK(CLK), .RN(n41), .Q(
        mux_reg2[11]) );
  DFFR_X1 \mux_reg2_reg[12]  ( .D(mux_2_out[12]), .CK(CLK), .RN(n41), .Q(
        mux_reg2[12]) );
  DFFR_X1 \mux_reg2_reg[13]  ( .D(mux_2_out[13]), .CK(CLK), .RN(n40), .Q(
        mux_reg2[13]) );
  DFFR_X1 \mux_reg2_reg[14]  ( .D(mux_2_out[14]), .CK(CLK), .RN(n40), .Q(
        mux_reg2[14]) );
  DFFR_X1 \mux_reg2_reg[15]  ( .D(mux_2_out[15]), .CK(CLK), .RN(n40), .Q(
        mux_reg2[15]) );
  DFFR_X1 \mux_reg2_reg[16]  ( .D(mux_2_out[16]), .CK(CLK), .RN(n40), .Q(
        mux_reg2[16]) );
  DFFR_X1 \mux_reg2_reg[17]  ( .D(mux_2_out[17]), .CK(CLK), .RN(n40), .Q(
        mux_reg2[17]) );
  DFFR_X1 \mux_reg2_reg[18]  ( .D(mux_2_out[18]), .CK(CLK), .RN(n40), .Q(
        mux_reg2[18]) );
  DFFR_X1 \mux_reg2_reg[19]  ( .D(mux_2_out[19]), .CK(CLK), .RN(n40), .Q(
        mux_reg2[19]) );
  DFFR_X1 \mux_reg2_reg[20]  ( .D(mux_2_out[20]), .CK(CLK), .RN(n40), .Q(
        mux_reg2[20]) );
  DFFR_X1 \mux_reg2_reg[21]  ( .D(mux_2_out[21]), .CK(CLK), .RN(n40), .Q(
        mux_reg2[21]) );
  DFFR_X1 \mux_reg2_reg[22]  ( .D(mux_2_out[22]), .CK(CLK), .RN(n40), .Q(
        mux_reg2[22]) );
  DFFR_X1 \mux_reg2_reg[23]  ( .D(mux_2_out[23]), .CK(CLK), .RN(n40), .Q(
        mux_reg2[23]) );
  DFFR_X1 \mux_reg2_reg[24]  ( .D(mux_2_out[24]), .CK(CLK), .RN(n39), .Q(
        mux_reg2[24]) );
  DFFR_X1 \mux_reg2_reg[25]  ( .D(mux_2_out[25]), .CK(CLK), .RN(n39), .Q(
        mux_reg2[25]) );
  DFFR_X1 \mux_reg2_reg[26]  ( .D(mux_2_out[26]), .CK(CLK), .RN(n39), .Q(
        mux_reg2[26]) );
  DFFR_X1 \mux_reg2_reg[27]  ( .D(mux_2_out[27]), .CK(CLK), .RN(n39), .Q(
        mux_reg2[27]) );
  DFFR_X1 \mux_reg2_reg[28]  ( .D(mux_2_out[28]), .CK(CLK), .RN(n39), .Q(
        mux_reg2[28]) );
  DFFR_X1 \mux_reg2_reg[29]  ( .D(mux_2_out[29]), .CK(CLK), .RN(n39), .Q(
        mux_reg2[29]) );
  DFFR_X1 \mux_reg2_reg[30]  ( .D(mux_2_out[30]), .CK(CLK), .RN(n39), .Q(
        mux_reg2[30]) );
  DFFR_X1 \mux_reg2_reg[31]  ( .D(mux_2_out[31]), .CK(CLK), .RN(n39), .Q(
        mux_reg2[31]) );
  DFFR_X1 \sum_reg3_reg[0]  ( .D(sum_3_out[0]), .CK(CLK), .RN(n39), .Q(
        sum_reg3[0]) );
  DFFR_X1 \sum_reg3_reg[1]  ( .D(sum_3_out[1]), .CK(CLK), .RN(n39), .Q(
        sum_reg3[1]) );
  DFFR_X1 \sum_reg3_reg[2]  ( .D(sum_3_out[2]), .CK(CLK), .RN(n39), .Q(
        sum_reg3[2]) );
  DFFR_X1 \sum_reg3_reg[3]  ( .D(sum_3_out[3]), .CK(CLK), .RN(n38), .Q(
        sum_reg3[3]) );
  DFFR_X1 \sum_reg3_reg[4]  ( .D(sum_3_out[4]), .CK(CLK), .RN(n38), .Q(
        sum_reg3[4]) );
  DFFR_X1 \sum_reg3_reg[5]  ( .D(sum_3_out[5]), .CK(CLK), .RN(n38), .Q(
        sum_reg3[5]) );
  DFFR_X1 \sum_reg3_reg[6]  ( .D(sum_3_out[6]), .CK(CLK), .RN(n38), .Q(
        sum_reg3[6]) );
  DFFR_X1 \sum_reg3_reg[7]  ( .D(sum_3_out[7]), .CK(CLK), .RN(n38), .Q(
        sum_reg3[7]) );
  DFFR_X1 \sum_reg3_reg[8]  ( .D(sum_3_out[8]), .CK(CLK), .RN(n38), .Q(
        sum_reg3[8]) );
  DFFR_X1 \sum_reg3_reg[9]  ( .D(sum_3_out[9]), .CK(CLK), .RN(n38), .Q(
        sum_reg3[9]) );
  DFFR_X1 \sum_reg3_reg[10]  ( .D(sum_3_out[10]), .CK(CLK), .RN(n38), .Q(
        sum_reg3[10]) );
  DFFR_X1 \sum_reg3_reg[11]  ( .D(sum_3_out[11]), .CK(CLK), .RN(n38), .Q(
        sum_reg3[11]) );
  DFFR_X1 \sum_reg3_reg[12]  ( .D(sum_3_out[12]), .CK(CLK), .RN(n38), .Q(
        sum_reg3[12]) );
  DFFR_X1 \sum_reg3_reg[13]  ( .D(sum_3_out[13]), .CK(CLK), .RN(n38), .Q(
        sum_reg3[13]) );
  DFFR_X1 \sum_reg3_reg[14]  ( .D(sum_3_out[14]), .CK(CLK), .RN(n37), .Q(
        sum_reg3[14]) );
  DFFR_X1 \sum_reg3_reg[15]  ( .D(sum_3_out[15]), .CK(CLK), .RN(n37), .Q(
        sum_reg3[15]) );
  DFFR_X1 \sum_reg3_reg[16]  ( .D(sum_3_out[16]), .CK(CLK), .RN(n37), .Q(
        sum_reg3[16]) );
  DFFR_X1 \sum_reg3_reg[17]  ( .D(sum_3_out[17]), .CK(CLK), .RN(n37), .Q(
        sum_reg3[17]) );
  DFFR_X1 \sum_reg3_reg[18]  ( .D(sum_3_out[18]), .CK(CLK), .RN(n37), .Q(
        sum_reg3[18]) );
  DFFR_X1 \sum_reg3_reg[19]  ( .D(sum_3_out[19]), .CK(CLK), .RN(n37), .Q(
        sum_reg3[19]) );
  DFFR_X1 \sum_reg3_reg[20]  ( .D(sum_3_out[20]), .CK(CLK), .RN(n37), .Q(
        sum_reg3[20]) );
  DFFR_X1 \sum_reg3_reg[21]  ( .D(sum_3_out[21]), .CK(CLK), .RN(n37), .Q(
        sum_reg3[21]) );
  DFFR_X1 \sum_reg3_reg[22]  ( .D(sum_3_out[22]), .CK(CLK), .RN(n37), .Q(
        sum_reg3[22]) );
  DFFR_X1 \sum_reg3_reg[23]  ( .D(sum_3_out[23]), .CK(CLK), .RN(n37), .Q(
        sum_reg3[23]) );
  DFFR_X1 \sum_reg3_reg[24]  ( .D(sum_3_out[24]), .CK(CLK), .RN(n37), .Q(
        sum_reg3[24]) );
  DFFR_X1 \sum_reg3_reg[25]  ( .D(sum_3_out[25]), .CK(CLK), .RN(n36), .Q(
        sum_reg3[25]) );
  DFFR_X1 \sum_reg3_reg[26]  ( .D(sum_3_out[26]), .CK(CLK), .RN(n36), .Q(
        sum_reg3[26]) );
  DFFR_X1 \sum_reg3_reg[27]  ( .D(sum_3_out[27]), .CK(CLK), .RN(n36), .Q(
        sum_reg3[27]) );
  DFFR_X1 \sum_reg3_reg[28]  ( .D(sum_3_out[28]), .CK(CLK), .RN(n36), .Q(
        sum_reg3[28]) );
  DFFR_X1 \sum_reg3_reg[29]  ( .D(sum_3_out[29]), .CK(CLK), .RN(n36), .Q(
        sum_reg3[29]) );
  DFFR_X1 \sum_reg3_reg[30]  ( .D(sum_3_out[30]), .CK(CLK), .RN(n36), .Q(
        sum_reg3[30]) );
  DFFR_X1 \sum_reg3_reg[31]  ( .D(sum_3_out[31]), .CK(CLK), .RN(n36), .Q(
        sum_reg3[31]) );
  DFFR_X1 \sum_reg3_reg[32]  ( .D(sum_3_out[32]), .CK(CLK), .RN(n36), .Q(
        sum_reg3[32]) );
  DFFR_X1 \sum_reg3_reg[33]  ( .D(sum_3_out[33]), .CK(CLK), .RN(n36), .Q(
        sum_reg3[33]) );
  DFFR_X1 \sum_reg3_reg[34]  ( .D(sum_3_out[34]), .CK(CLK), .RN(n36), .Q(
        sum_reg3[34]) );
  DFFR_X1 \sum_reg3_reg[35]  ( .D(sum_3_out[35]), .CK(CLK), .RN(n36), .Q(
        sum_reg3[35]) );
  DFFR_X1 \sum_reg3_reg[36]  ( .D(sum_3_out[36]), .CK(CLK), .RN(n35), .Q(
        sum_reg3[36]) );
  DFFR_X1 \sum_reg3_reg[37]  ( .D(sum_3_out[37]), .CK(CLK), .RN(n35), .Q(
        sum_reg3[37]) );
  DFFR_X1 \sum_reg3_reg[38]  ( .D(sum_3_out[38]), .CK(CLK), .RN(n35), .Q(
        sum_reg3[38]) );
  DFFR_X1 \sum_reg3_reg[39]  ( .D(sum_3_out[39]), .CK(CLK), .RN(n35), .Q(
        sum_reg3[39]) );
  DFFR_X1 \sum_reg3_reg[40]  ( .D(sum_3_out[40]), .CK(CLK), .RN(n35), .Q(
        sum_reg3[40]) );
  DFFR_X1 \sum_reg3_reg[41]  ( .D(sum_3_out[41]), .CK(CLK), .RN(n35), .Q(
        sum_reg3[41]) );
  DFFR_X1 \sum_reg3_reg[42]  ( .D(sum_3_out[42]), .CK(CLK), .RN(n35), .Q(
        sum_reg3[42]) );
  DFFR_X1 \sum_reg3_reg[43]  ( .D(sum_3_out[43]), .CK(CLK), .RN(n35), .Q(
        sum_reg3[43]) );
  DFFR_X1 \sum_reg3_reg[44]  ( .D(sum_3_out[44]), .CK(CLK), .RN(n35), .Q(
        sum_reg3[44]) );
  DFFR_X1 \sum_reg3_reg[45]  ( .D(sum_3_out[45]), .CK(CLK), .RN(n35), .Q(
        sum_reg3[45]) );
  DFFR_X1 \sum_reg3_reg[46]  ( .D(sum_3_out[46]), .CK(CLK), .RN(n35), .Q(
        sum_reg3[46]) );
  DFFR_X1 \sum_reg3_reg[47]  ( .D(sum_3_out[47]), .CK(CLK), .RN(n34), .Q(
        sum_reg3[47]) );
  DFFR_X1 \sum_reg3_reg[48]  ( .D(sum_3_out[48]), .CK(CLK), .RN(n34), .Q(
        sum_reg3[48]) );
  DFFR_X1 \sum_reg3_reg[49]  ( .D(sum_3_out[49]), .CK(CLK), .RN(n34), .Q(
        sum_reg3[49]) );
  DFFR_X1 \sum_reg3_reg[50]  ( .D(sum_3_out[50]), .CK(CLK), .RN(n34), .Q(
        sum_reg3[50]) );
  DFFR_X1 \sum_reg3_reg[51]  ( .D(sum_3_out[51]), .CK(CLK), .RN(n34), .Q(
        sum_reg3[51]) );
  DFFR_X1 \sum_reg3_reg[52]  ( .D(sum_3_out[52]), .CK(CLK), .RN(n34), .Q(
        sum_reg3[52]) );
  DFFR_X1 \sum_reg3_reg[53]  ( .D(sum_3_out[53]), .CK(CLK), .RN(n34), .Q(
        sum_reg3[53]) );
  DFFR_X1 \sum_reg3_reg[54]  ( .D(sum_3_out[54]), .CK(CLK), .RN(n34), .Q(
        sum_reg3[54]) );
  DFFR_X1 \sum_reg3_reg[55]  ( .D(sum_3_out[55]), .CK(CLK), .RN(n34), .Q(
        sum_reg3[55]) );
  DFFR_X1 \sum_reg3_reg[56]  ( .D(sum_3_out[56]), .CK(CLK), .RN(n34), .Q(
        sum_reg3[56]) );
  DFFR_X1 \sum_reg3_reg[57]  ( .D(sum_3_out[57]), .CK(CLK), .RN(n34), .Q(
        sum_reg3[57]) );
  DFFR_X1 \sum_reg3_reg[58]  ( .D(sum_3_out[58]), .CK(CLK), .RN(n33), .Q(
        sum_reg3[58]) );
  DFFR_X1 \sum_reg3_reg[59]  ( .D(sum_3_out[59]), .CK(CLK), .RN(n33), .Q(
        sum_reg3[59]) );
  DFFR_X1 \sum_reg3_reg[60]  ( .D(sum_3_out[60]), .CK(CLK), .RN(n33), .Q(
        sum_reg3[60]) );
  DFFR_X1 \sum_reg3_reg[61]  ( .D(sum_3_out[61]), .CK(CLK), .RN(n33), .Q(
        sum_reg3[61]) );
  DFFR_X1 \sum_reg3_reg[62]  ( .D(sum_3_out[62]), .CK(CLK), .RN(n33), .Q(
        sum_reg3[62]) );
  DFFR_X1 \sum_reg3_reg[63]  ( .D(sum_3_out[63]), .CK(CLK), .RN(n33), .Q(
        sum_reg3[63]) );
  DFFR_X1 \enc_reg31_reg[2]  ( .D(\s_sel[3][2] ), .CK(CLK), .RN(n33), .Q(
        enc_reg31[2]) );
  DFFR_X1 \enc_reg32_reg[2]  ( .D(enc_reg31[2]), .CK(CLK), .RN(n33), .Q(
        enc_reg32[2]) );
  DFFR_X1 \enc_reg31_reg[1]  ( .D(\s_sel[3][1] ), .CK(CLK), .RN(n33), .Q(
        enc_reg31[1]) );
  DFFR_X1 \enc_reg32_reg[1]  ( .D(enc_reg31[1]), .CK(CLK), .RN(n33), .Q(
        enc_reg32[1]) );
  DFFR_X1 \enc_reg31_reg[0]  ( .D(\s_sel[3][0] ), .CK(CLK), .RN(n33), .Q(
        enc_reg31[0]) );
  DFFR_X1 \enc_reg32_reg[0]  ( .D(enc_reg31[0]), .CK(CLK), .RN(n32), .Q(
        enc_reg32[0]) );
  DFFR_X1 \mux_reg3_reg[0]  ( .D(mux_3_out[0]), .CK(CLK), .RN(n32), .Q(
        mux_reg3[0]) );
  DFFR_X1 \mux_reg3_reg[1]  ( .D(mux_3_out[1]), .CK(CLK), .RN(n32), .Q(
        mux_reg3[1]) );
  DFFR_X1 \mux_reg3_reg[2]  ( .D(mux_3_out[2]), .CK(CLK), .RN(n32), .Q(
        mux_reg3[2]) );
  DFFR_X1 \mux_reg3_reg[3]  ( .D(mux_3_out[3]), .CK(CLK), .RN(n32), .Q(
        mux_reg3[3]) );
  DFFR_X1 \mux_reg3_reg[4]  ( .D(mux_3_out[4]), .CK(CLK), .RN(n32), .Q(
        mux_reg3[4]) );
  DFFR_X1 \mux_reg3_reg[5]  ( .D(mux_3_out[5]), .CK(CLK), .RN(n32), .Q(
        mux_reg3[5]) );
  DFFR_X1 \mux_reg3_reg[6]  ( .D(mux_3_out[6]), .CK(CLK), .RN(n32), .Q(
        mux_reg3[6]) );
  DFFR_X1 \mux_reg3_reg[7]  ( .D(mux_3_out[7]), .CK(CLK), .RN(n32), .Q(
        mux_reg3[7]) );
  DFFR_X1 \mux_reg3_reg[8]  ( .D(mux_3_out[8]), .CK(CLK), .RN(n32), .Q(
        mux_reg3[8]) );
  DFFR_X1 \mux_reg3_reg[9]  ( .D(mux_3_out[9]), .CK(CLK), .RN(n32), .Q(
        mux_reg3[9]) );
  DFFR_X1 \mux_reg3_reg[10]  ( .D(mux_3_out[10]), .CK(CLK), .RN(n31), .Q(
        mux_reg3[10]) );
  DFFR_X1 \mux_reg3_reg[11]  ( .D(mux_3_out[11]), .CK(CLK), .RN(n31), .Q(
        mux_reg3[11]) );
  DFFR_X1 \mux_reg3_reg[12]  ( .D(mux_3_out[12]), .CK(CLK), .RN(n31), .Q(
        mux_reg3[12]) );
  DFFR_X1 \mux_reg3_reg[13]  ( .D(mux_3_out[13]), .CK(CLK), .RN(n31), .Q(
        mux_reg3[13]) );
  DFFR_X1 \mux_reg3_reg[14]  ( .D(mux_3_out[14]), .CK(CLK), .RN(n31), .Q(
        mux_reg3[14]) );
  DFFR_X1 \mux_reg3_reg[15]  ( .D(mux_3_out[15]), .CK(CLK), .RN(n31), .Q(
        mux_reg3[15]) );
  DFFR_X1 \mux_reg3_reg[16]  ( .D(mux_3_out[16]), .CK(CLK), .RN(n31), .Q(
        mux_reg3[16]) );
  DFFR_X1 \mux_reg3_reg[17]  ( .D(mux_3_out[17]), .CK(CLK), .RN(n31), .Q(
        mux_reg3[17]) );
  DFFR_X1 \mux_reg3_reg[18]  ( .D(mux_3_out[18]), .CK(CLK), .RN(n31), .Q(
        mux_reg3[18]) );
  DFFR_X1 \mux_reg3_reg[19]  ( .D(mux_3_out[19]), .CK(CLK), .RN(n31), .Q(
        mux_reg3[19]) );
  DFFR_X1 \mux_reg3_reg[20]  ( .D(mux_3_out[20]), .CK(CLK), .RN(n31), .Q(
        mux_reg3[20]) );
  DFFR_X1 \mux_reg3_reg[21]  ( .D(mux_3_out[21]), .CK(CLK), .RN(n30), .Q(
        mux_reg3[21]) );
  DFFR_X1 \mux_reg3_reg[22]  ( .D(mux_3_out[22]), .CK(CLK), .RN(n30), .Q(
        mux_reg3[22]) );
  DFFR_X1 \mux_reg3_reg[23]  ( .D(mux_3_out[23]), .CK(CLK), .RN(n30), .Q(
        mux_reg3[23]) );
  DFFR_X1 \mux_reg3_reg[24]  ( .D(mux_3_out[24]), .CK(CLK), .RN(n30), .Q(
        mux_reg3[24]) );
  DFFR_X1 \mux_reg3_reg[25]  ( .D(mux_3_out[25]), .CK(CLK), .RN(n30), .Q(
        mux_reg3[25]) );
  DFFR_X1 \mux_reg3_reg[26]  ( .D(mux_3_out[26]), .CK(CLK), .RN(n30), .Q(
        mux_reg3[26]) );
  DFFR_X1 \mux_reg3_reg[27]  ( .D(mux_3_out[27]), .CK(CLK), .RN(n30), .Q(
        mux_reg3[27]) );
  DFFR_X1 \mux_reg3_reg[28]  ( .D(mux_3_out[28]), .CK(CLK), .RN(n30), .Q(
        mux_reg3[28]) );
  DFFR_X1 \mux_reg3_reg[29]  ( .D(mux_3_out[29]), .CK(CLK), .RN(n30), .Q(
        mux_reg3[29]) );
  DFFR_X1 \mux_reg3_reg[30]  ( .D(mux_3_out[30]), .CK(CLK), .RN(n30), .Q(
        mux_reg3[30]) );
  DFFR_X1 \mux_reg3_reg[31]  ( .D(mux_3_out[31]), .CK(CLK), .RN(n30), .Q(
        mux_reg3[31]) );
  enc33_0 enc_0 ( .A({B[1:0], 1'b0}), .Y({\s_sel[0][2] , \s_sel[0][1] , 
        \s_sel[0][0] }) );
  enc33_3 enc_1 ( .A(B[3:1]), .Y({\s_sel[1][2] , \s_sel[1][1] , \s_sel[1][0] }) );
  enc33_2 enc_2 ( .A(B[5:3]), .Y({\s_sel[2][2] , \s_sel[2][1] , \s_sel[2][0] }) );
  enc33_1 enc_3 ( .A(B[7:5]), .Y({\s_sel[3][2] , \s_sel[3][1] , \s_sel[3][0] }) );
  shl1_NBIT32_0 shift2A ( .A({n18, A[30:0]}), .Y({s_2A_1[31:1], 
        SYNOPSYS_UNCONNECTED__0}) );
  shl2_NBIT32_0 shift4A ( .A({n18, A[30:0]}), .Y({s_4A_1[31:2], 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2}) );
  shl3_NBIT32 shift8A ( .A({n18, A[30:0]}), .Y({s_8A_1[31:3], 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5}) );
  negate_NBIT32_0 neg1 ( .A({n18, A[30:0]}), .Y(s_A_neg) );
  negate_NBIT32_7 neg2 ( .A({s_2A_1[31:1], 1'b0}), .Y(s_2A_1_neg) );
  negate_NBIT32_6 neg3 ( .A({s_4A_1[31:2], 1'b0, 1'b0}), .Y(s_4A_1_neg) );
  negate_NBIT32_5 neg4 ( .A({s_8A_1[31:3], 1'b0, 1'b0, 1'b0}), .Y(s_8A_1_neg)
         );
  mux51_gen_NBIT32_0 mux1 ( .A0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .A1({n18, A[30:0]}), .A2(s_A_neg), .A3({s_2A_1[31:1], 1'b0}), 
        .A4(s_2A_1_neg), .SEL({\s_sel[0][2] , \s_sel[0][1] , \s_sel[0][0] }), 
        .Y(mux1_out) );
  mux51_gen_NBIT32_3 mux2 ( .A0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .A1({s_4A_1[31:2], 1'b0, 1'b0}), .A2(s_4A_1_neg), .A3({
        s_8A_1[31:3], 1'b0, 1'b0, 1'b0}), .A4(s_8A_1_neg), .SEL({\s_sel[1][2] , 
        \s_sel[1][1] , \s_sel[1][0] }), .Y(mux2_out) );
  shl1_NBIT32_2 shift2A_2 ( .A({A4_reg1[31:3], 1'b0, 1'b0, 1'b0}), .Y({
        s_A_2[31:1], SYNOPSYS_UNCONNECTED__6}) );
  shl2_NBIT32_2 shift4A_2 ( .A({A4_reg1[31:3], 1'b0, 1'b0, 1'b0}), .Y({
        s_2A_2[31:2], SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8}) );
  negate_NBIT32_4 neg5 ( .A({s_A_2[31:1], 1'b0}), .Y(s_A_2_neg) );
  negate_NBIT32_3 neg6 ( .A({s_2A_2[31:2], 1'b0, 1'b0}), .Y(s_2A_2_neg) );
  mux51_gen_NBIT32_2 mux3 ( .A0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .A1({s_A_2[31:1], 1'b0}), .A2(s_A_2_neg), .A3({s_2A_2[31:2], 
        1'b0, 1'b0}), .A4(s_2A_2_neg), .SEL(enc_reg21), .Y(mux_2_out) );
  P4_ADDER_NBIT64_0 SUM1 ( .A({n12, n12, n12, n12, n12, n13, n13, n13, n13, 
        n13, n13, n14, n14, n14, n14, n14, n14, n15, n15, n15, n15, n15, n15, 
        n16, n16, n16, n16, n16, n16, n17, n17, n17, n17, mux1_reg1[30:0]}), 
        .B({n9, n9, n9, n9, n9, n9, n9, n9, n9, n9, n9, n8, n8, n8, n8, n8, n8, 
        n8, n8, n8, n8, n8, n7, n7, n7, n7, n7, n7, n7, n7, n7, n7, n7, 
        mux2_reg1[30:0]}), .Cin(1'b0), .S(sum_2_out) );
  shl1_NBIT32_1 shift2A_3 ( .A({A4_reg2[31:2], 1'b0, 1'b0}), .Y({s_A_3[31:1], 
        SYNOPSYS_UNCONNECTED__9}) );
  shl2_NBIT32_1 shift4A_3 ( .A({A4_reg2[31:2], 1'b0, 1'b0}), .Y({s_2A_3[31:2], 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11}) );
  negate_NBIT32_2 neg7 ( .A({s_A_3[31:1], 1'b0}), .Y(s_A_3_neg) );
  negate_NBIT32_1 neg8 ( .A({s_2A_3[31:2], 1'b0, 1'b0}), .Y(s_2A_3_neg) );
  mux51_gen_NBIT32_1 mux4 ( .A0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .A1({s_A_3[31:1], 1'b0}), .A2(s_A_3_neg), .A3({s_2A_3[31:2], 
        1'b0, 1'b0}), .A4(s_2A_3_neg), .SEL(enc_reg32), .Y(mux_3_out) );
  P4_ADDER_NBIT64_2 SUM2 ( .A(sum_reg2), .B({n6, n6, n6, n6, n6, n6, n6, n6, 
        n6, n6, n6, n5, n5, n5, n5, n5, n5, n5, n5, n5, n5, n5, n4, n4, n4, n4, 
        n4, n4, n4, n4, n4, n4, n4, mux_reg2[30:0]}), .Cin(1'b0), .S(sum_3_out) );
  P4_ADDER_NBIT64_1 SUM3 ( .A(sum_reg3), .B({n3, n3, n3, n3, n3, n3, n3, n3, 
        n3, n3, n3, n2, n2, n2, n2, n2, n2, n2, n2, n2, n2, n2, n1, n1, n1, n1, 
        n1, n1, n1, n1, n1, n1, n1, mux_reg3[30:0]}), .Cin(1'b0), .S(P) );
  BUF_X1 U3 ( .A(n28), .Z(n21) );
  BUF_X1 U4 ( .A(n28), .Z(n22) );
  BUF_X1 U5 ( .A(n28), .Z(n23) );
  BUF_X1 U6 ( .A(n27), .Z(n24) );
  BUF_X1 U7 ( .A(n27), .Z(n25) );
  BUF_X1 U8 ( .A(n29), .Z(n19) );
  BUF_X1 U9 ( .A(n29), .Z(n20) );
  BUF_X1 U10 ( .A(n27), .Z(n26) );
  BUF_X1 U11 ( .A(RST), .Z(n28) );
  BUF_X1 U12 ( .A(RST), .Z(n27) );
  BUF_X1 U13 ( .A(RST), .Z(n29) );
  BUF_X2 U14 ( .A(n11), .Z(n15) );
  BUF_X2 U15 ( .A(n10), .Z(n13) );
  BUF_X2 U16 ( .A(n11), .Z(n16) );
  BUF_X2 U17 ( .A(n10), .Z(n14) );
  BUF_X2 U18 ( .A(n10), .Z(n12) );
  BUF_X2 U19 ( .A(n11), .Z(n17) );
  BUF_X1 U20 ( .A(A[31]), .Z(n18) );
  BUF_X1 U21 ( .A(mux_reg2[31]), .Z(n5) );
  BUF_X1 U22 ( .A(mux_reg2[31]), .Z(n4) );
  BUF_X1 U23 ( .A(mux2_reg1[31]), .Z(n7) );
  BUF_X1 U24 ( .A(mux2_reg1[31]), .Z(n8) );
  BUF_X1 U25 ( .A(mux2_reg1[31]), .Z(n9) );
  BUF_X1 U26 ( .A(mux_reg2[31]), .Z(n6) );
  BUF_X1 U27 ( .A(mux1_reg1[31]), .Z(n11) );
  BUF_X1 U28 ( .A(mux1_reg1[31]), .Z(n10) );
  BUF_X1 U29 ( .A(mux_reg3[31]), .Z(n1) );
  BUF_X1 U30 ( .A(mux_reg3[31]), .Z(n2) );
  BUF_X1 U31 ( .A(mux_reg3[31]), .Z(n3) );
  CLKBUF_X1 U37 ( .A(n19), .Z(n30) );
  CLKBUF_X1 U38 ( .A(n19), .Z(n31) );
  CLKBUF_X1 U39 ( .A(n19), .Z(n32) );
  CLKBUF_X1 U40 ( .A(n19), .Z(n33) );
  CLKBUF_X1 U41 ( .A(n20), .Z(n34) );
  CLKBUF_X1 U42 ( .A(n20), .Z(n35) );
  CLKBUF_X1 U43 ( .A(n20), .Z(n36) );
  CLKBUF_X1 U44 ( .A(n20), .Z(n37) );
  CLKBUF_X1 U45 ( .A(n21), .Z(n38) );
  CLKBUF_X1 U46 ( .A(n21), .Z(n39) );
  CLKBUF_X1 U47 ( .A(n21), .Z(n40) );
  CLKBUF_X1 U48 ( .A(n21), .Z(n41) );
  CLKBUF_X1 U49 ( .A(n22), .Z(n42) );
  CLKBUF_X1 U50 ( .A(n22), .Z(n43) );
  CLKBUF_X1 U51 ( .A(n22), .Z(n44) );
  CLKBUF_X1 U52 ( .A(n22), .Z(n45) );
  CLKBUF_X1 U53 ( .A(n23), .Z(n46) );
  CLKBUF_X1 U54 ( .A(n23), .Z(n47) );
  CLKBUF_X1 U55 ( .A(n23), .Z(n48) );
  CLKBUF_X1 U56 ( .A(n23), .Z(n49) );
  CLKBUF_X1 U57 ( .A(n24), .Z(n50) );
  CLKBUF_X1 U58 ( .A(n24), .Z(n51) );
  CLKBUF_X1 U59 ( .A(n24), .Z(n52) );
  CLKBUF_X1 U60 ( .A(n24), .Z(n53) );
  CLKBUF_X1 U61 ( .A(n25), .Z(n54) );
  CLKBUF_X1 U62 ( .A(n25), .Z(n55) );
  CLKBUF_X1 U63 ( .A(n25), .Z(n56) );
  CLKBUF_X1 U64 ( .A(n25), .Z(n57) );
  CLKBUF_X1 U65 ( .A(n26), .Z(n58) );
  CLKBUF_X1 U66 ( .A(n26), .Z(n59) );
  CLKBUF_X1 U67 ( .A(n26), .Z(n60) );
endmodule


module MUX21_424 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_423 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_422 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_421 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_420 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_419 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_418 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_417 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_416 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_415 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_414 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_413 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_412 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_411 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_410 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_409 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_408 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_407 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_406 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_405 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_404 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_403 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_402 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_401 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_400 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_399 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_398 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_397 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_396 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_395 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_394 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_393 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_GENERIC_NBIT32_1 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   n1, n2, n3;

  MUX21_424 MUXES_0 ( .A(A[0]), .B(B[0]), .S(n1), .Y(Y[0]) );
  MUX21_423 MUXES_1 ( .A(A[1]), .B(B[1]), .S(n1), .Y(Y[1]) );
  MUX21_422 MUXES_2 ( .A(A[2]), .B(B[2]), .S(n1), .Y(Y[2]) );
  MUX21_421 MUXES_3 ( .A(A[3]), .B(B[3]), .S(n1), .Y(Y[3]) );
  MUX21_420 MUXES_4 ( .A(A[4]), .B(B[4]), .S(n1), .Y(Y[4]) );
  MUX21_419 MUXES_5 ( .A(A[5]), .B(B[5]), .S(n1), .Y(Y[5]) );
  MUX21_418 MUXES_6 ( .A(A[6]), .B(B[6]), .S(n1), .Y(Y[6]) );
  MUX21_417 MUXES_7 ( .A(A[7]), .B(B[7]), .S(n1), .Y(Y[7]) );
  MUX21_416 MUXES_8 ( .A(A[8]), .B(B[8]), .S(n1), .Y(Y[8]) );
  MUX21_415 MUXES_9 ( .A(A[9]), .B(B[9]), .S(n1), .Y(Y[9]) );
  MUX21_414 MUXES_10 ( .A(A[10]), .B(B[10]), .S(n1), .Y(Y[10]) );
  MUX21_413 MUXES_11 ( .A(A[11]), .B(B[11]), .S(n1), .Y(Y[11]) );
  MUX21_412 MUXES_12 ( .A(A[12]), .B(B[12]), .S(n2), .Y(Y[12]) );
  MUX21_411 MUXES_13 ( .A(A[13]), .B(B[13]), .S(n2), .Y(Y[13]) );
  MUX21_410 MUXES_14 ( .A(A[14]), .B(B[14]), .S(n2), .Y(Y[14]) );
  MUX21_409 MUXES_15 ( .A(A[15]), .B(B[15]), .S(n2), .Y(Y[15]) );
  MUX21_408 MUXES_16 ( .A(A[16]), .B(B[16]), .S(n2), .Y(Y[16]) );
  MUX21_407 MUXES_17 ( .A(A[17]), .B(B[17]), .S(n2), .Y(Y[17]) );
  MUX21_406 MUXES_18 ( .A(A[18]), .B(B[18]), .S(n2), .Y(Y[18]) );
  MUX21_405 MUXES_19 ( .A(A[19]), .B(B[19]), .S(n2), .Y(Y[19]) );
  MUX21_404 MUXES_20 ( .A(A[20]), .B(B[20]), .S(n2), .Y(Y[20]) );
  MUX21_403 MUXES_21 ( .A(A[21]), .B(B[21]), .S(n2), .Y(Y[21]) );
  MUX21_402 MUXES_22 ( .A(A[22]), .B(B[22]), .S(n2), .Y(Y[22]) );
  MUX21_401 MUXES_23 ( .A(A[23]), .B(B[23]), .S(n2), .Y(Y[23]) );
  MUX21_400 MUXES_24 ( .A(A[24]), .B(B[24]), .S(n3), .Y(Y[24]) );
  MUX21_399 MUXES_25 ( .A(A[25]), .B(B[25]), .S(n3), .Y(Y[25]) );
  MUX21_398 MUXES_26 ( .A(A[26]), .B(B[26]), .S(n3), .Y(Y[26]) );
  MUX21_397 MUXES_27 ( .A(A[27]), .B(B[27]), .S(n3), .Y(Y[27]) );
  MUX21_396 MUXES_28 ( .A(A[28]), .B(B[28]), .S(n3), .Y(Y[28]) );
  MUX21_395 MUXES_29 ( .A(A[29]), .B(B[29]), .S(n3), .Y(Y[29]) );
  MUX21_394 MUXES_30 ( .A(A[30]), .B(B[30]), .S(n3), .Y(Y[30]) );
  MUX21_393 MUXES_31 ( .A(A[31]), .B(B[31]), .S(n3), .Y(Y[31]) );
  BUF_X1 U1 ( .A(SEL), .Z(n2) );
  BUF_X1 U2 ( .A(SEL), .Z(n1) );
  BUF_X1 U3 ( .A(SEL), .Z(n3) );
endmodule


module EXU_N32 ( DATA1, DATA2, FUNC, RD_in, SN, CLK, RST, OVF, stall_flag, 
        RD_sel_flag, OUTPUT, RD_stall, RD_out, H_MULOUT );
  input [31:0] DATA1;
  input [31:0] DATA2;
  input [3:0] FUNC;
  input [4:0] RD_in;
  output [31:0] OUTPUT;
  output [4:0] RD_stall;
  output [4:0] RD_out;
  output [31:0] H_MULOUT;
  input SN, CLK, RST;
  output OVF, stall_flag, RD_sel_flag;
  wire   mul_flag_reg1, N3, n1;
  wire   [4:0] RD_reg2;
  wire   [4:0] s_RD_in;
  wire   [31:0] s_ALUout;
  wire   [31:0] s_mul_out;

  DFFR_X1 \RD_reg1_reg[4]  ( .D(s_RD_in[4]), .CK(CLK), .RN(n1), .Q(RD_stall[4]) );
  DFFR_X1 \RD_reg1_reg[3]  ( .D(s_RD_in[3]), .CK(CLK), .RN(n1), .Q(RD_stall[3]) );
  DFFR_X1 \RD_reg1_reg[2]  ( .D(s_RD_in[2]), .CK(CLK), .RN(n1), .Q(RD_stall[2]) );
  DFFR_X1 \RD_reg1_reg[1]  ( .D(s_RD_in[1]), .CK(CLK), .RN(n1), .Q(RD_stall[1]) );
  DFFR_X1 \RD_reg1_reg[0]  ( .D(s_RD_in[0]), .CK(CLK), .RN(n1), .Q(RD_stall[0]) );
  DFFR_X1 \RD_reg2_reg[4]  ( .D(RD_stall[4]), .CK(CLK), .RN(n1), .Q(RD_reg2[4]) );
  DFFR_X1 \RD_reg2_reg[3]  ( .D(RD_stall[3]), .CK(CLK), .RN(n1), .Q(RD_reg2[3]) );
  DFFR_X1 \RD_reg2_reg[2]  ( .D(RD_stall[2]), .CK(CLK), .RN(n1), .Q(RD_reg2[2]) );
  DFFR_X1 \RD_reg2_reg[1]  ( .D(RD_stall[1]), .CK(CLK), .RN(n1), .Q(RD_reg2[1]) );
  DFFR_X1 \RD_reg2_reg[0]  ( .D(RD_stall[0]), .CK(CLK), .RN(n1), .Q(RD_reg2[0]) );
  DFFR_X1 \RD_reg3_reg[4]  ( .D(RD_reg2[4]), .CK(CLK), .RN(n1), .Q(RD_out[4])
         );
  DFFR_X1 \RD_reg3_reg[3]  ( .D(RD_reg2[3]), .CK(CLK), .RN(n1), .Q(RD_out[3])
         );
  DFFR_X1 \RD_reg3_reg[2]  ( .D(RD_reg2[2]), .CK(CLK), .RN(n1), .Q(RD_out[2])
         );
  DFFR_X1 \RD_reg3_reg[1]  ( .D(RD_reg2[1]), .CK(CLK), .RN(n1), .Q(RD_out[1])
         );
  DFFR_X1 \RD_reg3_reg[0]  ( .D(RD_reg2[0]), .CK(CLK), .RN(n1), .Q(RD_out[0])
         );
  DFFR_X1 mul_flag_reg1_reg ( .D(N3), .CK(CLK), .RN(n1), .Q(mul_flag_reg1) );
  DFFR_X1 mul_flag_reg2_reg ( .D(mul_flag_reg1), .CK(CLK), .RN(n1), .Q(
        stall_flag) );
  ALU_N32 ALU1 ( .DATA1(DATA1), .DATA2(DATA2), .FUNC(FUNC), .SN(SN), .OVF(OVF), 
        .OUTALU(s_ALUout) );
  boothmul_NBIT_in32 MUL ( .A(DATA1), .B(DATA2), .mulin_flag(N3), .CLK(CLK), 
        .RST(n1), .MULready(RD_sel_flag), .P({H_MULOUT, s_mul_out}) );
  MUX21_GENERIC_NBIT32_1 OUTPUT_MUX ( .A(s_ALUout), .B(s_mul_out), .SEL(
        RD_sel_flag), .Y(OUTPUT) );
  BUF_X1 U3 ( .A(RST), .Z(n1) );
  AND4_X1 U4 ( .A1(FUNC[3]), .A2(FUNC[2]), .A3(FUNC[1]), .A4(FUNC[0]), .ZN(N3)
         );
  AND2_X1 U5 ( .A1(RD_in[4]), .A2(N3), .ZN(s_RD_in[4]) );
  AND2_X1 U6 ( .A1(RD_in[2]), .A2(N3), .ZN(s_RD_in[2]) );
  AND2_X1 U7 ( .A1(RD_in[0]), .A2(N3), .ZN(s_RD_in[0]) );
  AND2_X1 U8 ( .A1(RD_in[1]), .A2(N3), .ZN(s_RD_in[1]) );
  AND2_X1 U9 ( .A1(RD_in[3]), .A2(N3), .ZN(s_RD_in[3]) );
endmodule


module MUX21_461 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_460 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_459 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_458 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_457 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_GENERIC_NBIT5_1 ( A, B, SEL, Y );
  input [4:0] A;
  input [4:0] B;
  output [4:0] Y;
  input SEL;


  MUX21_461 MUXES_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_460 MUXES_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_459 MUXES_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_458 MUXES_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
  MUX21_457 MUXES_4 ( .A(A[4]), .B(B[4]), .S(SEL), .Y(Y[4]) );
endmodule


module EXE ( CLK, RST, IMM, RA, RB, WA, RSA, RSB, ALU_outmem, WB_out, MEM_RD, 
        WB_RD, LD_EN, WB_EN, S1, S2, ALU3, ALU2, ALU1, ALU0, SN, RD_inmul, 
        flag_structHzd, flag_ismul, OVF, \output , ME, WAout );
  input [31:0] IMM;
  input [31:0] RA;
  input [31:0] RB;
  input [4:0] WA;
  input [4:0] RSA;
  input [4:0] RSB;
  input [31:0] ALU_outmem;
  input [31:0] WB_out;
  input [4:0] MEM_RD;
  input [4:0] WB_RD;
  output [4:0] RD_inmul;
  output [31:0] \output ;
  output [31:0] ME;
  output [4:0] WAout;
  input CLK, RST, LD_EN, WB_EN, S1, S2, ALU3, ALU2, ALU1, ALU0, SN;
  output flag_structHzd, flag_ismul, OVF;
  wire   N4, s_ovf, s_RD_sel2;
  wire   [1:0] s_S1;
  wire   [1:0] s_S2;
  wire   [1:0] s_S3;
  wire   [31:0] MUX1out;
  wire   [31:0] MUX2out;
  wire   [4:0] s_ALU_RD;
  wire   [4:0] s_mul_RD_out;
  assign flag_ismul = N4;

  forwarding_unit_WORD_size32_NREG32 FWU ( .RSA(RSA), .RSB(RSB), .ALU_outmem(
        ALU_outmem), .WB_out(WB_out), .MEM_RD(MEM_RD), .WB_RD(WB_RD), .LD_EN(
        LD_EN), .WB_EN(WB_EN), .S1(S1), .S2(S2), .SEL1(s_S1), .SEL2(s_S2), 
        .SEL3(s_S3) );
  MUX41_GENERIC_NBIT32_0 FW_MUX1 ( .A(IMM), .B(RA), .C(ALU_outmem), .D(WB_out), 
        .SEL(s_S1), .Y(MUX1out) );
  MUX41_GENERIC_NBIT32_2 FW_MUX2 ( .A(RB), .B(IMM), .C(ALU_outmem), .D(WB_out), 
        .SEL(s_S2), .Y(MUX2out) );
  MUX41_GENERIC_NBIT32_1 FW_MUX3 ( .A(IMM), .B(RB), .C(ALU_outmem), .D(WB_out), 
        .SEL(s_S3), .Y(ME) );
  MUX21_GENERIC_NBIT5_0 RD_MUX1 ( .A(WA), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
        .SEL(N4), .Y(s_ALU_RD) );
  EXU_N32 EXUx ( .DATA1(MUX1out), .DATA2(MUX2out), .FUNC({ALU3, ALU2, ALU1, 
        ALU0}), .RD_in(WA), .SN(SN), .CLK(CLK), .RST(RST), .OVF(s_ovf), 
        .stall_flag(flag_structHzd), .RD_sel_flag(s_RD_sel2), .OUTPUT(\output ), .RD_stall(RD_inmul), .RD_out(s_mul_RD_out) );
  MUX21_GENERIC_NBIT5_1 RD_MUX2 ( .A(s_ALU_RD), .B(s_mul_RD_out), .SEL(
        s_RD_sel2), .Y(WAout) );
  AND2_X1 U2 ( .A1(s_ovf), .A2(SN), .ZN(OVF) );
  AND4_X1 U3 ( .A1(ALU3), .A2(ALU2), .A3(ALU1), .A4(ALU0), .ZN(N4) );
endmodule


module MMU_WORD_size32 ( Wrd, BHU0, wdata_size );
  output [1:0] wdata_size;
  input Wrd, BHU0;
  wire   Wrd, N3;
  assign wdata_size[1] = Wrd;
  assign wdata_size[0] = N3;

  OR2_X1 U2 ( .A1(BHU0), .A2(Wrd), .ZN(N3) );
endmodule


module MUX51_0 ( A, B, C, D, E, S, Y );
  input [2:0] S;
  input A, B, C, D, E;
  output Y;
  wire   n5, n6, n7, n8, n1, n2, n3;

  AOI22_X1 U1 ( .A1(C), .A2(n1), .B1(D), .B2(S[0]), .ZN(n7) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S[0]), .B2(B), .ZN(n8) );
  INV_X1 U3 ( .A(n5), .ZN(Y) );
  AOI22_X1 U4 ( .A1(n6), .A2(n3), .B1(S[2]), .B2(E), .ZN(n5) );
  OAI22_X1 U5 ( .A1(n7), .A2(n2), .B1(S[1]), .B2(n8), .ZN(n6) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
  INV_X1 U8 ( .A(S[2]), .ZN(n3) );
endmodule


module MUX51_31 ( A, B, C, D, E, S, Y );
  input [2:0] S;
  input A, B, C, D, E;
  output Y;
  wire   n1, n2, n3, n9, n10, n11, n12;

  AOI22_X1 U1 ( .A1(A), .A2(n1), .B1(S[0]), .B2(B), .ZN(n9) );
  AOI22_X1 U2 ( .A1(C), .A2(n1), .B1(D), .B2(S[0]), .ZN(n10) );
  INV_X1 U3 ( .A(n12), .ZN(Y) );
  AOI22_X1 U4 ( .A1(n11), .A2(n3), .B1(S[2]), .B2(E), .ZN(n12) );
  OAI22_X1 U5 ( .A1(n10), .A2(n2), .B1(S[1]), .B2(n9), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
  INV_X1 U8 ( .A(S[2]), .ZN(n3) );
endmodule


module MUX51_30 ( A, B, C, D, E, S, Y );
  input [2:0] S;
  input A, B, C, D, E;
  output Y;
  wire   n1, n2, n3, n9, n10, n11, n12;

  AOI22_X1 U1 ( .A1(A), .A2(n1), .B1(S[0]), .B2(B), .ZN(n9) );
  AOI22_X1 U2 ( .A1(C), .A2(n1), .B1(D), .B2(S[0]), .ZN(n10) );
  INV_X1 U3 ( .A(n12), .ZN(Y) );
  AOI22_X1 U4 ( .A1(n11), .A2(n3), .B1(S[2]), .B2(E), .ZN(n12) );
  OAI22_X1 U5 ( .A1(n10), .A2(n2), .B1(S[1]), .B2(n9), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
  INV_X1 U8 ( .A(S[2]), .ZN(n3) );
endmodule


module MUX51_29 ( A, B, C, D, E, S, Y );
  input [2:0] S;
  input A, B, C, D, E;
  output Y;
  wire   n1, n2, n3, n9, n10, n11, n12;

  AOI22_X1 U1 ( .A1(A), .A2(n1), .B1(S[0]), .B2(B), .ZN(n9) );
  AOI22_X1 U2 ( .A1(C), .A2(n1), .B1(D), .B2(S[0]), .ZN(n10) );
  INV_X1 U3 ( .A(n12), .ZN(Y) );
  AOI22_X1 U4 ( .A1(n11), .A2(n3), .B1(S[2]), .B2(E), .ZN(n12) );
  OAI22_X1 U5 ( .A1(n10), .A2(n2), .B1(S[1]), .B2(n9), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
  INV_X1 U8 ( .A(S[2]), .ZN(n3) );
endmodule


module MUX51_28 ( A, B, C, D, E, S, Y );
  input [2:0] S;
  input A, B, C, D, E;
  output Y;
  wire   n1, n2, n3, n9, n10, n11, n12;

  AOI22_X1 U1 ( .A1(A), .A2(n1), .B1(S[0]), .B2(B), .ZN(n9) );
  AOI22_X1 U2 ( .A1(C), .A2(n1), .B1(D), .B2(S[0]), .ZN(n10) );
  INV_X1 U3 ( .A(n12), .ZN(Y) );
  AOI22_X1 U4 ( .A1(n11), .A2(n3), .B1(S[2]), .B2(E), .ZN(n12) );
  OAI22_X1 U5 ( .A1(n10), .A2(n2), .B1(S[1]), .B2(n9), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
  INV_X1 U8 ( .A(S[2]), .ZN(n3) );
endmodule


module MUX51_27 ( A, B, C, D, E, S, Y );
  input [2:0] S;
  input A, B, C, D, E;
  output Y;
  wire   n1, n2, n3, n9, n10, n11, n12;

  AOI22_X1 U1 ( .A1(A), .A2(n1), .B1(S[0]), .B2(B), .ZN(n9) );
  AOI22_X1 U2 ( .A1(C), .A2(n1), .B1(D), .B2(S[0]), .ZN(n10) );
  INV_X1 U3 ( .A(n12), .ZN(Y) );
  AOI22_X1 U4 ( .A1(n11), .A2(n3), .B1(S[2]), .B2(E), .ZN(n12) );
  OAI22_X1 U5 ( .A1(n10), .A2(n2), .B1(S[1]), .B2(n9), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
  INV_X1 U8 ( .A(S[2]), .ZN(n3) );
endmodule


module MUX51_26 ( A, B, C, D, E, S, Y );
  input [2:0] S;
  input A, B, C, D, E;
  output Y;
  wire   n1, n2, n3, n9, n10, n11, n12;

  AOI22_X1 U1 ( .A1(A), .A2(n1), .B1(S[0]), .B2(B), .ZN(n9) );
  AOI22_X1 U2 ( .A1(C), .A2(n1), .B1(D), .B2(S[0]), .ZN(n10) );
  INV_X1 U3 ( .A(n12), .ZN(Y) );
  AOI22_X1 U4 ( .A1(n11), .A2(n3), .B1(S[2]), .B2(E), .ZN(n12) );
  OAI22_X1 U5 ( .A1(n10), .A2(n2), .B1(S[1]), .B2(n9), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
  INV_X1 U8 ( .A(S[2]), .ZN(n3) );
endmodule


module MUX51_25 ( A, B, C, D, E, S, Y );
  input [2:0] S;
  input A, B, C, D, E;
  output Y;
  wire   n1, n2, n3, n9, n10, n11, n12;

  AOI22_X1 U1 ( .A1(A), .A2(n1), .B1(S[0]), .B2(B), .ZN(n9) );
  AOI22_X1 U2 ( .A1(C), .A2(n1), .B1(D), .B2(S[0]), .ZN(n10) );
  INV_X1 U3 ( .A(n12), .ZN(Y) );
  AOI22_X1 U4 ( .A1(n11), .A2(n3), .B1(S[2]), .B2(E), .ZN(n12) );
  OAI22_X1 U5 ( .A1(n10), .A2(n2), .B1(S[1]), .B2(n9), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
  INV_X1 U8 ( .A(S[2]), .ZN(n3) );
endmodule


module MUX51_24 ( A, B, C, D, E, S, Y );
  input [2:0] S;
  input A, B, C, D, E;
  output Y;
  wire   n1, n2, n3, n9, n10, n11, n12;

  AOI22_X1 U1 ( .A1(C), .A2(n1), .B1(D), .B2(S[0]), .ZN(n10) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S[0]), .B2(B), .ZN(n9) );
  INV_X1 U3 ( .A(n12), .ZN(Y) );
  AOI22_X1 U4 ( .A1(n11), .A2(n3), .B1(S[2]), .B2(E), .ZN(n12) );
  OAI22_X1 U5 ( .A1(n10), .A2(n2), .B1(S[1]), .B2(n9), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
  INV_X1 U8 ( .A(S[2]), .ZN(n3) );
endmodule


module MUX51_23 ( A, B, C, D, E, S, Y );
  input [2:0] S;
  input A, B, C, D, E;
  output Y;
  wire   n1, n2, n3, n9, n10, n11, n12;

  AOI22_X1 U1 ( .A1(C), .A2(n1), .B1(D), .B2(S[0]), .ZN(n10) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S[0]), .B2(B), .ZN(n9) );
  INV_X1 U3 ( .A(n12), .ZN(Y) );
  AOI22_X1 U4 ( .A1(n11), .A2(n3), .B1(S[2]), .B2(E), .ZN(n12) );
  OAI22_X1 U5 ( .A1(n10), .A2(n2), .B1(S[1]), .B2(n9), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
  INV_X1 U8 ( .A(S[2]), .ZN(n3) );
endmodule


module MUX51_22 ( A, B, C, D, E, S, Y );
  input [2:0] S;
  input A, B, C, D, E;
  output Y;
  wire   n1, n2, n3, n9, n10, n11, n12;

  AOI22_X1 U1 ( .A1(C), .A2(n1), .B1(D), .B2(S[0]), .ZN(n10) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S[0]), .B2(B), .ZN(n9) );
  INV_X1 U3 ( .A(n12), .ZN(Y) );
  AOI22_X1 U4 ( .A1(n11), .A2(n3), .B1(S[2]), .B2(E), .ZN(n12) );
  OAI22_X1 U5 ( .A1(n10), .A2(n2), .B1(S[1]), .B2(n9), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
  INV_X1 U8 ( .A(S[2]), .ZN(n3) );
endmodule


module MUX51_21 ( A, B, C, D, E, S, Y );
  input [2:0] S;
  input A, B, C, D, E;
  output Y;
  wire   n1, n2, n3, n9, n10, n11, n12;

  AOI22_X1 U1 ( .A1(C), .A2(n1), .B1(D), .B2(S[0]), .ZN(n10) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S[0]), .B2(B), .ZN(n9) );
  INV_X1 U3 ( .A(n12), .ZN(Y) );
  AOI22_X1 U4 ( .A1(n11), .A2(n3), .B1(S[2]), .B2(E), .ZN(n12) );
  OAI22_X1 U5 ( .A1(n10), .A2(n2), .B1(S[1]), .B2(n9), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
  INV_X1 U8 ( .A(S[2]), .ZN(n3) );
endmodule


module MUX51_20 ( A, B, C, D, E, S, Y );
  input [2:0] S;
  input A, B, C, D, E;
  output Y;
  wire   n1, n2, n3, n9, n10, n11, n12;

  AOI22_X1 U1 ( .A1(C), .A2(n1), .B1(D), .B2(S[0]), .ZN(n10) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S[0]), .B2(B), .ZN(n9) );
  INV_X1 U3 ( .A(n12), .ZN(Y) );
  AOI22_X1 U4 ( .A1(n11), .A2(n3), .B1(S[2]), .B2(E), .ZN(n12) );
  OAI22_X1 U5 ( .A1(n10), .A2(n2), .B1(S[1]), .B2(n9), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
  INV_X1 U8 ( .A(S[2]), .ZN(n3) );
endmodule


module MUX51_19 ( A, B, C, D, E, S, Y );
  input [2:0] S;
  input A, B, C, D, E;
  output Y;
  wire   n1, n2, n3, n9, n10, n11, n12;

  AOI22_X1 U1 ( .A1(C), .A2(n1), .B1(D), .B2(S[0]), .ZN(n10) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S[0]), .B2(B), .ZN(n9) );
  INV_X1 U3 ( .A(n12), .ZN(Y) );
  AOI22_X1 U4 ( .A1(n11), .A2(n3), .B1(S[2]), .B2(E), .ZN(n12) );
  OAI22_X1 U5 ( .A1(n10), .A2(n2), .B1(S[1]), .B2(n9), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
  INV_X1 U8 ( .A(S[2]), .ZN(n3) );
endmodule


module MUX51_18 ( A, B, C, D, E, S, Y );
  input [2:0] S;
  input A, B, C, D, E;
  output Y;
  wire   n1, n2, n3, n9, n10, n11, n12;

  AOI22_X1 U1 ( .A1(C), .A2(n1), .B1(D), .B2(S[0]), .ZN(n10) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S[0]), .B2(B), .ZN(n9) );
  INV_X1 U3 ( .A(n12), .ZN(Y) );
  AOI22_X1 U4 ( .A1(n11), .A2(n3), .B1(S[2]), .B2(E), .ZN(n12) );
  OAI22_X1 U5 ( .A1(n10), .A2(n2), .B1(S[1]), .B2(n9), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
  INV_X1 U8 ( .A(S[2]), .ZN(n3) );
endmodule


module MUX51_17 ( A, B, C, D, E, S, Y );
  input [2:0] S;
  input A, B, C, D, E;
  output Y;
  wire   n1, n2, n3, n9, n10, n11, n12;

  AOI22_X1 U1 ( .A1(C), .A2(n1), .B1(D), .B2(S[0]), .ZN(n10) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S[0]), .B2(B), .ZN(n9) );
  INV_X1 U3 ( .A(n12), .ZN(Y) );
  AOI22_X1 U4 ( .A1(n11), .A2(n3), .B1(S[2]), .B2(E), .ZN(n12) );
  OAI22_X1 U5 ( .A1(n10), .A2(n2), .B1(S[1]), .B2(n9), .ZN(n11) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
  INV_X1 U8 ( .A(S[2]), .ZN(n3) );
endmodule


module MUX51_16 ( A, B, C, D, E, S, Y );
  input [2:0] S;
  input A, B, C, D, E;
  output Y;
  wire   n1, n2, n3, n9, n10, n11, n12;

  AOI22_X1 U1 ( .A1(C), .A2(n1), .B1(D), .B2(S[0]), .ZN(n10) );
  INV_X1 U2 ( .A(n12), .ZN(Y) );
  AOI22_X1 U3 ( .A1(n11), .A2(n3), .B1(S[2]), .B2(E), .ZN(n12) );
  OAI22_X1 U4 ( .A1(n10), .A2(n2), .B1(S[1]), .B2(n9), .ZN(n11) );
  AOI22_X1 U5 ( .A1(A), .A2(n1), .B1(S[0]), .B2(B), .ZN(n9) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
  INV_X1 U8 ( .A(S[2]), .ZN(n3) );
endmodule


module MUX51_15 ( A, B, C, D, E, S, Y );
  input [2:0] S;
  input A, B, C, D, E;
  output Y;
  wire   n1, n2, n3, n9, n10, n11, n12;

  AOI22_X1 U1 ( .A1(C), .A2(n1), .B1(D), .B2(S[0]), .ZN(n10) );
  INV_X1 U2 ( .A(n12), .ZN(Y) );
  AOI22_X1 U3 ( .A1(n11), .A2(n3), .B1(S[2]), .B2(E), .ZN(n12) );
  OAI22_X1 U4 ( .A1(n10), .A2(n2), .B1(S[1]), .B2(n9), .ZN(n11) );
  AOI22_X1 U5 ( .A1(A), .A2(n1), .B1(S[0]), .B2(B), .ZN(n9) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
  INV_X1 U8 ( .A(S[2]), .ZN(n3) );
endmodule


module MUX51_14 ( A, B, C, D, E, S, Y );
  input [2:0] S;
  input A, B, C, D, E;
  output Y;
  wire   n1, n2, n3, n9, n10, n11, n12;

  AOI22_X1 U1 ( .A1(C), .A2(n1), .B1(D), .B2(S[0]), .ZN(n10) );
  INV_X1 U2 ( .A(n12), .ZN(Y) );
  AOI22_X1 U3 ( .A1(n11), .A2(n3), .B1(S[2]), .B2(E), .ZN(n12) );
  OAI22_X1 U4 ( .A1(n10), .A2(n2), .B1(S[1]), .B2(n9), .ZN(n11) );
  AOI22_X1 U5 ( .A1(A), .A2(n1), .B1(S[0]), .B2(B), .ZN(n9) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
  INV_X1 U8 ( .A(S[2]), .ZN(n3) );
endmodule


module MUX51_13 ( A, B, C, D, E, S, Y );
  input [2:0] S;
  input A, B, C, D, E;
  output Y;
  wire   n1, n2, n3, n9, n10, n11, n12;

  AOI22_X1 U1 ( .A1(C), .A2(n1), .B1(D), .B2(S[0]), .ZN(n10) );
  INV_X1 U2 ( .A(n12), .ZN(Y) );
  AOI22_X1 U3 ( .A1(n11), .A2(n3), .B1(S[2]), .B2(E), .ZN(n12) );
  OAI22_X1 U4 ( .A1(n10), .A2(n2), .B1(S[1]), .B2(n9), .ZN(n11) );
  AOI22_X1 U5 ( .A1(A), .A2(n1), .B1(S[0]), .B2(B), .ZN(n9) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
  INV_X1 U8 ( .A(S[2]), .ZN(n3) );
endmodule


module MUX51_12 ( A, B, C, D, E, S, Y );
  input [2:0] S;
  input A, B, C, D, E;
  output Y;
  wire   n1, n2, n3, n9, n10, n11, n12;

  AOI22_X1 U1 ( .A1(C), .A2(n1), .B1(D), .B2(S[0]), .ZN(n10) );
  INV_X1 U2 ( .A(n12), .ZN(Y) );
  AOI22_X1 U3 ( .A1(n11), .A2(n3), .B1(S[2]), .B2(E), .ZN(n12) );
  OAI22_X1 U4 ( .A1(n10), .A2(n2), .B1(S[1]), .B2(n9), .ZN(n11) );
  AOI22_X1 U5 ( .A1(A), .A2(n1), .B1(S[0]), .B2(B), .ZN(n9) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
  INV_X1 U8 ( .A(S[2]), .ZN(n3) );
endmodule


module MUX51_11 ( A, B, C, D, E, S, Y );
  input [2:0] S;
  input A, B, C, D, E;
  output Y;
  wire   n1, n2, n3, n9, n10, n11, n12;

  AOI22_X1 U1 ( .A1(C), .A2(n1), .B1(D), .B2(S[0]), .ZN(n10) );
  INV_X1 U2 ( .A(n12), .ZN(Y) );
  AOI22_X1 U3 ( .A1(n11), .A2(n3), .B1(S[2]), .B2(E), .ZN(n12) );
  OAI22_X1 U4 ( .A1(n10), .A2(n2), .B1(S[1]), .B2(n9), .ZN(n11) );
  AOI22_X1 U5 ( .A1(A), .A2(n1), .B1(S[0]), .B2(B), .ZN(n9) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
  INV_X1 U8 ( .A(S[2]), .ZN(n3) );
endmodule


module MUX51_10 ( A, B, C, D, E, S, Y );
  input [2:0] S;
  input A, B, C, D, E;
  output Y;
  wire   n1, n2, n3, n9, n10, n11, n12;

  AOI22_X1 U1 ( .A1(C), .A2(n1), .B1(D), .B2(S[0]), .ZN(n10) );
  INV_X1 U2 ( .A(n12), .ZN(Y) );
  AOI22_X1 U3 ( .A1(n11), .A2(n3), .B1(S[2]), .B2(E), .ZN(n12) );
  OAI22_X1 U4 ( .A1(n10), .A2(n2), .B1(S[1]), .B2(n9), .ZN(n11) );
  AOI22_X1 U5 ( .A1(A), .A2(n1), .B1(S[0]), .B2(B), .ZN(n9) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
  INV_X1 U8 ( .A(S[2]), .ZN(n3) );
endmodule


module MUX51_9 ( A, B, C, D, E, S, Y );
  input [2:0] S;
  input A, B, C, D, E;
  output Y;
  wire   n1, n2, n3, n9, n10, n11, n12;

  AOI22_X1 U1 ( .A1(C), .A2(n1), .B1(D), .B2(S[0]), .ZN(n10) );
  INV_X1 U2 ( .A(n12), .ZN(Y) );
  AOI22_X1 U3 ( .A1(n11), .A2(n3), .B1(S[2]), .B2(E), .ZN(n12) );
  OAI22_X1 U4 ( .A1(n10), .A2(n2), .B1(S[1]), .B2(n9), .ZN(n11) );
  AOI22_X1 U5 ( .A1(A), .A2(n1), .B1(S[0]), .B2(B), .ZN(n9) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
  INV_X1 U8 ( .A(S[2]), .ZN(n3) );
endmodule


module MUX51_8 ( A, B, C, D, E, S, Y );
  input [2:0] S;
  input A, B, C, D, E;
  output Y;
  wire   n1, n2, n3, n9, n10, n11, n12;

  AOI22_X1 U1 ( .A1(C), .A2(n1), .B1(D), .B2(S[0]), .ZN(n10) );
  INV_X1 U2 ( .A(n12), .ZN(Y) );
  AOI22_X1 U3 ( .A1(n11), .A2(n3), .B1(S[2]), .B2(E), .ZN(n12) );
  OAI22_X1 U4 ( .A1(n10), .A2(n2), .B1(S[1]), .B2(n9), .ZN(n11) );
  AOI22_X1 U5 ( .A1(A), .A2(n1), .B1(S[0]), .B2(B), .ZN(n9) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
  INV_X1 U8 ( .A(S[2]), .ZN(n3) );
endmodule


module MUX51_7 ( A, B, C, D, E, S, Y );
  input [2:0] S;
  input A, B, C, D, E;
  output Y;
  wire   n1, n2, n3, n9, n10, n11, n12;

  AOI22_X1 U1 ( .A1(C), .A2(n1), .B1(D), .B2(S[0]), .ZN(n10) );
  INV_X1 U2 ( .A(n12), .ZN(Y) );
  AOI22_X1 U3 ( .A1(n11), .A2(n3), .B1(S[2]), .B2(E), .ZN(n12) );
  OAI22_X1 U4 ( .A1(n10), .A2(n2), .B1(S[1]), .B2(n9), .ZN(n11) );
  AOI22_X1 U5 ( .A1(A), .A2(n1), .B1(S[0]), .B2(B), .ZN(n9) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
  INV_X1 U8 ( .A(S[2]), .ZN(n3) );
endmodule


module MUX51_6 ( A, B, C, D, E, S, Y );
  input [2:0] S;
  input A, B, C, D, E;
  output Y;
  wire   n1, n2, n3, n9, n10, n11, n12;

  AOI22_X1 U1 ( .A1(C), .A2(n1), .B1(D), .B2(S[0]), .ZN(n10) );
  INV_X1 U2 ( .A(n12), .ZN(Y) );
  AOI22_X1 U3 ( .A1(n11), .A2(n3), .B1(S[2]), .B2(E), .ZN(n12) );
  OAI22_X1 U4 ( .A1(n10), .A2(n2), .B1(S[1]), .B2(n9), .ZN(n11) );
  AOI22_X1 U5 ( .A1(A), .A2(n1), .B1(S[0]), .B2(B), .ZN(n9) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
  INV_X1 U8 ( .A(S[2]), .ZN(n3) );
endmodule


module MUX51_5 ( A, B, C, D, E, S, Y );
  input [2:0] S;
  input A, B, C, D, E;
  output Y;
  wire   n1, n2, n3, n9, n10, n11, n12;

  AOI22_X1 U1 ( .A1(C), .A2(n1), .B1(D), .B2(S[0]), .ZN(n10) );
  INV_X1 U2 ( .A(n12), .ZN(Y) );
  AOI22_X1 U3 ( .A1(n11), .A2(n3), .B1(S[2]), .B2(E), .ZN(n12) );
  OAI22_X1 U4 ( .A1(n10), .A2(n2), .B1(S[1]), .B2(n9), .ZN(n11) );
  AOI22_X1 U5 ( .A1(A), .A2(n1), .B1(S[0]), .B2(B), .ZN(n9) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
  INV_X1 U8 ( .A(S[2]), .ZN(n3) );
endmodule


module MUX51_4 ( A, B, C, D, E, S, Y );
  input [2:0] S;
  input A, B, C, D, E;
  output Y;
  wire   n1, n2, n3, n9, n10, n11, n12;

  AOI22_X1 U1 ( .A1(C), .A2(n1), .B1(D), .B2(S[0]), .ZN(n10) );
  INV_X1 U2 ( .A(n12), .ZN(Y) );
  AOI22_X1 U3 ( .A1(n11), .A2(n3), .B1(S[2]), .B2(E), .ZN(n12) );
  OAI22_X1 U4 ( .A1(n10), .A2(n2), .B1(S[1]), .B2(n9), .ZN(n11) );
  AOI22_X1 U5 ( .A1(A), .A2(n1), .B1(S[0]), .B2(B), .ZN(n9) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
  INV_X1 U8 ( .A(S[2]), .ZN(n3) );
endmodule


module MUX51_3 ( A, B, C, D, E, S, Y );
  input [2:0] S;
  input A, B, C, D, E;
  output Y;
  wire   n1, n2, n3, n9, n10, n11, n12;

  AOI22_X1 U1 ( .A1(C), .A2(n1), .B1(D), .B2(S[0]), .ZN(n10) );
  INV_X1 U2 ( .A(n12), .ZN(Y) );
  AOI22_X1 U3 ( .A1(n11), .A2(n3), .B1(S[2]), .B2(E), .ZN(n12) );
  OAI22_X1 U4 ( .A1(n10), .A2(n2), .B1(S[1]), .B2(n9), .ZN(n11) );
  AOI22_X1 U5 ( .A1(A), .A2(n1), .B1(S[0]), .B2(B), .ZN(n9) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
  INV_X1 U8 ( .A(S[2]), .ZN(n3) );
endmodule


module MUX51_2 ( A, B, C, D, E, S, Y );
  input [2:0] S;
  input A, B, C, D, E;
  output Y;
  wire   n1, n2, n3, n9, n10, n11, n12;

  AOI22_X1 U1 ( .A1(C), .A2(n1), .B1(D), .B2(S[0]), .ZN(n10) );
  INV_X1 U2 ( .A(n12), .ZN(Y) );
  AOI22_X1 U3 ( .A1(n11), .A2(n3), .B1(S[2]), .B2(E), .ZN(n12) );
  OAI22_X1 U4 ( .A1(n10), .A2(n2), .B1(S[1]), .B2(n9), .ZN(n11) );
  AOI22_X1 U5 ( .A1(A), .A2(n1), .B1(S[0]), .B2(B), .ZN(n9) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
  INV_X1 U8 ( .A(S[2]), .ZN(n3) );
endmodule


module MUX51_1 ( A, B, C, D, E, S, Y );
  input [2:0] S;
  input A, B, C, D, E;
  output Y;
  wire   n1, n2, n3, n9, n10, n11, n12;

  AOI22_X1 U1 ( .A1(C), .A2(n1), .B1(D), .B2(S[0]), .ZN(n10) );
  INV_X1 U2 ( .A(n12), .ZN(Y) );
  AOI22_X1 U3 ( .A1(n11), .A2(n3), .B1(S[2]), .B2(E), .ZN(n12) );
  OAI22_X1 U4 ( .A1(n10), .A2(n2), .B1(S[1]), .B2(n9), .ZN(n11) );
  AOI22_X1 U5 ( .A1(A), .A2(n1), .B1(S[0]), .B2(B), .ZN(n9) );
  INV_X1 U6 ( .A(S[0]), .ZN(n1) );
  INV_X1 U7 ( .A(S[1]), .ZN(n2) );
  INV_X1 U8 ( .A(S[2]), .ZN(n3) );
endmodule


module MUX51_GENERIC_NBIT32 ( A, B, C, D, E, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [31:0] D;
  input [31:0] E;
  input [2:0] SEL;
  output [31:0] Y;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9;

  MUX51_0 MUXES_0 ( .A(A[0]), .B(B[0]), .C(C[0]), .D(D[0]), .E(E[0]), .S({n9, 
        n6, n3}), .Y(Y[0]) );
  MUX51_31 MUXES_1 ( .A(A[1]), .B(B[1]), .C(C[1]), .D(D[1]), .E(E[1]), .S({n7, 
        n4, n1}), .Y(Y[1]) );
  MUX51_30 MUXES_2 ( .A(A[2]), .B(B[2]), .C(C[2]), .D(D[2]), .E(E[2]), .S({n7, 
        n4, n1}), .Y(Y[2]) );
  MUX51_29 MUXES_3 ( .A(A[3]), .B(B[3]), .C(C[3]), .D(D[3]), .E(E[3]), .S({n7, 
        n4, n1}), .Y(Y[3]) );
  MUX51_28 MUXES_4 ( .A(A[4]), .B(B[4]), .C(C[4]), .D(D[4]), .E(E[4]), .S({n7, 
        n4, n1}), .Y(Y[4]) );
  MUX51_27 MUXES_5 ( .A(A[5]), .B(B[5]), .C(C[5]), .D(D[5]), .E(E[5]), .S({n7, 
        n4, n1}), .Y(Y[5]) );
  MUX51_26 MUXES_6 ( .A(A[6]), .B(B[6]), .C(C[6]), .D(D[6]), .E(E[6]), .S({n7, 
        n4, n1}), .Y(Y[6]) );
  MUX51_25 MUXES_7 ( .A(A[7]), .B(B[7]), .C(C[7]), .D(D[7]), .E(E[7]), .S({n7, 
        n4, n1}), .Y(Y[7]) );
  MUX51_24 MUXES_8 ( .A(A[8]), .B(B[8]), .C(C[8]), .D(D[8]), .E(E[8]), .S({n7, 
        n4, n1}), .Y(Y[8]) );
  MUX51_23 MUXES_9 ( .A(A[9]), .B(B[9]), .C(C[9]), .D(D[9]), .E(E[9]), .S({n7, 
        n4, n1}), .Y(Y[9]) );
  MUX51_22 MUXES_10 ( .A(A[10]), .B(B[10]), .C(C[10]), .D(D[10]), .E(E[10]), 
        .S({n7, n4, n1}), .Y(Y[10]) );
  MUX51_21 MUXES_11 ( .A(A[11]), .B(B[11]), .C(C[11]), .D(D[11]), .E(E[11]), 
        .S({n7, n4, n1}), .Y(Y[11]) );
  MUX51_20 MUXES_12 ( .A(A[12]), .B(B[12]), .C(C[12]), .D(D[12]), .E(E[12]), 
        .S({n7, n4, n1}), .Y(Y[12]) );
  MUX51_19 MUXES_13 ( .A(A[13]), .B(B[13]), .C(C[13]), .D(D[13]), .E(E[13]), 
        .S({n8, n5, n2}), .Y(Y[13]) );
  MUX51_18 MUXES_14 ( .A(A[14]), .B(B[14]), .C(C[14]), .D(D[14]), .E(E[14]), 
        .S({n8, n5, n2}), .Y(Y[14]) );
  MUX51_17 MUXES_15 ( .A(A[15]), .B(B[15]), .C(C[15]), .D(D[15]), .E(E[15]), 
        .S({n8, n5, n2}), .Y(Y[15]) );
  MUX51_16 MUXES_16 ( .A(A[16]), .B(B[16]), .C(C[16]), .D(D[16]), .E(E[16]), 
        .S({n8, n5, n2}), .Y(Y[16]) );
  MUX51_15 MUXES_17 ( .A(A[17]), .B(B[17]), .C(C[17]), .D(D[17]), .E(E[17]), 
        .S({n8, n5, n2}), .Y(Y[17]) );
  MUX51_14 MUXES_18 ( .A(A[18]), .B(B[18]), .C(C[18]), .D(D[18]), .E(E[18]), 
        .S({n8, n5, n2}), .Y(Y[18]) );
  MUX51_13 MUXES_19 ( .A(A[19]), .B(B[19]), .C(C[19]), .D(D[19]), .E(E[19]), 
        .S({n8, n5, n2}), .Y(Y[19]) );
  MUX51_12 MUXES_20 ( .A(A[20]), .B(B[20]), .C(C[20]), .D(D[20]), .E(E[20]), 
        .S({n8, n5, n2}), .Y(Y[20]) );
  MUX51_11 MUXES_21 ( .A(A[21]), .B(B[21]), .C(C[21]), .D(D[21]), .E(E[21]), 
        .S({n8, n5, n2}), .Y(Y[21]) );
  MUX51_10 MUXES_22 ( .A(A[22]), .B(B[22]), .C(C[22]), .D(D[22]), .E(E[22]), 
        .S({n8, n5, n2}), .Y(Y[22]) );
  MUX51_9 MUXES_23 ( .A(A[23]), .B(B[23]), .C(C[23]), .D(D[23]), .E(E[23]), 
        .S({n8, n5, n2}), .Y(Y[23]) );
  MUX51_8 MUXES_24 ( .A(A[24]), .B(B[24]), .C(C[24]), .D(D[24]), .E(E[24]), 
        .S({n8, n5, n2}), .Y(Y[24]) );
  MUX51_7 MUXES_25 ( .A(A[25]), .B(B[25]), .C(C[25]), .D(D[25]), .E(E[25]), 
        .S({n9, n6, n3}), .Y(Y[25]) );
  MUX51_6 MUXES_26 ( .A(A[26]), .B(B[26]), .C(C[26]), .D(D[26]), .E(E[26]), 
        .S({n9, n6, n3}), .Y(Y[26]) );
  MUX51_5 MUXES_27 ( .A(A[27]), .B(B[27]), .C(C[27]), .D(D[27]), .E(E[27]), 
        .S({n9, n6, n3}), .Y(Y[27]) );
  MUX51_4 MUXES_28 ( .A(A[28]), .B(B[28]), .C(C[28]), .D(D[28]), .E(E[28]), 
        .S({n9, n6, n3}), .Y(Y[28]) );
  MUX51_3 MUXES_29 ( .A(A[29]), .B(B[29]), .C(C[29]), .D(D[29]), .E(E[29]), 
        .S({n9, n6, n3}), .Y(Y[29]) );
  MUX51_2 MUXES_30 ( .A(A[30]), .B(B[30]), .C(C[30]), .D(D[30]), .E(E[30]), 
        .S({n9, n6, n3}), .Y(Y[30]) );
  MUX51_1 MUXES_31 ( .A(A[31]), .B(B[31]), .C(C[31]), .D(D[31]), .E(E[31]), 
        .S({n9, n6, n3}), .Y(Y[31]) );
  BUF_X1 U1 ( .A(SEL[0]), .Z(n3) );
  BUF_X2 U2 ( .A(SEL[0]), .Z(n2) );
  BUF_X2 U3 ( .A(SEL[0]), .Z(n1) );
  BUF_X1 U4 ( .A(SEL[1]), .Z(n5) );
  BUF_X1 U5 ( .A(SEL[1]), .Z(n4) );
  BUF_X1 U6 ( .A(SEL[2]), .Z(n8) );
  BUF_X1 U7 ( .A(SEL[2]), .Z(n7) );
  BUF_X1 U8 ( .A(SEL[1]), .Z(n6) );
  BUF_X1 U9 ( .A(SEL[2]), .Z(n9) );
endmodule


module MEM_MEMORY_SIZE128 ( CLK, RST, ALUout, MEout, RDin, DRAM_data_out, LnS, 
        Wrd, BHU1, BHU0, EN3, DRAM_addr, DRAM_data_in, MMU_out, \output , 
        alu_out, RDout );
  input [31:0] ALUout;
  input [31:0] MEout;
  input [4:0] RDin;
  input [31:0] DRAM_data_out;
  output [8:0] DRAM_addr;
  output [31:0] DRAM_data_in;
  output [1:0] MMU_out;
  output [31:0] \output ;
  output [31:0] alu_out;
  output [4:0] RDout;
  input CLK, RST, LnS, Wrd, BHU1, BHU0, EN3;
  wire   n1, n2, n3, n4, n5, n6;
  assign DRAM_data_in[31] = MEout[31];
  assign DRAM_data_in[30] = MEout[30];
  assign DRAM_data_in[29] = MEout[29];
  assign DRAM_data_in[28] = MEout[28];
  assign DRAM_data_in[27] = MEout[27];
  assign DRAM_data_in[26] = MEout[26];
  assign DRAM_data_in[25] = MEout[25];
  assign DRAM_data_in[24] = MEout[24];
  assign DRAM_data_in[23] = MEout[23];
  assign DRAM_data_in[22] = MEout[22];
  assign DRAM_data_in[21] = MEout[21];
  assign DRAM_data_in[20] = MEout[20];
  assign DRAM_data_in[19] = MEout[19];
  assign DRAM_data_in[18] = MEout[18];
  assign DRAM_data_in[17] = MEout[17];
  assign DRAM_data_in[16] = MEout[16];
  assign DRAM_data_in[15] = MEout[15];
  assign DRAM_data_in[14] = MEout[14];
  assign DRAM_data_in[13] = MEout[13];
  assign DRAM_data_in[12] = MEout[12];
  assign DRAM_data_in[11] = MEout[11];
  assign DRAM_data_in[10] = MEout[10];
  assign DRAM_data_in[9] = MEout[9];
  assign DRAM_data_in[8] = MEout[8];
  assign DRAM_data_in[7] = MEout[7];
  assign DRAM_data_in[6] = MEout[6];
  assign DRAM_data_in[5] = MEout[5];
  assign DRAM_data_in[4] = MEout[4];
  assign DRAM_data_in[3] = MEout[3];
  assign DRAM_data_in[2] = MEout[2];
  assign DRAM_data_in[1] = MEout[1];
  assign DRAM_data_in[0] = MEout[0];
  assign alu_out[31] = ALUout[31];
  assign alu_out[30] = ALUout[30];
  assign alu_out[29] = ALUout[29];
  assign alu_out[28] = ALUout[28];
  assign alu_out[27] = ALUout[27];
  assign alu_out[26] = ALUout[26];
  assign alu_out[25] = ALUout[25];
  assign alu_out[24] = ALUout[24];
  assign alu_out[23] = ALUout[23];
  assign alu_out[22] = ALUout[22];
  assign alu_out[21] = ALUout[21];
  assign alu_out[20] = ALUout[20];
  assign alu_out[19] = ALUout[19];
  assign alu_out[18] = ALUout[18];
  assign alu_out[17] = ALUout[17];
  assign alu_out[16] = ALUout[16];
  assign alu_out[15] = ALUout[15];
  assign alu_out[14] = ALUout[14];
  assign alu_out[13] = ALUout[13];
  assign alu_out[12] = ALUout[12];
  assign alu_out[11] = ALUout[11];
  assign alu_out[10] = ALUout[10];
  assign alu_out[9] = ALUout[9];
  assign alu_out[8] = ALUout[8];
  assign DRAM_addr[8] = ALUout[8];
  assign alu_out[7] = ALUout[7];
  assign DRAM_addr[7] = ALUout[7];
  assign alu_out[6] = ALUout[6];
  assign DRAM_addr[6] = ALUout[6];
  assign alu_out[5] = ALUout[5];
  assign DRAM_addr[5] = ALUout[5];
  assign alu_out[4] = ALUout[4];
  assign DRAM_addr[4] = ALUout[4];
  assign alu_out[3] = ALUout[3];
  assign DRAM_addr[3] = ALUout[3];
  assign alu_out[2] = ALUout[2];
  assign DRAM_addr[2] = ALUout[2];
  assign alu_out[1] = ALUout[1];
  assign DRAM_addr[1] = ALUout[1];
  assign alu_out[0] = ALUout[0];
  assign DRAM_addr[0] = ALUout[0];
  assign RDout[4] = RDin[4];
  assign RDout[3] = RDin[3];
  assign RDout[2] = RDin[2];
  assign RDout[1] = RDin[1];
  assign RDout[0] = RDin[0];

  MMU_WORD_size32 mem_MU ( .Wrd(Wrd), .BHU0(BHU0), .wdata_size(MMU_out) );
  MUX51_GENERIC_NBIT32 mux ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, n4, DRAM_data_out[30:24]}), .B({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, n3, DRAM_data_out[30:16]}), .C({n3, n3, n3, n3, n3, 
        n3, n3, n3, n3, n3, n4, n4, n4, n4, n4, n4, n4, n4, n4, n4, n4, n5, n5, 
        n5, n5, DRAM_data_out[30:24]}), .D({n5, n5, n5, n5, n5, n5, n5, n5, n5, 
        n6, n6, n6, n6, n6, n6, n6, n6, DRAM_data_out[30:16]}), .E({n3, 
        DRAM_data_out[30:0]}), .SEL({Wrd, BHU1, BHU0}), .Y(\output ) );
  BUF_X1 U2 ( .A(n2), .Z(n5) );
  BUF_X1 U3 ( .A(n1), .Z(n3) );
  BUF_X1 U4 ( .A(n1), .Z(n4) );
  BUF_X1 U5 ( .A(n2), .Z(n6) );
  BUF_X1 U6 ( .A(DRAM_data_out[31]), .Z(n1) );
  BUF_X1 U7 ( .A(DRAM_data_out[31]), .Z(n2) );
endmodule


module MUX21_456 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_455 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_454 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_453 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_452 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_451 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_450 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_449 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_448 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_447 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_446 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_445 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_444 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_443 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_442 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_441 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_440 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_439 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_438 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_437 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_436 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_435 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_434 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_433 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_432 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_431 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_430 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_429 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_428 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_427 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_426 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_425 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n4;

  INV_X1 U1 ( .A(n4), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n4) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_GENERIC_NBIT32_2 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   n1, n2, n3;

  MUX21_456 MUXES_0 ( .A(A[0]), .B(B[0]), .S(n1), .Y(Y[0]) );
  MUX21_455 MUXES_1 ( .A(A[1]), .B(B[1]), .S(n1), .Y(Y[1]) );
  MUX21_454 MUXES_2 ( .A(A[2]), .B(B[2]), .S(n1), .Y(Y[2]) );
  MUX21_453 MUXES_3 ( .A(A[3]), .B(B[3]), .S(n1), .Y(Y[3]) );
  MUX21_452 MUXES_4 ( .A(A[4]), .B(B[4]), .S(n1), .Y(Y[4]) );
  MUX21_451 MUXES_5 ( .A(A[5]), .B(B[5]), .S(n1), .Y(Y[5]) );
  MUX21_450 MUXES_6 ( .A(A[6]), .B(B[6]), .S(n1), .Y(Y[6]) );
  MUX21_449 MUXES_7 ( .A(A[7]), .B(B[7]), .S(n1), .Y(Y[7]) );
  MUX21_448 MUXES_8 ( .A(A[8]), .B(B[8]), .S(n1), .Y(Y[8]) );
  MUX21_447 MUXES_9 ( .A(A[9]), .B(B[9]), .S(n1), .Y(Y[9]) );
  MUX21_446 MUXES_10 ( .A(A[10]), .B(B[10]), .S(n1), .Y(Y[10]) );
  MUX21_445 MUXES_11 ( .A(A[11]), .B(B[11]), .S(n1), .Y(Y[11]) );
  MUX21_444 MUXES_12 ( .A(A[12]), .B(B[12]), .S(n2), .Y(Y[12]) );
  MUX21_443 MUXES_13 ( .A(A[13]), .B(B[13]), .S(n2), .Y(Y[13]) );
  MUX21_442 MUXES_14 ( .A(A[14]), .B(B[14]), .S(n2), .Y(Y[14]) );
  MUX21_441 MUXES_15 ( .A(A[15]), .B(B[15]), .S(n2), .Y(Y[15]) );
  MUX21_440 MUXES_16 ( .A(A[16]), .B(B[16]), .S(n2), .Y(Y[16]) );
  MUX21_439 MUXES_17 ( .A(A[17]), .B(B[17]), .S(n2), .Y(Y[17]) );
  MUX21_438 MUXES_18 ( .A(A[18]), .B(B[18]), .S(n2), .Y(Y[18]) );
  MUX21_437 MUXES_19 ( .A(A[19]), .B(B[19]), .S(n2), .Y(Y[19]) );
  MUX21_436 MUXES_20 ( .A(A[20]), .B(B[20]), .S(n2), .Y(Y[20]) );
  MUX21_435 MUXES_21 ( .A(A[21]), .B(B[21]), .S(n2), .Y(Y[21]) );
  MUX21_434 MUXES_22 ( .A(A[22]), .B(B[22]), .S(n2), .Y(Y[22]) );
  MUX21_433 MUXES_23 ( .A(A[23]), .B(B[23]), .S(n2), .Y(Y[23]) );
  MUX21_432 MUXES_24 ( .A(A[24]), .B(B[24]), .S(n3), .Y(Y[24]) );
  MUX21_431 MUXES_25 ( .A(A[25]), .B(B[25]), .S(n3), .Y(Y[25]) );
  MUX21_430 MUXES_26 ( .A(A[26]), .B(B[26]), .S(n3), .Y(Y[26]) );
  MUX21_429 MUXES_27 ( .A(A[27]), .B(B[27]), .S(n3), .Y(Y[27]) );
  MUX21_428 MUXES_28 ( .A(A[28]), .B(B[28]), .S(n3), .Y(Y[28]) );
  MUX21_427 MUXES_29 ( .A(A[29]), .B(B[29]), .S(n3), .Y(Y[29]) );
  MUX21_426 MUXES_30 ( .A(A[30]), .B(B[30]), .S(n3), .Y(Y[30]) );
  MUX21_425 MUXES_31 ( .A(A[31]), .B(B[31]), .S(n3), .Y(Y[31]) );
  BUF_X1 U1 ( .A(SEL), .Z(n1) );
  BUF_X1 U2 ( .A(SEL), .Z(n2) );
  BUF_X1 U3 ( .A(SEL), .Z(n3) );
endmodule


module WB ( mem_out, alu_out, S3, \output  );
  input [31:0] mem_out;
  input [31:0] alu_out;
  output [31:0] \output ;
  input S3;


  MUX21_GENERIC_NBIT32_2 MUX ( .A(mem_out), .B(alu_out), .SEL(S3), .Y(\output ) );
endmodule


module DataPath_MEM_SIZE128_WORD_size32_NREG32 ( CLK, RST, RF1, RF2, EN1, S1, 
        S2, ALU3, ALU2, ALU1, ALU0, SN, LnS, BHU1, BHU0, Wrd, EN3, S3, WF1, Ld, 
        instr, IRAM_addr, DRAM_data_out, MMU_out, DRAM_addr, DRAM_data_in, 
        opcode, func, OVF );
  input [31:0] instr;
  output [31:0] IRAM_addr;
  input [31:0] DRAM_data_out;
  output [1:0] MMU_out;
  output [8:0] DRAM_addr;
  output [31:0] DRAM_data_in;
  output [5:0] opcode;
  output [10:0] func;
  input CLK, RST, RF1, RF2, EN1, S1, S2, ALU3, ALU2, ALU1, ALU0, SN, LnS, BHU1,
         BHU0, Wrd, EN3, S3, WF1, Ld;
  output OVF;
  wire   flag_signal, hazard_NPC_sel, s_flag_structHzd, s_flag_ismul, n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12;
  wire   [31:0] PC_reg;
  wire   [31:0] NPC_reg;
  wire   [31:0] IR_reg;
  wire   [31:0] Imm_reg;
  wire   [31:0] RA_reg;
  wire   [31:0] RB_reg;
  wire   [4:0] RSA_reg;
  wire   [4:0] RSB_reg;
  wire   [4:0] RD_regexe;
  wire   [31:0] ALU_reg;
  wire   [31:0] ME_reg;
  wire   [4:0] RD_regmem;
  wire   [31:0] LMD_reg;
  wire   [31:0] ALU_regmem;
  wire   [4:0] RD_regwb;
  wire   [31:0] PC_muxout;
  wire   [31:0] NPC_fetchout;
  wire   [31:0] NOP_MUX_OUT;
  wire   [31:0] IMM_decout;
  wire   [31:0] RA_decout;
  wire   [31:0] RB_decout;
  wire   [4:0] RD_decout;
  wire   [4:0] RSA_decout;
  wire   [4:0] RSB_decout;
  wire   [31:0] ALU_exeout;
  wire   [31:0] ME_exeout;
  wire   [4:0] RD_exeout;
  wire   [31:0] mem_out;
  wire   [31:0] ALU_memout;
  wire   [4:0] RD_memout;
  wire   [31:0] s_NPC_jump;
  wire   [31:0] hazard_NPC;
  wire   [31:0] WB_data;
  wire   [4:0] s_RD_inmul;

  DFFR_X1 \ALU_regmem_reg[0]  ( .D(ALU_memout[0]), .CK(CLK), .RN(n8), .Q(
        ALU_regmem[0]) );
  DFFR_X1 \IR_reg_reg[0]  ( .D(NOP_MUX_OUT[0]), .CK(CLK), .RN(n4), .Q(
        IR_reg[0]) );
  DFFR_X1 \IR_reg_reg[1]  ( .D(NOP_MUX_OUT[1]), .CK(CLK), .RN(n8), .Q(
        IR_reg[1]) );
  DFFR_X1 \IR_reg_reg[2]  ( .D(NOP_MUX_OUT[2]), .CK(CLK), .RN(n8), .Q(
        IR_reg[2]) );
  DFFR_X1 \IR_reg_reg[3]  ( .D(NOP_MUX_OUT[3]), .CK(CLK), .RN(n8), .Q(
        IR_reg[3]) );
  DFFR_X1 \IR_reg_reg[4]  ( .D(NOP_MUX_OUT[4]), .CK(CLK), .RN(n8), .Q(
        IR_reg[4]) );
  DFFR_X1 \IR_reg_reg[5]  ( .D(NOP_MUX_OUT[5]), .CK(CLK), .RN(n8), .Q(
        IR_reg[5]) );
  DFFR_X1 \IR_reg_reg[6]  ( .D(NOP_MUX_OUT[6]), .CK(CLK), .RN(n8), .Q(
        IR_reg[6]) );
  DFFR_X1 \IR_reg_reg[7]  ( .D(NOP_MUX_OUT[7]), .CK(CLK), .RN(n8), .Q(
        IR_reg[7]) );
  DFFR_X1 \IR_reg_reg[8]  ( .D(NOP_MUX_OUT[8]), .CK(CLK), .RN(n8), .Q(
        IR_reg[8]) );
  DFFR_X1 \IR_reg_reg[9]  ( .D(NOP_MUX_OUT[9]), .CK(CLK), .RN(n8), .Q(
        IR_reg[9]) );
  DFFR_X1 \IR_reg_reg[10]  ( .D(NOP_MUX_OUT[10]), .CK(CLK), .RN(n8), .Q(
        IR_reg[10]) );
  DFFR_X1 \IR_reg_reg[11]  ( .D(NOP_MUX_OUT[11]), .CK(CLK), .RN(n8), .Q(
        IR_reg[11]) );
  DFFR_X1 \IR_reg_reg[12]  ( .D(NOP_MUX_OUT[12]), .CK(CLK), .RN(n8), .Q(
        IR_reg[12]) );
  DFFR_X1 \IR_reg_reg[13]  ( .D(NOP_MUX_OUT[13]), .CK(CLK), .RN(n7), .Q(
        IR_reg[13]) );
  DFFR_X1 \IR_reg_reg[14]  ( .D(NOP_MUX_OUT[14]), .CK(CLK), .RN(n7), .Q(
        IR_reg[14]) );
  DFFR_X1 \IR_reg_reg[15]  ( .D(NOP_MUX_OUT[15]), .CK(CLK), .RN(n7), .Q(
        IR_reg[15]) );
  DFFR_X1 \IR_reg_reg[16]  ( .D(NOP_MUX_OUT[16]), .CK(CLK), .RN(n7), .Q(
        IR_reg[16]) );
  DFFR_X1 \IR_reg_reg[17]  ( .D(NOP_MUX_OUT[17]), .CK(CLK), .RN(n7), .Q(
        IR_reg[17]) );
  DFFR_X1 \IR_reg_reg[18]  ( .D(NOP_MUX_OUT[18]), .CK(CLK), .RN(n7), .Q(
        IR_reg[18]) );
  DFFR_X1 \IR_reg_reg[19]  ( .D(NOP_MUX_OUT[19]), .CK(CLK), .RN(n7), .Q(
        IR_reg[19]) );
  DFFR_X1 \IR_reg_reg[20]  ( .D(NOP_MUX_OUT[20]), .CK(CLK), .RN(n7), .Q(
        IR_reg[20]) );
  DFFR_X1 \IR_reg_reg[21]  ( .D(NOP_MUX_OUT[21]), .CK(CLK), .RN(n7), .Q(
        IR_reg[21]) );
  DFFR_X1 \IR_reg_reg[22]  ( .D(NOP_MUX_OUT[22]), .CK(CLK), .RN(n7), .Q(
        IR_reg[22]) );
  DFFR_X1 \IR_reg_reg[23]  ( .D(NOP_MUX_OUT[23]), .CK(CLK), .RN(n7), .Q(
        IR_reg[23]) );
  DFFR_X1 \IR_reg_reg[24]  ( .D(NOP_MUX_OUT[24]), .CK(CLK), .RN(n7), .Q(
        IR_reg[24]) );
  DFFR_X1 \IR_reg_reg[25]  ( .D(NOP_MUX_OUT[25]), .CK(CLK), .RN(n7), .Q(
        IR_reg[25]) );
  DFFS_X1 \IR_reg_reg[26]  ( .D(NOP_MUX_OUT[26]), .CK(CLK), .SN(n12), .Q(
        IR_reg[26]) );
  DFFR_X1 \IR_reg_reg[27]  ( .D(NOP_MUX_OUT[27]), .CK(CLK), .RN(n7), .Q(
        IR_reg[27]) );
  DFFR_X1 \IR_reg_reg[29]  ( .D(NOP_MUX_OUT[29]), .CK(CLK), .RN(n7), .Q(
        IR_reg[29]) );
  DFFR_X1 \IR_reg_reg[31]  ( .D(NOP_MUX_OUT[31]), .CK(CLK), .RN(n7), .Q(
        IR_reg[31]) );
  DFFR_X1 \NPC_reg_reg[0]  ( .D(NPC_fetchout[0]), .CK(CLK), .RN(n7), .Q(
        NPC_reg[0]) );
  DFFR_X1 \NPC_reg_reg[1]  ( .D(NPC_fetchout[1]), .CK(CLK), .RN(n7), .Q(
        NPC_reg[1]) );
  DFFR_X1 \NPC_reg_reg[2]  ( .D(NPC_fetchout[2]), .CK(CLK), .RN(n7), .Q(
        NPC_reg[2]) );
  DFFR_X1 \NPC_reg_reg[3]  ( .D(NPC_fetchout[3]), .CK(CLK), .RN(n7), .Q(
        NPC_reg[3]) );
  DFFR_X1 \NPC_reg_reg[4]  ( .D(NPC_fetchout[4]), .CK(CLK), .RN(n7), .Q(
        NPC_reg[4]) );
  DFFR_X1 \NPC_reg_reg[5]  ( .D(NPC_fetchout[5]), .CK(CLK), .RN(n7), .Q(
        NPC_reg[5]) );
  DFFR_X1 \NPC_reg_reg[6]  ( .D(NPC_fetchout[6]), .CK(CLK), .RN(n7), .Q(
        NPC_reg[6]) );
  DFFR_X1 \NPC_reg_reg[7]  ( .D(NPC_fetchout[7]), .CK(CLK), .RN(n7), .Q(
        NPC_reg[7]) );
  DFFR_X1 \NPC_reg_reg[8]  ( .D(NPC_fetchout[8]), .CK(CLK), .RN(n7), .Q(
        NPC_reg[8]) );
  DFFR_X1 \NPC_reg_reg[9]  ( .D(NPC_fetchout[9]), .CK(CLK), .RN(n7), .Q(
        NPC_reg[9]) );
  DFFR_X1 \NPC_reg_reg[10]  ( .D(NPC_fetchout[10]), .CK(CLK), .RN(n7), .Q(
        NPC_reg[10]) );
  DFFR_X1 \NPC_reg_reg[11]  ( .D(NPC_fetchout[11]), .CK(CLK), .RN(n7), .Q(
        NPC_reg[11]) );
  DFFR_X1 \NPC_reg_reg[12]  ( .D(NPC_fetchout[12]), .CK(CLK), .RN(n7), .Q(
        NPC_reg[12]) );
  DFFR_X1 \NPC_reg_reg[13]  ( .D(NPC_fetchout[13]), .CK(CLK), .RN(n7), .Q(
        NPC_reg[13]) );
  DFFR_X1 \NPC_reg_reg[14]  ( .D(NPC_fetchout[14]), .CK(CLK), .RN(n7), .Q(
        NPC_reg[14]) );
  DFFR_X1 \NPC_reg_reg[15]  ( .D(NPC_fetchout[15]), .CK(CLK), .RN(n7), .Q(
        NPC_reg[15]) );
  DFFR_X1 \NPC_reg_reg[16]  ( .D(NPC_fetchout[16]), .CK(CLK), .RN(n7), .Q(
        NPC_reg[16]) );
  DFFR_X1 \NPC_reg_reg[17]  ( .D(NPC_fetchout[17]), .CK(CLK), .RN(n7), .Q(
        NPC_reg[17]) );
  DFFR_X1 \NPC_reg_reg[18]  ( .D(NPC_fetchout[18]), .CK(CLK), .RN(n7), .Q(
        NPC_reg[18]) );
  DFFR_X1 \NPC_reg_reg[19]  ( .D(NPC_fetchout[19]), .CK(CLK), .RN(n7), .Q(
        NPC_reg[19]) );
  DFFR_X1 \NPC_reg_reg[20]  ( .D(NPC_fetchout[20]), .CK(CLK), .RN(n7), .Q(
        NPC_reg[20]) );
  DFFR_X1 \NPC_reg_reg[21]  ( .D(NPC_fetchout[21]), .CK(CLK), .RN(n7), .Q(
        NPC_reg[21]) );
  DFFR_X1 \NPC_reg_reg[22]  ( .D(NPC_fetchout[22]), .CK(CLK), .RN(n7), .Q(
        NPC_reg[22]) );
  DFFR_X1 \NPC_reg_reg[23]  ( .D(NPC_fetchout[23]), .CK(CLK), .RN(n7), .Q(
        NPC_reg[23]) );
  DFFR_X1 \NPC_reg_reg[24]  ( .D(NPC_fetchout[24]), .CK(CLK), .RN(n7), .Q(
        NPC_reg[24]) );
  DFFR_X1 \NPC_reg_reg[25]  ( .D(NPC_fetchout[25]), .CK(CLK), .RN(n7), .Q(
        NPC_reg[25]) );
  DFFR_X1 \NPC_reg_reg[26]  ( .D(NPC_fetchout[26]), .CK(CLK), .RN(n6), .Q(
        NPC_reg[26]) );
  DFFR_X1 \NPC_reg_reg[27]  ( .D(NPC_fetchout[27]), .CK(CLK), .RN(n6), .Q(
        NPC_reg[27]) );
  DFFR_X1 \NPC_reg_reg[28]  ( .D(NPC_fetchout[28]), .CK(CLK), .RN(n6), .Q(
        NPC_reg[28]) );
  DFFR_X1 \NPC_reg_reg[29]  ( .D(NPC_fetchout[29]), .CK(CLK), .RN(n6), .Q(
        NPC_reg[29]) );
  DFFR_X1 \NPC_reg_reg[30]  ( .D(NPC_fetchout[30]), .CK(CLK), .RN(n6), .Q(
        NPC_reg[30]) );
  DFFR_X1 \NPC_reg_reg[31]  ( .D(NPC_fetchout[31]), .CK(CLK), .RN(n6), .Q(
        NPC_reg[31]) );
  DFFR_X1 \PC_reg_reg[0]  ( .D(PC_muxout[0]), .CK(CLK), .RN(n6), .Q(PC_reg[0])
         );
  DFFR_X1 \PC_reg_reg[1]  ( .D(PC_muxout[1]), .CK(CLK), .RN(n6), .Q(PC_reg[1])
         );
  DFFR_X1 \PC_reg_reg[2]  ( .D(PC_muxout[2]), .CK(CLK), .RN(n6), .Q(PC_reg[2])
         );
  DFFR_X1 \PC_reg_reg[3]  ( .D(PC_muxout[3]), .CK(CLK), .RN(n6), .Q(PC_reg[3])
         );
  DFFR_X1 \PC_reg_reg[4]  ( .D(PC_muxout[4]), .CK(CLK), .RN(n6), .Q(PC_reg[4])
         );
  DFFR_X1 \PC_reg_reg[5]  ( .D(PC_muxout[5]), .CK(CLK), .RN(n6), .Q(PC_reg[5])
         );
  DFFR_X1 \PC_reg_reg[6]  ( .D(PC_muxout[6]), .CK(CLK), .RN(n6), .Q(PC_reg[6])
         );
  DFFR_X1 \PC_reg_reg[7]  ( .D(PC_muxout[7]), .CK(CLK), .RN(n6), .Q(PC_reg[7])
         );
  DFFR_X1 \PC_reg_reg[8]  ( .D(PC_muxout[8]), .CK(CLK), .RN(n6), .Q(PC_reg[8])
         );
  DFFR_X1 \PC_reg_reg[9]  ( .D(PC_muxout[9]), .CK(CLK), .RN(n6), .Q(PC_reg[9])
         );
  DFFR_X1 \PC_reg_reg[10]  ( .D(PC_muxout[10]), .CK(CLK), .RN(n6), .Q(
        PC_reg[10]) );
  DFFR_X1 \PC_reg_reg[11]  ( .D(PC_muxout[11]), .CK(CLK), .RN(n6), .Q(
        PC_reg[11]) );
  DFFR_X1 \PC_reg_reg[12]  ( .D(PC_muxout[12]), .CK(CLK), .RN(n6), .Q(
        PC_reg[12]) );
  DFFR_X1 \PC_reg_reg[13]  ( .D(PC_muxout[13]), .CK(CLK), .RN(n6), .Q(
        PC_reg[13]) );
  DFFR_X1 \PC_reg_reg[14]  ( .D(PC_muxout[14]), .CK(CLK), .RN(n6), .Q(
        PC_reg[14]) );
  DFFR_X1 \PC_reg_reg[15]  ( .D(PC_muxout[15]), .CK(CLK), .RN(n6), .Q(
        PC_reg[15]) );
  DFFR_X1 \PC_reg_reg[16]  ( .D(PC_muxout[16]), .CK(CLK), .RN(n6), .Q(
        PC_reg[16]) );
  DFFR_X1 \PC_reg_reg[17]  ( .D(PC_muxout[17]), .CK(CLK), .RN(n6), .Q(
        PC_reg[17]) );
  DFFR_X1 \PC_reg_reg[18]  ( .D(PC_muxout[18]), .CK(CLK), .RN(n6), .Q(
        PC_reg[18]) );
  DFFR_X1 \PC_reg_reg[19]  ( .D(PC_muxout[19]), .CK(CLK), .RN(n6), .Q(
        PC_reg[19]) );
  DFFR_X1 \PC_reg_reg[20]  ( .D(PC_muxout[20]), .CK(CLK), .RN(n6), .Q(
        PC_reg[20]) );
  DFFR_X1 \PC_reg_reg[21]  ( .D(PC_muxout[21]), .CK(CLK), .RN(n6), .Q(
        PC_reg[21]) );
  DFFR_X1 \PC_reg_reg[22]  ( .D(PC_muxout[22]), .CK(CLK), .RN(n6), .Q(
        PC_reg[22]) );
  DFFR_X1 \PC_reg_reg[23]  ( .D(PC_muxout[23]), .CK(CLK), .RN(n6), .Q(
        PC_reg[23]) );
  DFFR_X1 \PC_reg_reg[24]  ( .D(PC_muxout[24]), .CK(CLK), .RN(n6), .Q(
        PC_reg[24]) );
  DFFR_X1 \PC_reg_reg[25]  ( .D(PC_muxout[25]), .CK(CLK), .RN(n6), .Q(
        PC_reg[25]) );
  DFFR_X1 \PC_reg_reg[26]  ( .D(PC_muxout[26]), .CK(CLK), .RN(n6), .Q(
        PC_reg[26]) );
  DFFR_X1 \PC_reg_reg[27]  ( .D(PC_muxout[27]), .CK(CLK), .RN(n6), .Q(
        PC_reg[27]) );
  DFFR_X1 \PC_reg_reg[28]  ( .D(PC_muxout[28]), .CK(CLK), .RN(n6), .Q(
        PC_reg[28]) );
  DFFR_X1 \PC_reg_reg[29]  ( .D(PC_muxout[29]), .CK(CLK), .RN(n6), .Q(
        PC_reg[29]) );
  DFFR_X1 \PC_reg_reg[30]  ( .D(PC_muxout[30]), .CK(CLK), .RN(n6), .Q(
        PC_reg[30]) );
  DFFR_X1 \PC_reg_reg[31]  ( .D(PC_muxout[31]), .CK(CLK), .RN(n6), .Q(
        PC_reg[31]) );
  DFFR_X1 \RD_regexe_reg[0]  ( .D(RD_decout[0]), .CK(CLK), .RN(n6), .Q(
        RD_regexe[0]) );
  DFFR_X1 \RD_regexe_reg[1]  ( .D(RD_decout[1]), .CK(CLK), .RN(n6), .Q(
        RD_regexe[1]) );
  DFFR_X1 \RD_regexe_reg[2]  ( .D(RD_decout[2]), .CK(CLK), .RN(n6), .Q(
        RD_regexe[2]) );
  DFFR_X1 \RD_regexe_reg[3]  ( .D(RD_decout[3]), .CK(CLK), .RN(n5), .Q(
        RD_regexe[3]) );
  DFFR_X1 \RD_regexe_reg[4]  ( .D(RD_decout[4]), .CK(CLK), .RN(n5), .Q(
        RD_regexe[4]) );
  DFFR_X1 \RSB_reg_reg[0]  ( .D(RSB_decout[0]), .CK(CLK), .RN(n5), .Q(
        RSB_reg[0]) );
  DFFR_X1 \RSB_reg_reg[1]  ( .D(RSB_decout[1]), .CK(CLK), .RN(n5), .Q(
        RSB_reg[1]) );
  DFFR_X1 \RSB_reg_reg[2]  ( .D(RSB_decout[2]), .CK(CLK), .RN(n5), .Q(
        RSB_reg[2]) );
  DFFR_X1 \RSB_reg_reg[3]  ( .D(RSB_decout[3]), .CK(CLK), .RN(n5), .Q(
        RSB_reg[3]) );
  DFFR_X1 \RSB_reg_reg[4]  ( .D(RSB_decout[4]), .CK(CLK), .RN(n5), .Q(
        RSB_reg[4]) );
  DFFR_X1 \RSA_reg_reg[0]  ( .D(RSA_decout[0]), .CK(CLK), .RN(n5), .Q(
        RSA_reg[0]) );
  DFFR_X1 \RSA_reg_reg[1]  ( .D(RSA_decout[1]), .CK(CLK), .RN(n5), .Q(
        RSA_reg[1]) );
  DFFR_X1 \RSA_reg_reg[2]  ( .D(RSA_decout[2]), .CK(CLK), .RN(n5), .Q(
        RSA_reg[2]) );
  DFFR_X1 \RSA_reg_reg[3]  ( .D(RSA_decout[3]), .CK(CLK), .RN(n5), .Q(
        RSA_reg[3]) );
  DFFR_X1 \RSA_reg_reg[4]  ( .D(RSA_decout[4]), .CK(CLK), .RN(n5), .Q(
        RSA_reg[4]) );
  DFFR_X1 \RB_reg_reg[0]  ( .D(RB_decout[0]), .CK(CLK), .RN(n5), .Q(RB_reg[0])
         );
  DFFR_X1 \RB_reg_reg[1]  ( .D(RB_decout[1]), .CK(CLK), .RN(n5), .Q(RB_reg[1])
         );
  DFFR_X1 \RB_reg_reg[2]  ( .D(RB_decout[2]), .CK(CLK), .RN(n5), .Q(RB_reg[2])
         );
  DFFR_X1 \RB_reg_reg[3]  ( .D(RB_decout[3]), .CK(CLK), .RN(n5), .Q(RB_reg[3])
         );
  DFFR_X1 \RB_reg_reg[4]  ( .D(RB_decout[4]), .CK(CLK), .RN(n5), .Q(RB_reg[4])
         );
  DFFR_X1 \RB_reg_reg[5]  ( .D(RB_decout[5]), .CK(CLK), .RN(n5), .Q(RB_reg[5])
         );
  DFFR_X1 \RB_reg_reg[6]  ( .D(RB_decout[6]), .CK(CLK), .RN(n5), .Q(RB_reg[6])
         );
  DFFR_X1 \RB_reg_reg[7]  ( .D(RB_decout[7]), .CK(CLK), .RN(n5), .Q(RB_reg[7])
         );
  DFFR_X1 \RB_reg_reg[8]  ( .D(RB_decout[8]), .CK(CLK), .RN(n5), .Q(RB_reg[8])
         );
  DFFR_X1 \RB_reg_reg[9]  ( .D(RB_decout[9]), .CK(CLK), .RN(n5), .Q(RB_reg[9])
         );
  DFFR_X1 \RB_reg_reg[10]  ( .D(RB_decout[10]), .CK(CLK), .RN(n5), .Q(
        RB_reg[10]) );
  DFFR_X1 \RB_reg_reg[11]  ( .D(RB_decout[11]), .CK(CLK), .RN(n5), .Q(
        RB_reg[11]) );
  DFFR_X1 \RB_reg_reg[12]  ( .D(RB_decout[12]), .CK(CLK), .RN(n5), .Q(
        RB_reg[12]) );
  DFFR_X1 \RB_reg_reg[13]  ( .D(RB_decout[13]), .CK(CLK), .RN(n5), .Q(
        RB_reg[13]) );
  DFFR_X1 \RB_reg_reg[14]  ( .D(RB_decout[14]), .CK(CLK), .RN(n5), .Q(
        RB_reg[14]) );
  DFFR_X1 \RB_reg_reg[15]  ( .D(RB_decout[15]), .CK(CLK), .RN(n5), .Q(
        RB_reg[15]) );
  DFFR_X1 \RB_reg_reg[16]  ( .D(RB_decout[16]), .CK(CLK), .RN(n5), .Q(
        RB_reg[16]) );
  DFFR_X1 \RB_reg_reg[17]  ( .D(RB_decout[17]), .CK(CLK), .RN(n5), .Q(
        RB_reg[17]) );
  DFFR_X1 \RB_reg_reg[18]  ( .D(RB_decout[18]), .CK(CLK), .RN(n5), .Q(
        RB_reg[18]) );
  DFFR_X1 \RB_reg_reg[19]  ( .D(RB_decout[19]), .CK(CLK), .RN(n5), .Q(
        RB_reg[19]) );
  DFFR_X1 \RB_reg_reg[20]  ( .D(RB_decout[20]), .CK(CLK), .RN(n5), .Q(
        RB_reg[20]) );
  DFFR_X1 \RB_reg_reg[21]  ( .D(RB_decout[21]), .CK(CLK), .RN(n5), .Q(
        RB_reg[21]) );
  DFFR_X1 \RB_reg_reg[22]  ( .D(RB_decout[22]), .CK(CLK), .RN(n5), .Q(
        RB_reg[22]) );
  DFFR_X1 \RB_reg_reg[23]  ( .D(RB_decout[23]), .CK(CLK), .RN(n5), .Q(
        RB_reg[23]) );
  DFFR_X1 \RB_reg_reg[24]  ( .D(RB_decout[24]), .CK(CLK), .RN(n5), .Q(
        RB_reg[24]) );
  DFFR_X1 \RB_reg_reg[25]  ( .D(RB_decout[25]), .CK(CLK), .RN(n5), .Q(
        RB_reg[25]) );
  DFFR_X1 \RB_reg_reg[26]  ( .D(RB_decout[26]), .CK(CLK), .RN(n5), .Q(
        RB_reg[26]) );
  DFFR_X1 \RB_reg_reg[27]  ( .D(RB_decout[27]), .CK(CLK), .RN(n5), .Q(
        RB_reg[27]) );
  DFFR_X1 \RB_reg_reg[28]  ( .D(RB_decout[28]), .CK(CLK), .RN(n5), .Q(
        RB_reg[28]) );
  DFFR_X1 \RB_reg_reg[29]  ( .D(RB_decout[29]), .CK(CLK), .RN(n5), .Q(
        RB_reg[29]) );
  DFFR_X1 \RB_reg_reg[30]  ( .D(RB_decout[30]), .CK(CLK), .RN(n4), .Q(
        RB_reg[30]) );
  DFFR_X1 \RB_reg_reg[31]  ( .D(RB_decout[31]), .CK(CLK), .RN(n4), .Q(
        RB_reg[31]) );
  DFFR_X1 \RA_reg_reg[0]  ( .D(RA_decout[0]), .CK(CLK), .RN(n4), .Q(RA_reg[0])
         );
  DFFR_X1 \RA_reg_reg[1]  ( .D(RA_decout[1]), .CK(CLK), .RN(n4), .Q(RA_reg[1])
         );
  DFFR_X1 \RA_reg_reg[2]  ( .D(RA_decout[2]), .CK(CLK), .RN(n4), .Q(RA_reg[2])
         );
  DFFR_X1 \RA_reg_reg[3]  ( .D(RA_decout[3]), .CK(CLK), .RN(n4), .Q(RA_reg[3])
         );
  DFFR_X1 \RA_reg_reg[4]  ( .D(RA_decout[4]), .CK(CLK), .RN(n4), .Q(RA_reg[4])
         );
  DFFR_X1 \RA_reg_reg[5]  ( .D(RA_decout[5]), .CK(CLK), .RN(n4), .Q(RA_reg[5])
         );
  DFFR_X1 \RA_reg_reg[6]  ( .D(RA_decout[6]), .CK(CLK), .RN(n4), .Q(RA_reg[6])
         );
  DFFR_X1 \RA_reg_reg[7]  ( .D(RA_decout[7]), .CK(CLK), .RN(n4), .Q(RA_reg[7])
         );
  DFFR_X1 \RA_reg_reg[8]  ( .D(RA_decout[8]), .CK(CLK), .RN(n4), .Q(RA_reg[8])
         );
  DFFR_X1 \RA_reg_reg[9]  ( .D(RA_decout[9]), .CK(CLK), .RN(n4), .Q(RA_reg[9])
         );
  DFFR_X1 \RA_reg_reg[10]  ( .D(RA_decout[10]), .CK(CLK), .RN(n4), .Q(
        RA_reg[10]) );
  DFFR_X1 \RA_reg_reg[11]  ( .D(RA_decout[11]), .CK(CLK), .RN(n4), .Q(
        RA_reg[11]) );
  DFFR_X1 \RA_reg_reg[12]  ( .D(RA_decout[12]), .CK(CLK), .RN(n4), .Q(
        RA_reg[12]) );
  DFFR_X1 \RA_reg_reg[13]  ( .D(RA_decout[13]), .CK(CLK), .RN(n4), .Q(
        RA_reg[13]) );
  DFFR_X1 \RA_reg_reg[14]  ( .D(RA_decout[14]), .CK(CLK), .RN(n4), .Q(
        RA_reg[14]) );
  DFFR_X1 \RA_reg_reg[15]  ( .D(RA_decout[15]), .CK(CLK), .RN(n4), .Q(
        RA_reg[15]) );
  DFFR_X1 \RA_reg_reg[16]  ( .D(RA_decout[16]), .CK(CLK), .RN(n4), .Q(
        RA_reg[16]) );
  DFFR_X1 \RA_reg_reg[17]  ( .D(RA_decout[17]), .CK(CLK), .RN(n4), .Q(
        RA_reg[17]) );
  DFFR_X1 \RA_reg_reg[18]  ( .D(RA_decout[18]), .CK(CLK), .RN(n4), .Q(
        RA_reg[18]) );
  DFFR_X1 \RA_reg_reg[19]  ( .D(RA_decout[19]), .CK(CLK), .RN(n4), .Q(
        RA_reg[19]) );
  DFFR_X1 \RA_reg_reg[20]  ( .D(RA_decout[20]), .CK(CLK), .RN(n4), .Q(
        RA_reg[20]) );
  DFFR_X1 \RA_reg_reg[21]  ( .D(RA_decout[21]), .CK(CLK), .RN(n4), .Q(
        RA_reg[21]) );
  DFFR_X1 \RA_reg_reg[22]  ( .D(RA_decout[22]), .CK(CLK), .RN(n4), .Q(
        RA_reg[22]) );
  DFFR_X1 \RA_reg_reg[23]  ( .D(RA_decout[23]), .CK(CLK), .RN(n4), .Q(
        RA_reg[23]) );
  DFFR_X1 \RA_reg_reg[24]  ( .D(RA_decout[24]), .CK(CLK), .RN(n4), .Q(
        RA_reg[24]) );
  DFFR_X1 \RA_reg_reg[25]  ( .D(RA_decout[25]), .CK(CLK), .RN(n4), .Q(
        RA_reg[25]) );
  DFFR_X1 \RA_reg_reg[26]  ( .D(RA_decout[26]), .CK(CLK), .RN(n4), .Q(
        RA_reg[26]) );
  DFFR_X1 \RA_reg_reg[27]  ( .D(RA_decout[27]), .CK(CLK), .RN(n4), .Q(
        RA_reg[27]) );
  DFFR_X1 \RA_reg_reg[28]  ( .D(RA_decout[28]), .CK(CLK), .RN(n4), .Q(
        RA_reg[28]) );
  DFFR_X1 \RA_reg_reg[29]  ( .D(RA_decout[29]), .CK(CLK), .RN(n4), .Q(
        RA_reg[29]) );
  DFFR_X1 \RA_reg_reg[30]  ( .D(RA_decout[30]), .CK(CLK), .RN(n6), .Q(
        RA_reg[30]) );
  DFFR_X1 \RA_reg_reg[31]  ( .D(RA_decout[31]), .CK(CLK), .RN(n12), .Q(
        RA_reg[31]) );
  DFFR_X1 \Imm_reg_reg[0]  ( .D(IMM_decout[0]), .CK(CLK), .RN(n12), .Q(
        Imm_reg[0]) );
  DFFR_X1 \Imm_reg_reg[1]  ( .D(IMM_decout[1]), .CK(CLK), .RN(n12), .Q(
        Imm_reg[1]) );
  DFFR_X1 \Imm_reg_reg[2]  ( .D(IMM_decout[2]), .CK(CLK), .RN(n12), .Q(
        Imm_reg[2]) );
  DFFR_X1 \Imm_reg_reg[3]  ( .D(IMM_decout[3]), .CK(CLK), .RN(n12), .Q(
        Imm_reg[3]) );
  DFFR_X1 \Imm_reg_reg[4]  ( .D(IMM_decout[4]), .CK(CLK), .RN(n12), .Q(
        Imm_reg[4]) );
  DFFR_X1 \Imm_reg_reg[5]  ( .D(IMM_decout[5]), .CK(CLK), .RN(n12), .Q(
        Imm_reg[5]) );
  DFFR_X1 \Imm_reg_reg[6]  ( .D(IMM_decout[6]), .CK(CLK), .RN(n12), .Q(
        Imm_reg[6]) );
  DFFR_X1 \Imm_reg_reg[7]  ( .D(IMM_decout[7]), .CK(CLK), .RN(n12), .Q(
        Imm_reg[7]) );
  DFFR_X1 \Imm_reg_reg[8]  ( .D(IMM_decout[8]), .CK(CLK), .RN(n12), .Q(
        Imm_reg[8]) );
  DFFR_X1 \Imm_reg_reg[9]  ( .D(IMM_decout[9]), .CK(CLK), .RN(n12), .Q(
        Imm_reg[9]) );
  DFFR_X1 \Imm_reg_reg[10]  ( .D(IMM_decout[10]), .CK(CLK), .RN(n12), .Q(
        Imm_reg[10]) );
  DFFR_X1 \Imm_reg_reg[11]  ( .D(IMM_decout[11]), .CK(CLK), .RN(n11), .Q(
        Imm_reg[11]) );
  DFFR_X1 \Imm_reg_reg[12]  ( .D(IMM_decout[12]), .CK(CLK), .RN(n12), .Q(
        Imm_reg[12]) );
  DFFR_X1 \Imm_reg_reg[13]  ( .D(IMM_decout[13]), .CK(CLK), .RN(n12), .Q(
        Imm_reg[13]) );
  DFFR_X1 \Imm_reg_reg[14]  ( .D(IMM_decout[14]), .CK(CLK), .RN(n11), .Q(
        Imm_reg[14]) );
  DFFR_X1 \Imm_reg_reg[15]  ( .D(IMM_decout[15]), .CK(CLK), .RN(n12), .Q(
        Imm_reg[15]) );
  DFFR_X1 \Imm_reg_reg[16]  ( .D(IMM_decout[16]), .CK(CLK), .RN(n11), .Q(
        Imm_reg[16]) );
  DFFR_X1 \Imm_reg_reg[17]  ( .D(IMM_decout[17]), .CK(CLK), .RN(n11), .Q(
        Imm_reg[17]) );
  DFFR_X1 \Imm_reg_reg[18]  ( .D(IMM_decout[18]), .CK(CLK), .RN(n11), .Q(
        Imm_reg[18]) );
  DFFR_X1 \Imm_reg_reg[19]  ( .D(IMM_decout[19]), .CK(CLK), .RN(n11), .Q(
        Imm_reg[19]) );
  DFFR_X1 \Imm_reg_reg[20]  ( .D(IMM_decout[20]), .CK(CLK), .RN(n11), .Q(
        Imm_reg[20]) );
  DFFR_X1 \Imm_reg_reg[21]  ( .D(IMM_decout[21]), .CK(CLK), .RN(n11), .Q(
        Imm_reg[21]) );
  DFFR_X1 \Imm_reg_reg[22]  ( .D(IMM_decout[22]), .CK(CLK), .RN(n11), .Q(
        Imm_reg[22]) );
  DFFR_X1 \Imm_reg_reg[23]  ( .D(IMM_decout[23]), .CK(CLK), .RN(n11), .Q(
        Imm_reg[23]) );
  DFFR_X1 \Imm_reg_reg[24]  ( .D(IMM_decout[24]), .CK(CLK), .RN(n11), .Q(
        Imm_reg[24]) );
  DFFR_X1 \Imm_reg_reg[25]  ( .D(IMM_decout[25]), .CK(CLK), .RN(n11), .Q(
        Imm_reg[25]) );
  DFFR_X1 \Imm_reg_reg[26]  ( .D(IMM_decout[26]), .CK(CLK), .RN(n11), .Q(
        Imm_reg[26]) );
  DFFR_X1 \Imm_reg_reg[27]  ( .D(IMM_decout[27]), .CK(CLK), .RN(n11), .Q(
        Imm_reg[27]) );
  DFFR_X1 \Imm_reg_reg[28]  ( .D(IMM_decout[28]), .CK(CLK), .RN(n11), .Q(
        Imm_reg[28]) );
  DFFR_X1 \Imm_reg_reg[29]  ( .D(IMM_decout[29]), .CK(CLK), .RN(n11), .Q(
        Imm_reg[29]) );
  DFFR_X1 \Imm_reg_reg[30]  ( .D(IMM_decout[30]), .CK(CLK), .RN(n11), .Q(
        Imm_reg[30]) );
  DFFR_X1 \Imm_reg_reg[31]  ( .D(IMM_decout[31]), .CK(CLK), .RN(n11), .Q(
        Imm_reg[31]) );
  DFFR_X1 \RD_regmem_reg[0]  ( .D(RD_exeout[0]), .CK(CLK), .RN(n11), .Q(
        RD_regmem[0]) );
  DFFR_X1 \RD_regmem_reg[1]  ( .D(RD_exeout[1]), .CK(CLK), .RN(n11), .Q(
        RD_regmem[1]) );
  DFFR_X1 \RD_regmem_reg[2]  ( .D(RD_exeout[2]), .CK(CLK), .RN(n11), .Q(
        RD_regmem[2]) );
  DFFR_X1 \RD_regmem_reg[3]  ( .D(RD_exeout[3]), .CK(CLK), .RN(n11), .Q(
        RD_regmem[3]) );
  DFFR_X1 \RD_regmem_reg[4]  ( .D(RD_exeout[4]), .CK(CLK), .RN(n11), .Q(
        RD_regmem[4]) );
  DFFR_X1 \ME_reg_reg[0]  ( .D(ME_exeout[0]), .CK(CLK), .RN(n11), .Q(ME_reg[0]) );
  DFFR_X1 \ME_reg_reg[1]  ( .D(ME_exeout[1]), .CK(CLK), .RN(n11), .Q(ME_reg[1]) );
  DFFR_X1 \ME_reg_reg[2]  ( .D(ME_exeout[2]), .CK(CLK), .RN(n11), .Q(ME_reg[2]) );
  DFFR_X1 \ME_reg_reg[3]  ( .D(ME_exeout[3]), .CK(CLK), .RN(n11), .Q(ME_reg[3]) );
  DFFR_X1 \ME_reg_reg[4]  ( .D(ME_exeout[4]), .CK(CLK), .RN(n11), .Q(ME_reg[4]) );
  DFFR_X1 \ME_reg_reg[5]  ( .D(ME_exeout[5]), .CK(CLK), .RN(n11), .Q(ME_reg[5]) );
  DFFR_X1 \ME_reg_reg[6]  ( .D(ME_exeout[6]), .CK(CLK), .RN(n11), .Q(ME_reg[6]) );
  DFFR_X1 \ME_reg_reg[7]  ( .D(ME_exeout[7]), .CK(CLK), .RN(n11), .Q(ME_reg[7]) );
  DFFR_X1 \ME_reg_reg[8]  ( .D(ME_exeout[8]), .CK(CLK), .RN(n11), .Q(ME_reg[8]) );
  DFFR_X1 \ME_reg_reg[9]  ( .D(ME_exeout[9]), .CK(CLK), .RN(n11), .Q(ME_reg[9]) );
  DFFR_X1 \ME_reg_reg[10]  ( .D(ME_exeout[10]), .CK(CLK), .RN(n11), .Q(
        ME_reg[10]) );
  DFFR_X1 \ME_reg_reg[11]  ( .D(ME_exeout[11]), .CK(CLK), .RN(n11), .Q(
        ME_reg[11]) );
  DFFR_X1 \ME_reg_reg[12]  ( .D(ME_exeout[12]), .CK(CLK), .RN(n11), .Q(
        ME_reg[12]) );
  DFFR_X1 \ME_reg_reg[13]  ( .D(ME_exeout[13]), .CK(CLK), .RN(n11), .Q(
        ME_reg[13]) );
  DFFR_X1 \ME_reg_reg[14]  ( .D(ME_exeout[14]), .CK(CLK), .RN(n11), .Q(
        ME_reg[14]) );
  DFFR_X1 \ME_reg_reg[15]  ( .D(ME_exeout[15]), .CK(CLK), .RN(n11), .Q(
        ME_reg[15]) );
  DFFR_X1 \ME_reg_reg[16]  ( .D(ME_exeout[16]), .CK(CLK), .RN(n11), .Q(
        ME_reg[16]) );
  DFFR_X1 \ME_reg_reg[17]  ( .D(ME_exeout[17]), .CK(CLK), .RN(n11), .Q(
        ME_reg[17]) );
  DFFR_X1 \ME_reg_reg[18]  ( .D(ME_exeout[18]), .CK(CLK), .RN(n11), .Q(
        ME_reg[18]) );
  DFFR_X1 \ME_reg_reg[19]  ( .D(ME_exeout[19]), .CK(CLK), .RN(n10), .Q(
        ME_reg[19]) );
  DFFR_X1 \ME_reg_reg[20]  ( .D(ME_exeout[20]), .CK(CLK), .RN(n10), .Q(
        ME_reg[20]) );
  DFFR_X1 \ME_reg_reg[21]  ( .D(ME_exeout[21]), .CK(CLK), .RN(n10), .Q(
        ME_reg[21]) );
  DFFR_X1 \ME_reg_reg[22]  ( .D(ME_exeout[22]), .CK(CLK), .RN(n10), .Q(
        ME_reg[22]) );
  DFFR_X1 \ME_reg_reg[23]  ( .D(ME_exeout[23]), .CK(CLK), .RN(n10), .Q(
        ME_reg[23]) );
  DFFR_X1 \ME_reg_reg[24]  ( .D(ME_exeout[24]), .CK(CLK), .RN(n10), .Q(
        ME_reg[24]) );
  DFFR_X1 \ME_reg_reg[25]  ( .D(ME_exeout[25]), .CK(CLK), .RN(n10), .Q(
        ME_reg[25]) );
  DFFR_X1 \ME_reg_reg[26]  ( .D(ME_exeout[26]), .CK(CLK), .RN(n10), .Q(
        ME_reg[26]) );
  DFFR_X1 \ME_reg_reg[27]  ( .D(ME_exeout[27]), .CK(CLK), .RN(n10), .Q(
        ME_reg[27]) );
  DFFR_X1 \ME_reg_reg[28]  ( .D(ME_exeout[28]), .CK(CLK), .RN(n10), .Q(
        ME_reg[28]) );
  DFFR_X1 \ME_reg_reg[29]  ( .D(ME_exeout[29]), .CK(CLK), .RN(n10), .Q(
        ME_reg[29]) );
  DFFR_X1 \ME_reg_reg[30]  ( .D(ME_exeout[30]), .CK(CLK), .RN(n10), .Q(
        ME_reg[30]) );
  DFFR_X1 \ME_reg_reg[31]  ( .D(ME_exeout[31]), .CK(CLK), .RN(n10), .Q(
        ME_reg[31]) );
  DFFR_X1 \ALU_reg_reg[0]  ( .D(ALU_exeout[0]), .CK(CLK), .RN(n10), .Q(
        ALU_reg[0]) );
  DFFR_X1 \ALU_reg_reg[1]  ( .D(ALU_exeout[1]), .CK(CLK), .RN(n10), .Q(
        ALU_reg[1]) );
  DFFR_X1 \ALU_reg_reg[2]  ( .D(ALU_exeout[2]), .CK(CLK), .RN(n10), .Q(
        ALU_reg[2]) );
  DFFR_X1 \ALU_reg_reg[3]  ( .D(ALU_exeout[3]), .CK(CLK), .RN(n10), .Q(
        ALU_reg[3]) );
  DFFR_X1 \ALU_reg_reg[4]  ( .D(ALU_exeout[4]), .CK(CLK), .RN(n10), .Q(
        ALU_reg[4]) );
  DFFR_X1 \ALU_reg_reg[5]  ( .D(ALU_exeout[5]), .CK(CLK), .RN(n10), .Q(
        ALU_reg[5]) );
  DFFR_X1 \ALU_reg_reg[6]  ( .D(ALU_exeout[6]), .CK(CLK), .RN(n10), .Q(
        ALU_reg[6]) );
  DFFR_X1 \ALU_reg_reg[7]  ( .D(ALU_exeout[7]), .CK(CLK), .RN(n10), .Q(
        ALU_reg[7]) );
  DFFR_X1 \ALU_reg_reg[8]  ( .D(ALU_exeout[8]), .CK(CLK), .RN(n10), .Q(
        ALU_reg[8]) );
  DFFR_X1 \ALU_reg_reg[9]  ( .D(ALU_exeout[9]), .CK(CLK), .RN(n10), .Q(
        ALU_reg[9]) );
  DFFR_X1 \ALU_reg_reg[10]  ( .D(ALU_exeout[10]), .CK(CLK), .RN(n10), .Q(
        ALU_reg[10]) );
  DFFR_X1 \ALU_reg_reg[11]  ( .D(ALU_exeout[11]), .CK(CLK), .RN(n10), .Q(
        ALU_reg[11]) );
  DFFR_X1 \ALU_reg_reg[12]  ( .D(ALU_exeout[12]), .CK(CLK), .RN(n10), .Q(
        ALU_reg[12]) );
  DFFR_X1 \ALU_reg_reg[13]  ( .D(ALU_exeout[13]), .CK(CLK), .RN(n10), .Q(
        ALU_reg[13]) );
  DFFR_X1 \ALU_reg_reg[14]  ( .D(ALU_exeout[14]), .CK(CLK), .RN(n10), .Q(
        ALU_reg[14]) );
  DFFR_X1 \ALU_reg_reg[15]  ( .D(ALU_exeout[15]), .CK(CLK), .RN(n10), .Q(
        ALU_reg[15]) );
  DFFR_X1 \ALU_reg_reg[16]  ( .D(ALU_exeout[16]), .CK(CLK), .RN(n10), .Q(
        ALU_reg[16]) );
  DFFR_X1 \ALU_reg_reg[17]  ( .D(ALU_exeout[17]), .CK(CLK), .RN(n10), .Q(
        ALU_reg[17]) );
  DFFR_X1 \ALU_reg_reg[18]  ( .D(ALU_exeout[18]), .CK(CLK), .RN(n10), .Q(
        ALU_reg[18]) );
  DFFR_X1 \ALU_reg_reg[19]  ( .D(ALU_exeout[19]), .CK(CLK), .RN(n10), .Q(
        ALU_reg[19]) );
  DFFR_X1 \ALU_reg_reg[20]  ( .D(ALU_exeout[20]), .CK(CLK), .RN(n10), .Q(
        ALU_reg[20]) );
  DFFR_X1 \ALU_reg_reg[21]  ( .D(ALU_exeout[21]), .CK(CLK), .RN(n10), .Q(
        ALU_reg[21]) );
  DFFR_X1 \ALU_reg_reg[22]  ( .D(ALU_exeout[22]), .CK(CLK), .RN(n10), .Q(
        ALU_reg[22]) );
  DFFR_X1 \ALU_reg_reg[23]  ( .D(ALU_exeout[23]), .CK(CLK), .RN(n10), .Q(
        ALU_reg[23]) );
  DFFR_X1 \ALU_reg_reg[24]  ( .D(ALU_exeout[24]), .CK(CLK), .RN(n10), .Q(
        ALU_reg[24]) );
  DFFR_X1 \ALU_reg_reg[25]  ( .D(ALU_exeout[25]), .CK(CLK), .RN(n10), .Q(
        ALU_reg[25]) );
  DFFR_X1 \ALU_reg_reg[26]  ( .D(ALU_exeout[26]), .CK(CLK), .RN(n10), .Q(
        ALU_reg[26]) );
  DFFR_X1 \ALU_reg_reg[27]  ( .D(ALU_exeout[27]), .CK(CLK), .RN(n10), .Q(
        ALU_reg[27]) );
  DFFR_X1 \ALU_reg_reg[28]  ( .D(ALU_exeout[28]), .CK(CLK), .RN(n9), .Q(
        ALU_reg[28]) );
  DFFR_X1 \ALU_reg_reg[29]  ( .D(ALU_exeout[29]), .CK(CLK), .RN(n9), .Q(
        ALU_reg[29]) );
  DFFR_X1 \ALU_reg_reg[30]  ( .D(ALU_exeout[30]), .CK(CLK), .RN(n9), .Q(
        ALU_reg[30]) );
  DFFR_X1 \ALU_reg_reg[31]  ( .D(ALU_exeout[31]), .CK(CLK), .RN(n9), .Q(
        ALU_reg[31]) );
  DFFR_X1 \RD_regwb_reg[0]  ( .D(RD_memout[0]), .CK(CLK), .RN(n9), .Q(
        RD_regwb[0]) );
  DFFR_X1 \RD_regwb_reg[1]  ( .D(RD_memout[1]), .CK(CLK), .RN(n9), .Q(
        RD_regwb[1]) );
  DFFR_X1 \RD_regwb_reg[2]  ( .D(RD_memout[2]), .CK(CLK), .RN(n9), .Q(
        RD_regwb[2]) );
  DFFR_X1 \RD_regwb_reg[3]  ( .D(RD_memout[3]), .CK(CLK), .RN(n9), .Q(
        RD_regwb[3]) );
  DFFR_X1 \RD_regwb_reg[4]  ( .D(RD_memout[4]), .CK(CLK), .RN(n9), .Q(
        RD_regwb[4]) );
  DFFR_X1 \ALU_regmem_reg[1]  ( .D(ALU_memout[1]), .CK(CLK), .RN(n9), .Q(
        ALU_regmem[1]) );
  DFFR_X1 \ALU_regmem_reg[2]  ( .D(ALU_memout[2]), .CK(CLK), .RN(n9), .Q(
        ALU_regmem[2]) );
  DFFR_X1 \ALU_regmem_reg[3]  ( .D(ALU_memout[3]), .CK(CLK), .RN(n9), .Q(
        ALU_regmem[3]) );
  DFFR_X1 \ALU_regmem_reg[4]  ( .D(ALU_memout[4]), .CK(CLK), .RN(n9), .Q(
        ALU_regmem[4]) );
  DFFR_X1 \ALU_regmem_reg[5]  ( .D(ALU_memout[5]), .CK(CLK), .RN(n9), .Q(
        ALU_regmem[5]) );
  DFFR_X1 \ALU_regmem_reg[6]  ( .D(ALU_memout[6]), .CK(CLK), .RN(n9), .Q(
        ALU_regmem[6]) );
  DFFR_X1 \ALU_regmem_reg[7]  ( .D(ALU_memout[7]), .CK(CLK), .RN(n9), .Q(
        ALU_regmem[7]) );
  DFFR_X1 \ALU_regmem_reg[8]  ( .D(ALU_memout[8]), .CK(CLK), .RN(n9), .Q(
        ALU_regmem[8]) );
  DFFR_X1 \ALU_regmem_reg[9]  ( .D(ALU_memout[9]), .CK(CLK), .RN(n9), .Q(
        ALU_regmem[9]) );
  DFFR_X1 \ALU_regmem_reg[10]  ( .D(ALU_memout[10]), .CK(CLK), .RN(n9), .Q(
        ALU_regmem[10]) );
  DFFR_X1 \ALU_regmem_reg[11]  ( .D(ALU_memout[11]), .CK(CLK), .RN(n9), .Q(
        ALU_regmem[11]) );
  DFFR_X1 \ALU_regmem_reg[12]  ( .D(ALU_memout[12]), .CK(CLK), .RN(n9), .Q(
        ALU_regmem[12]) );
  DFFR_X1 \ALU_regmem_reg[13]  ( .D(ALU_memout[13]), .CK(CLK), .RN(n9), .Q(
        ALU_regmem[13]) );
  DFFR_X1 \ALU_regmem_reg[14]  ( .D(ALU_memout[14]), .CK(CLK), .RN(n9), .Q(
        ALU_regmem[14]) );
  DFFR_X1 \ALU_regmem_reg[15]  ( .D(ALU_memout[15]), .CK(CLK), .RN(n9), .Q(
        ALU_regmem[15]) );
  DFFR_X1 \ALU_regmem_reg[16]  ( .D(ALU_memout[16]), .CK(CLK), .RN(n9), .Q(
        ALU_regmem[16]) );
  DFFR_X1 \ALU_regmem_reg[17]  ( .D(ALU_memout[17]), .CK(CLK), .RN(n9), .Q(
        ALU_regmem[17]) );
  DFFR_X1 \ALU_regmem_reg[18]  ( .D(ALU_memout[18]), .CK(CLK), .RN(n9), .Q(
        ALU_regmem[18]) );
  DFFR_X1 \ALU_regmem_reg[19]  ( .D(ALU_memout[19]), .CK(CLK), .RN(n9), .Q(
        ALU_regmem[19]) );
  DFFR_X1 \ALU_regmem_reg[20]  ( .D(ALU_memout[20]), .CK(CLK), .RN(n9), .Q(
        ALU_regmem[20]) );
  DFFR_X1 \ALU_regmem_reg[21]  ( .D(ALU_memout[21]), .CK(CLK), .RN(n9), .Q(
        ALU_regmem[21]) );
  DFFR_X1 \ALU_regmem_reg[22]  ( .D(ALU_memout[22]), .CK(CLK), .RN(n9), .Q(
        ALU_regmem[22]) );
  DFFR_X1 \ALU_regmem_reg[23]  ( .D(ALU_memout[23]), .CK(CLK), .RN(n9), .Q(
        ALU_regmem[23]) );
  DFFR_X1 \ALU_regmem_reg[24]  ( .D(ALU_memout[24]), .CK(CLK), .RN(n9), .Q(
        ALU_regmem[24]) );
  DFFR_X1 \ALU_regmem_reg[25]  ( .D(ALU_memout[25]), .CK(CLK), .RN(n10), .Q(
        ALU_regmem[25]) );
  DFFR_X1 \ALU_regmem_reg[26]  ( .D(ALU_memout[26]), .CK(CLK), .RN(n9), .Q(
        ALU_regmem[26]) );
  DFFR_X1 \ALU_regmem_reg[27]  ( .D(ALU_memout[27]), .CK(CLK), .RN(n9), .Q(
        ALU_regmem[27]) );
  DFFR_X1 \ALU_regmem_reg[28]  ( .D(ALU_memout[28]), .CK(CLK), .RN(n9), .Q(
        ALU_regmem[28]) );
  DFFR_X1 \ALU_regmem_reg[29]  ( .D(ALU_memout[29]), .CK(CLK), .RN(n9), .Q(
        ALU_regmem[29]) );
  DFFR_X1 \ALU_regmem_reg[30]  ( .D(ALU_memout[30]), .CK(CLK), .RN(n9), .Q(
        ALU_regmem[30]) );
  DFFR_X1 \ALU_regmem_reg[31]  ( .D(ALU_memout[31]), .CK(CLK), .RN(n9), .Q(
        ALU_regmem[31]) );
  DFFR_X1 \LMD_reg_reg[0]  ( .D(mem_out[0]), .CK(CLK), .RN(n9), .Q(LMD_reg[0])
         );
  DFFR_X1 \LMD_reg_reg[1]  ( .D(mem_out[1]), .CK(CLK), .RN(n9), .Q(LMD_reg[1])
         );
  DFFR_X1 \LMD_reg_reg[2]  ( .D(mem_out[2]), .CK(CLK), .RN(n9), .Q(LMD_reg[2])
         );
  DFFR_X1 \LMD_reg_reg[3]  ( .D(mem_out[3]), .CK(CLK), .RN(n8), .Q(LMD_reg[3])
         );
  DFFR_X1 \LMD_reg_reg[4]  ( .D(mem_out[4]), .CK(CLK), .RN(n8), .Q(LMD_reg[4])
         );
  DFFR_X1 \LMD_reg_reg[5]  ( .D(mem_out[5]), .CK(CLK), .RN(n8), .Q(LMD_reg[5])
         );
  DFFR_X1 \LMD_reg_reg[6]  ( .D(mem_out[6]), .CK(CLK), .RN(n8), .Q(LMD_reg[6])
         );
  DFFR_X1 \LMD_reg_reg[7]  ( .D(mem_out[7]), .CK(CLK), .RN(n8), .Q(LMD_reg[7])
         );
  DFFR_X1 \LMD_reg_reg[8]  ( .D(mem_out[8]), .CK(CLK), .RN(n8), .Q(LMD_reg[8])
         );
  DFFR_X1 \LMD_reg_reg[9]  ( .D(mem_out[9]), .CK(CLK), .RN(n8), .Q(LMD_reg[9])
         );
  DFFR_X1 \LMD_reg_reg[10]  ( .D(mem_out[10]), .CK(CLK), .RN(n8), .Q(
        LMD_reg[10]) );
  DFFR_X1 \LMD_reg_reg[11]  ( .D(mem_out[11]), .CK(CLK), .RN(n8), .Q(
        LMD_reg[11]) );
  DFFR_X1 \LMD_reg_reg[12]  ( .D(mem_out[12]), .CK(CLK), .RN(n8), .Q(
        LMD_reg[12]) );
  DFFR_X1 \LMD_reg_reg[13]  ( .D(mem_out[13]), .CK(CLK), .RN(n8), .Q(
        LMD_reg[13]) );
  DFFR_X1 \LMD_reg_reg[14]  ( .D(mem_out[14]), .CK(CLK), .RN(n8), .Q(
        LMD_reg[14]) );
  DFFR_X1 \LMD_reg_reg[15]  ( .D(mem_out[15]), .CK(CLK), .RN(n8), .Q(
        LMD_reg[15]) );
  DFFR_X1 \LMD_reg_reg[16]  ( .D(mem_out[16]), .CK(CLK), .RN(n8), .Q(
        LMD_reg[16]) );
  DFFR_X1 \LMD_reg_reg[17]  ( .D(mem_out[17]), .CK(CLK), .RN(n8), .Q(
        LMD_reg[17]) );
  DFFR_X1 \LMD_reg_reg[18]  ( .D(mem_out[18]), .CK(CLK), .RN(n8), .Q(
        LMD_reg[18]) );
  DFFR_X1 \LMD_reg_reg[19]  ( .D(mem_out[19]), .CK(CLK), .RN(n8), .Q(
        LMD_reg[19]) );
  DFFR_X1 \LMD_reg_reg[20]  ( .D(mem_out[20]), .CK(CLK), .RN(n8), .Q(
        LMD_reg[20]) );
  DFFR_X1 \LMD_reg_reg[21]  ( .D(mem_out[21]), .CK(CLK), .RN(n8), .Q(
        LMD_reg[21]) );
  DFFR_X1 \LMD_reg_reg[22]  ( .D(mem_out[22]), .CK(CLK), .RN(n8), .Q(
        LMD_reg[22]) );
  DFFR_X1 \LMD_reg_reg[23]  ( .D(mem_out[23]), .CK(CLK), .RN(n8), .Q(
        LMD_reg[23]) );
  DFFR_X1 \LMD_reg_reg[24]  ( .D(mem_out[24]), .CK(CLK), .RN(n8), .Q(
        LMD_reg[24]) );
  DFFR_X1 \LMD_reg_reg[25]  ( .D(mem_out[25]), .CK(CLK), .RN(n8), .Q(
        LMD_reg[25]) );
  DFFR_X1 \LMD_reg_reg[26]  ( .D(mem_out[26]), .CK(CLK), .RN(n8), .Q(
        LMD_reg[26]) );
  DFFR_X1 \LMD_reg_reg[27]  ( .D(mem_out[27]), .CK(CLK), .RN(n8), .Q(
        LMD_reg[27]) );
  DFFR_X1 \LMD_reg_reg[28]  ( .D(mem_out[28]), .CK(CLK), .RN(n8), .Q(
        LMD_reg[28]) );
  DFFR_X1 \LMD_reg_reg[29]  ( .D(mem_out[29]), .CK(CLK), .RN(n8), .Q(
        LMD_reg[29]) );
  DFFR_X1 \LMD_reg_reg[30]  ( .D(mem_out[30]), .CK(CLK), .RN(n8), .Q(
        LMD_reg[30]) );
  DFFR_X1 \LMD_reg_reg[31]  ( .D(mem_out[31]), .CK(CLK), .RN(n8), .Q(
        LMD_reg[31]) );
  MUX21_GENERIC_NBIT32_0 MUX ( .A(NPC_fetchout), .B(s_NPC_jump), .SEL(
        flag_signal), .Y(PC_muxout) );
  FETCH fetch_stage ( .PC(PC_reg), .hazard_PC(hazard_NPC), .PC_sel(
        hazard_NPC_sel), .IRAM_addr(IRAM_addr), .NPC(NPC_fetchout) );
  MUX21_GENERIC_NBIT32_5 NOP_MUX ( .A(instr), .B({1'b0, 1'b1, 1'b0, 1'b1, 1'b0, 
        1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .SEL(flag_signal), .Y(NOP_MUX_OUT) );
  DEC dec_stage ( .instr(IR_reg), .RST(n4), .RFdata_in(WB_data), .RFWA(
        RD_regwb), .NPC_in(NPC_reg), .EXE_RD(RD_regexe), .Ld(Ld), .ALU_regout(
        ALU_reg), .MEM_RD(RD_regmem), .WB_RD(RD_regwb), .RD_inmul(s_RD_inmul), 
        .flag_structHzd(s_flag_structHzd), .flag_ismul(s_flag_ismul), .RF1(RF1), .RF2(RF2), .WF1(WF1), .EN1(EN1), .opcode(opcode), .func(func), .IMM(
        IMM_decout), .RA(RA_decout), .RB(RB_decout), .RSA(RSA_decout), .RSB(
        RSB_decout), .RD(RD_decout), .stall_NPC(hazard_NPC), .PC_sel(
        hazard_NPC_sel), .dec_flag(flag_signal), .NPC_jump(s_NPC_jump) );
  EXE exe_stage ( .CLK(CLK), .RST(n4), .IMM(Imm_reg), .RA(RA_reg), .RB(RB_reg), 
        .WA(RD_regexe), .RSA(RSA_reg), .RSB(RSB_reg), .ALU_outmem(ALU_reg), 
        .WB_out(WB_data), .MEM_RD(RD_regmem), .WB_RD(RD_regwb), .LD_EN(EN3), 
        .WB_EN(WF1), .S1(S1), .S2(S2), .ALU3(ALU3), .ALU2(ALU2), .ALU1(ALU1), 
        .ALU0(ALU0), .SN(SN), .RD_inmul(s_RD_inmul), .flag_structHzd(
        s_flag_structHzd), .flag_ismul(s_flag_ismul), .OVF(OVF), .\output (
        ALU_exeout), .ME(ME_exeout), .WAout(RD_exeout) );
  MEM_MEMORY_SIZE128 mem_stage ( .CLK(CLK), .RST(n12), .ALUout(ALU_reg), 
        .MEout(ME_reg), .RDin(RD_regmem), .DRAM_data_out(DRAM_data_out), .LnS(
        LnS), .Wrd(Wrd), .BHU1(BHU1), .BHU0(BHU0), .EN3(EN3), .DRAM_addr(
        DRAM_addr), .DRAM_data_in(DRAM_data_in), .MMU_out(MMU_out), .\output (
        mem_out), .alu_out(ALU_memout), .RDout(RD_memout) );
  WB wb_stage ( .mem_out(LMD_reg), .alu_out(ALU_regmem), .S3(S3), .\output (
        WB_data) );
  DFFS_X2 \IR_reg_reg[30]  ( .D(NOP_MUX_OUT[30]), .CK(CLK), .SN(n12), .Q(
        IR_reg[30]) );
  DFFS_X1 \IR_reg_reg[28]  ( .D(NOP_MUX_OUT[28]), .CK(CLK), .SN(n12), .Q(
        IR_reg[28]) );
  BUF_X2 U3 ( .A(n2), .Z(n9) );
  BUF_X2 U4 ( .A(n3), .Z(n10) );
  BUF_X2 U5 ( .A(n3), .Z(n11) );
  BUF_X2 U6 ( .A(n1), .Z(n5) );
  BUF_X2 U7 ( .A(n1), .Z(n6) );
  BUF_X2 U8 ( .A(n2), .Z(n7) );
  BUF_X2 U9 ( .A(n2), .Z(n8) );
  BUF_X2 U10 ( .A(n1), .Z(n4) );
  BUF_X1 U11 ( .A(n3), .Z(n12) );
  BUF_X1 U12 ( .A(RST), .Z(n1) );
  BUF_X1 U13 ( .A(RST), .Z(n3) );
  BUF_X1 U14 ( .A(RST), .Z(n2) );
endmodule


module DLX_MEM_SIZE128_WORD_size32_NREG32 ( CLK, RST, from_DRAM_data, 
        IRAM_data, DRAM_addr, IRAM_addr, to_DRAM_data, DRAM_EN, DRAM_LnS, 
        MMU_out );
  input [31:0] from_DRAM_data;
  input [31:0] IRAM_data;
  output [8:0] DRAM_addr;
  output [7:0] IRAM_addr;
  output [31:0] to_DRAM_data;
  output [1:0] MMU_out;
  input CLK, RST;
  output DRAM_EN, DRAM_LnS;
  wire   s_RF1, s_RF2, s_EN1, s_S1, s_S2, s_ALU3, s_ALU2, s_ALU1, s_ALU0, s_SN,
         s_Wrd, s_BHU1, s_BHU0, s_S3, s_WF1, s_Ld;
  wire   [5:0] s_opcode;
  wire   [10:0] s_func;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23;

  hardwired_CU control_unit ( .clk(CLK), .rst(RST), .opcode(s_opcode), .func(
        s_func), .RF1(s_RF1), .RF2(s_RF2), .EN1(s_EN1), .S1(s_S1), .S2(s_S2), 
        .ALU3(s_ALU3), .ALU2(s_ALU2), .ALU1(s_ALU1), .ALU0(s_ALU0), .SN(s_SN), 
        .LnS(DRAM_LnS), .Wrd(s_Wrd), .BHU1(s_BHU1), .BHU0(s_BHU0), .EN3(
        DRAM_EN), .S3(s_S3), .WF1(s_WF1), .Ld(s_Ld) );
  DataPath_MEM_SIZE128_WORD_size32_NREG32 data_path ( .CLK(CLK), .RST(RST), 
        .RF1(s_RF1), .RF2(s_RF2), .EN1(s_EN1), .S1(s_S1), .S2(s_S2), .ALU3(
        s_ALU3), .ALU2(s_ALU2), .ALU1(s_ALU1), .ALU0(s_ALU0), .SN(s_SN), .LnS(
        DRAM_LnS), .BHU1(s_BHU1), .BHU0(s_BHU0), .Wrd(s_Wrd), .EN3(DRAM_EN), 
        .S3(s_S3), .WF1(s_WF1), .Ld(s_Ld), .instr(IRAM_data), .IRAM_addr({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, IRAM_addr}), 
        .DRAM_data_out(from_DRAM_data), .MMU_out(MMU_out), .DRAM_addr(
        DRAM_addr), .DRAM_data_in(to_DRAM_data), .opcode(s_opcode), .func(
        s_func) );
endmodule

