
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32 is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FETCH_DW01_add_0 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end FETCH_DW01_add_0;

architecture SYN_rpl of FETCH_DW01_add_0 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, SUM_26_port, 
      SUM_27_port, SUM_30_port, SUM_29_port, SUM_28_port, SUM_25_port, 
      SUM_24_port, SUM_23_port, SUM_22_port, SUM_21_port, SUM_20_port, 
      SUM_31_port, SUM_10_port, SUM_11_port, SUM_19_port, SUM_18_port, 
      SUM_17_port, SUM_16_port, SUM_15_port, SUM_14_port, SUM_13_port, 
      SUM_12_port, SUM_9_port, SUM_3_port, SUM_4_port, SUM_8_port, SUM_7_port, 
      SUM_6_port, SUM_5_port, n57, SUM_2_port : std_logic;

begin
   SUM <= ( SUM_31_port, SUM_30_port, SUM_29_port, SUM_28_port, SUM_27_port, 
      SUM_26_port, SUM_25_port, SUM_24_port, SUM_23_port, SUM_22_port, 
      SUM_21_port, SUM_20_port, SUM_19_port, SUM_18_port, SUM_17_port, 
      SUM_16_port, SUM_15_port, SUM_14_port, SUM_13_port, SUM_12_port, 
      SUM_11_port, SUM_10_port, SUM_9_port, SUM_8_port, SUM_7_port, SUM_6_port,
      SUM_5_port, SUM_4_port, SUM_3_port, SUM_2_port, A(1), A(0) );
   
   U1 : AND2_X1 port map( A1 => A(3), A2 => A(2), ZN => n1);
   U2 : AND2_X1 port map( A1 => A(10), A2 => n12, ZN => n2);
   U3 : AND2_X1 port map( A1 => A(26), A2 => n7, ZN => n3);
   U4 : AND2_X1 port map( A1 => A(6), A2 => n27, ZN => n4);
   U5 : AND2_X1 port map( A1 => A(7), A2 => n4, ZN => n5);
   U6 : AND2_X1 port map( A1 => A(24), A2 => n25, ZN => n6);
   U7 : AND2_X1 port map( A1 => A(25), A2 => n6, ZN => n7);
   U8 : AND2_X1 port map( A1 => A(27), A2 => n3, ZN => n8);
   U9 : AND2_X1 port map( A1 => A(28), A2 => n8, ZN => n9);
   U10 : AND2_X1 port map( A1 => A(29), A2 => n9, ZN => n10);
   U11 : AND2_X1 port map( A1 => A(8), A2 => n5, ZN => n11);
   U12 : AND2_X1 port map( A1 => A(9), A2 => n11, ZN => n12);
   U13 : AND2_X1 port map( A1 => A(11), A2 => n2, ZN => n13);
   U14 : AND2_X1 port map( A1 => A(12), A2 => n13, ZN => n14);
   U15 : AND2_X1 port map( A1 => A(13), A2 => n14, ZN => n15);
   U16 : AND2_X1 port map( A1 => A(14), A2 => n15, ZN => n16);
   U17 : AND2_X1 port map( A1 => A(15), A2 => n16, ZN => n17);
   U18 : AND2_X1 port map( A1 => A(16), A2 => n17, ZN => n18);
   U19 : AND2_X1 port map( A1 => A(17), A2 => n18, ZN => n19);
   U20 : AND2_X1 port map( A1 => A(18), A2 => n19, ZN => n20);
   U21 : AND2_X1 port map( A1 => A(19), A2 => n20, ZN => n21);
   U22 : AND2_X1 port map( A1 => A(20), A2 => n21, ZN => n22);
   U23 : AND2_X1 port map( A1 => A(21), A2 => n22, ZN => n23);
   U24 : AND2_X1 port map( A1 => A(22), A2 => n23, ZN => n24);
   U25 : AND2_X1 port map( A1 => A(23), A2 => n24, ZN => n25);
   U26 : AND2_X1 port map( A1 => A(4), A2 => n1, ZN => n26);
   U27 : AND2_X1 port map( A1 => A(5), A2 => n26, ZN => n27);
   U28 : NAND2_X1 port map( A1 => A(30), A2 => n10, ZN => n57);
   U29 : XOR2_X1 port map( A => A(26), B => n7, Z => SUM_26_port);
   U30 : XOR2_X1 port map( A => A(27), B => n3, Z => SUM_27_port);
   U31 : XOR2_X1 port map( A => A(30), B => n10, Z => SUM_30_port);
   U32 : XOR2_X1 port map( A => A(29), B => n9, Z => SUM_29_port);
   U33 : XOR2_X1 port map( A => A(28), B => n8, Z => SUM_28_port);
   U34 : XOR2_X1 port map( A => A(25), B => n6, Z => SUM_25_port);
   U35 : XOR2_X1 port map( A => A(24), B => n25, Z => SUM_24_port);
   U36 : XOR2_X1 port map( A => A(23), B => n24, Z => SUM_23_port);
   U37 : XOR2_X1 port map( A => A(22), B => n23, Z => SUM_22_port);
   U38 : XOR2_X1 port map( A => A(21), B => n22, Z => SUM_21_port);
   U39 : XOR2_X1 port map( A => A(20), B => n21, Z => SUM_20_port);
   U40 : XNOR2_X1 port map( A => A(31), B => n57, ZN => SUM_31_port);
   U41 : XOR2_X1 port map( A => A(10), B => n12, Z => SUM_10_port);
   U42 : XOR2_X1 port map( A => A(11), B => n2, Z => SUM_11_port);
   U43 : XOR2_X1 port map( A => A(19), B => n20, Z => SUM_19_port);
   U44 : XOR2_X1 port map( A => A(18), B => n19, Z => SUM_18_port);
   U45 : XOR2_X1 port map( A => A(17), B => n18, Z => SUM_17_port);
   U46 : XOR2_X1 port map( A => A(16), B => n17, Z => SUM_16_port);
   U47 : XOR2_X1 port map( A => A(15), B => n16, Z => SUM_15_port);
   U48 : XOR2_X1 port map( A => A(14), B => n15, Z => SUM_14_port);
   U49 : XOR2_X1 port map( A => A(13), B => n14, Z => SUM_13_port);
   U50 : XOR2_X1 port map( A => A(12), B => n13, Z => SUM_12_port);
   U51 : XOR2_X1 port map( A => A(9), B => n11, Z => SUM_9_port);
   U52 : INV_X1 port map( A => A(2), ZN => SUM_2_port);
   U53 : XOR2_X1 port map( A => A(3), B => A(2), Z => SUM_3_port);
   U54 : XOR2_X1 port map( A => A(4), B => n1, Z => SUM_4_port);
   U55 : XOR2_X1 port map( A => A(8), B => n5, Z => SUM_8_port);
   U56 : XOR2_X1 port map( A => A(7), B => n4, Z => SUM_7_port);
   U57 : XOR2_X1 port map( A => A(6), B => n27, Z => SUM_6_port);
   U58 : XOR2_X1 port map( A => A(5), B => n26, Z => SUM_5_port);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity 
   stall_detection_unit_op_code_size6_func_size11_PC_reg_size32_reg_file_size32_DW01_sub_3 
   is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end 
   stall_detection_unit_op_code_size6_func_size11_PC_reg_size32_reg_file_size32_DW01_sub_3;

architecture SYN_rpl of 
   stall_detection_unit_op_code_size6_func_size11_PC_reg_size32_reg_file_size32_DW01_sub_3 
   is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal DIFF_31_port, DIFF_30_port, DIFF_29_port, DIFF_28_port, DIFF_27_port,
      DIFF_26_port, DIFF_25_port, DIFF_24_port, DIFF_23_port, DIFF_22_port, 
      DIFF_21_port, DIFF_20_port, DIFF_19_port, DIFF_18_port, DIFF_17_port, 
      DIFF_16_port, DIFF_15_port, DIFF_14_port, DIFF_13_port, DIFF_12_port, 
      DIFF_11_port, DIFF_10_port, DIFF_9_port, DIFF_8_port, DIFF_7_port, 
      DIFF_6_port, DIFF_5_port, DIFF_4_port, DIFF_3_port, carry_31_port, 
      carry_30_port, carry_29_port, carry_28_port, carry_27_port, carry_26_port
      , carry_25_port, carry_24_port, carry_23_port, carry_22_port, 
      carry_21_port, carry_20_port, carry_19_port, carry_18_port, carry_17_port
      , carry_16_port, carry_15_port, carry_14_port, carry_13_port, 
      carry_12_port, carry_11_port, carry_10_port, carry_9_port, carry_8_port, 
      carry_7_port, carry_6_port, carry_5_port, carry_4_port, n1, n2, 
      DIFF_2_port : std_logic;

begin
   DIFF <= ( DIFF_31_port, DIFF_30_port, DIFF_29_port, DIFF_28_port, 
      DIFF_27_port, DIFF_26_port, DIFF_25_port, DIFF_24_port, DIFF_23_port, 
      DIFF_22_port, DIFF_21_port, DIFF_20_port, DIFF_19_port, DIFF_18_port, 
      DIFF_17_port, DIFF_16_port, DIFF_15_port, DIFF_14_port, DIFF_13_port, 
      DIFF_12_port, DIFF_11_port, DIFF_10_port, DIFF_9_port, DIFF_8_port, 
      DIFF_7_port, DIFF_6_port, DIFF_5_port, DIFF_4_port, DIFF_3_port, 
      DIFF_2_port, A(1), A(0) );
   
   U1 : XNOR2_X1 port map( A => A(10), B => carry_10_port, ZN => DIFF_10_port);
   U2 : XNOR2_X1 port map( A => A(11), B => carry_11_port, ZN => DIFF_11_port);
   U3 : XNOR2_X1 port map( A => A(13), B => carry_13_port, ZN => DIFF_13_port);
   U4 : XNOR2_X1 port map( A => A(15), B => carry_15_port, ZN => DIFF_15_port);
   U5 : XNOR2_X1 port map( A => A(16), B => carry_16_port, ZN => DIFF_16_port);
   U6 : XNOR2_X1 port map( A => A(17), B => carry_17_port, ZN => DIFF_17_port);
   U7 : XNOR2_X1 port map( A => A(18), B => carry_18_port, ZN => DIFF_18_port);
   U8 : XNOR2_X1 port map( A => A(19), B => carry_19_port, ZN => DIFF_19_port);
   U9 : XNOR2_X1 port map( A => A(5), B => carry_5_port, ZN => DIFF_5_port);
   U10 : XNOR2_X1 port map( A => A(8), B => carry_8_port, ZN => DIFF_8_port);
   U11 : XNOR2_X1 port map( A => A(9), B => carry_9_port, ZN => DIFF_9_port);
   U12 : XNOR2_X1 port map( A => A(20), B => carry_20_port, ZN => DIFF_20_port)
                           ;
   U13 : XNOR2_X1 port map( A => A(21), B => carry_21_port, ZN => DIFF_21_port)
                           ;
   U14 : XNOR2_X1 port map( A => A(22), B => carry_22_port, ZN => DIFF_22_port)
                           ;
   U15 : XNOR2_X1 port map( A => A(23), B => carry_23_port, ZN => DIFF_23_port)
                           ;
   U16 : XNOR2_X1 port map( A => A(24), B => carry_24_port, ZN => DIFF_24_port)
                           ;
   U17 : XNOR2_X1 port map( A => A(25), B => carry_25_port, ZN => DIFF_25_port)
                           ;
   U18 : XNOR2_X1 port map( A => A(26), B => carry_26_port, ZN => DIFF_26_port)
                           ;
   U19 : XNOR2_X1 port map( A => A(27), B => carry_27_port, ZN => DIFF_27_port)
                           ;
   U20 : XNOR2_X1 port map( A => A(28), B => carry_28_port, ZN => DIFF_28_port)
                           ;
   U21 : XNOR2_X1 port map( A => A(29), B => carry_29_port, ZN => DIFF_29_port)
                           ;
   U22 : XNOR2_X1 port map( A => A(30), B => carry_30_port, ZN => DIFF_30_port)
                           ;
   U23 : XNOR2_X1 port map( A => A(7), B => carry_7_port, ZN => DIFF_7_port);
   U24 : INV_X1 port map( A => A(2), ZN => DIFF_2_port);
   U25 : XNOR2_X1 port map( A => A(3), B => A(2), ZN => DIFF_3_port);
   U26 : XNOR2_X1 port map( A => A(4), B => carry_4_port, ZN => DIFF_4_port);
   U27 : XNOR2_X1 port map( A => A(12), B => carry_12_port, ZN => DIFF_12_port)
                           ;
   U28 : XNOR2_X1 port map( A => A(14), B => carry_14_port, ZN => DIFF_14_port)
                           ;
   U29 : XNOR2_X1 port map( A => A(6), B => carry_6_port, ZN => DIFF_6_port);
   U30 : OR2_X1 port map( A1 => A(3), A2 => A(2), ZN => carry_4_port);
   U31 : XNOR2_X1 port map( A => A(31), B => carry_31_port, ZN => DIFF_31_port)
                           ;
   U32 : NAND2_X1 port map( A1 => n1, A2 => n2, ZN => carry_31_port);
   U33 : INV_X1 port map( A => A(30), ZN => n1);
   U34 : INV_X1 port map( A => carry_30_port, ZN => n2);
   U35 : OR2_X1 port map( A1 => A(4), A2 => carry_4_port, ZN => carry_5_port);
   U36 : OR2_X1 port map( A1 => A(7), A2 => carry_7_port, ZN => carry_8_port);
   U37 : OR2_X1 port map( A1 => A(8), A2 => carry_8_port, ZN => carry_9_port);
   U38 : OR2_X1 port map( A1 => A(9), A2 => carry_9_port, ZN => carry_10_port);
   U39 : OR2_X1 port map( A1 => A(10), A2 => carry_10_port, ZN => carry_11_port
                           );
   U40 : OR2_X1 port map( A1 => A(11), A2 => carry_11_port, ZN => carry_12_port
                           );
   U41 : OR2_X1 port map( A1 => A(12), A2 => carry_12_port, ZN => carry_13_port
                           );
   U42 : OR2_X1 port map( A1 => A(13), A2 => carry_13_port, ZN => carry_14_port
                           );
   U43 : OR2_X1 port map( A1 => A(14), A2 => carry_14_port, ZN => carry_15_port
                           );
   U44 : OR2_X1 port map( A1 => A(15), A2 => carry_15_port, ZN => carry_16_port
                           );
   U45 : OR2_X1 port map( A1 => A(16), A2 => carry_16_port, ZN => carry_17_port
                           );
   U46 : OR2_X1 port map( A1 => A(23), A2 => carry_23_port, ZN => carry_24_port
                           );
   U47 : OR2_X1 port map( A1 => A(24), A2 => carry_24_port, ZN => carry_25_port
                           );
   U48 : OR2_X1 port map( A1 => A(25), A2 => carry_25_port, ZN => carry_26_port
                           );
   U49 : OR2_X1 port map( A1 => A(26), A2 => carry_26_port, ZN => carry_27_port
                           );
   U50 : OR2_X1 port map( A1 => A(27), A2 => carry_27_port, ZN => carry_28_port
                           );
   U51 : OR2_X1 port map( A1 => A(28), A2 => carry_28_port, ZN => carry_29_port
                           );
   U52 : OR2_X1 port map( A1 => A(29), A2 => carry_29_port, ZN => carry_30_port
                           );
   U53 : OR2_X1 port map( A1 => A(5), A2 => carry_5_port, ZN => carry_6_port);
   U54 : OR2_X1 port map( A1 => A(6), A2 => carry_6_port, ZN => carry_7_port);
   U55 : OR2_X1 port map( A1 => A(17), A2 => carry_17_port, ZN => carry_18_port
                           );
   U56 : OR2_X1 port map( A1 => A(18), A2 => carry_18_port, ZN => carry_19_port
                           );
   U57 : OR2_X1 port map( A1 => A(19), A2 => carry_19_port, ZN => carry_20_port
                           );
   U58 : OR2_X1 port map( A1 => A(20), A2 => carry_20_port, ZN => carry_21_port
                           );
   U59 : OR2_X1 port map( A1 => A(21), A2 => carry_21_port, ZN => carry_22_port
                           );
   U60 : OR2_X1 port map( A1 => A(22), A2 => carry_22_port, ZN => carry_23_port
                           );

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity 
   stall_detection_unit_op_code_size6_func_size11_PC_reg_size32_reg_file_size32_DW01_sub_2 
   is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end 
   stall_detection_unit_op_code_size6_func_size11_PC_reg_size32_reg_file_size32_DW01_sub_2;

architecture SYN_rpl of 
   stall_detection_unit_op_code_size6_func_size11_PC_reg_size32_reg_file_size32_DW01_sub_2 
   is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal DIFF_31_port, DIFF_30_port, DIFF_29_port, DIFF_28_port, DIFF_27_port,
      DIFF_26_port, DIFF_25_port, DIFF_24_port, DIFF_23_port, DIFF_22_port, 
      DIFF_21_port, DIFF_20_port, DIFF_19_port, DIFF_18_port, DIFF_17_port, 
      DIFF_16_port, DIFF_15_port, DIFF_14_port, DIFF_13_port, DIFF_12_port, 
      DIFF_11_port, DIFF_10_port, DIFF_9_port, DIFF_8_port, DIFF_7_port, 
      DIFF_6_port, DIFF_5_port, DIFF_4_port, DIFF_3_port, DIFF_2_port, 
      carry_31_port, carry_30_port, carry_29_port, carry_28_port, carry_27_port
      , carry_26_port, carry_25_port, carry_24_port, carry_23_port, 
      carry_22_port, carry_21_port, carry_20_port, carry_19_port, carry_18_port
      , carry_17_port, carry_16_port, carry_15_port, carry_14_port, 
      carry_13_port, carry_12_port, carry_11_port, carry_10_port, carry_9_port,
      carry_8_port, carry_7_port, carry_6_port, carry_5_port, carry_4_port, 
      carry_3_port, n1, n2, n3 : std_logic;

begin
   DIFF <= ( DIFF_31_port, DIFF_30_port, DIFF_29_port, DIFF_28_port, 
      DIFF_27_port, DIFF_26_port, DIFF_25_port, DIFF_24_port, DIFF_23_port, 
      DIFF_22_port, DIFF_21_port, DIFF_20_port, DIFF_19_port, DIFF_18_port, 
      DIFF_17_port, DIFF_16_port, DIFF_15_port, DIFF_14_port, DIFF_13_port, 
      DIFF_12_port, DIFF_11_port, DIFF_10_port, DIFF_9_port, DIFF_8_port, 
      DIFF_7_port, DIFF_6_port, DIFF_5_port, DIFF_4_port, DIFF_3_port, 
      DIFF_2_port, A(1), A(0) );
   
   U1 : XNOR2_X1 port map( A => A(10), B => carry_10_port, ZN => DIFF_10_port);
   U2 : XNOR2_X1 port map( A => A(11), B => carry_11_port, ZN => DIFF_11_port);
   U3 : XNOR2_X1 port map( A => A(13), B => carry_13_port, ZN => DIFF_13_port);
   U4 : XNOR2_X1 port map( A => A(15), B => carry_15_port, ZN => DIFF_15_port);
   U5 : XNOR2_X1 port map( A => A(16), B => carry_16_port, ZN => DIFF_16_port);
   U6 : XNOR2_X1 port map( A => A(17), B => carry_17_port, ZN => DIFF_17_port);
   U7 : XNOR2_X1 port map( A => A(18), B => carry_18_port, ZN => DIFF_18_port);
   U8 : XNOR2_X1 port map( A => A(19), B => carry_19_port, ZN => DIFF_19_port);
   U9 : XNOR2_X1 port map( A => A(5), B => carry_5_port, ZN => DIFF_5_port);
   U10 : XNOR2_X1 port map( A => A(8), B => carry_8_port, ZN => DIFF_8_port);
   U11 : XNOR2_X1 port map( A => A(9), B => carry_9_port, ZN => DIFF_9_port);
   U12 : XNOR2_X1 port map( A => A(20), B => carry_20_port, ZN => DIFF_20_port)
                           ;
   U13 : XNOR2_X1 port map( A => A(21), B => carry_21_port, ZN => DIFF_21_port)
                           ;
   U14 : XNOR2_X1 port map( A => A(22), B => carry_22_port, ZN => DIFF_22_port)
                           ;
   U15 : XNOR2_X1 port map( A => A(23), B => carry_23_port, ZN => DIFF_23_port)
                           ;
   U16 : XNOR2_X1 port map( A => A(24), B => carry_24_port, ZN => DIFF_24_port)
                           ;
   U17 : XNOR2_X1 port map( A => A(25), B => carry_25_port, ZN => DIFF_25_port)
                           ;
   U18 : XNOR2_X1 port map( A => A(26), B => carry_26_port, ZN => DIFF_26_port)
                           ;
   U19 : XNOR2_X1 port map( A => A(27), B => carry_27_port, ZN => DIFF_27_port)
                           ;
   U20 : XNOR2_X1 port map( A => A(28), B => carry_28_port, ZN => DIFF_28_port)
                           ;
   U21 : XNOR2_X1 port map( A => A(29), B => carry_29_port, ZN => DIFF_29_port)
                           ;
   U22 : XNOR2_X1 port map( A => A(30), B => carry_30_port, ZN => DIFF_30_port)
                           ;
   U23 : XNOR2_X1 port map( A => A(7), B => carry_7_port, ZN => DIFF_7_port);
   U24 : XNOR2_X1 port map( A => n3, B => A(2), ZN => DIFF_2_port);
   U25 : XNOR2_X1 port map( A => A(3), B => carry_3_port, ZN => DIFF_3_port);
   U26 : XNOR2_X1 port map( A => A(4), B => carry_4_port, ZN => DIFF_4_port);
   U27 : XNOR2_X1 port map( A => A(12), B => carry_12_port, ZN => DIFF_12_port)
                           ;
   U28 : XNOR2_X1 port map( A => A(14), B => carry_14_port, ZN => DIFF_14_port)
                           ;
   U29 : XNOR2_X1 port map( A => A(6), B => carry_6_port, ZN => DIFF_6_port);
   U30 : XNOR2_X1 port map( A => A(31), B => carry_31_port, ZN => DIFF_31_port)
                           ;
   U31 : NAND2_X1 port map( A1 => n1, A2 => n2, ZN => carry_31_port);
   U32 : INV_X1 port map( A => A(30), ZN => n1);
   U33 : INV_X1 port map( A => carry_30_port, ZN => n2);
   U34 : OR2_X1 port map( A1 => n3, A2 => A(2), ZN => carry_3_port);
   U35 : OR2_X1 port map( A1 => A(3), A2 => carry_3_port, ZN => carry_4_port);
   U36 : OR2_X1 port map( A1 => A(4), A2 => carry_4_port, ZN => carry_5_port);
   U37 : OR2_X1 port map( A1 => A(5), A2 => carry_5_port, ZN => carry_6_port);
   U38 : OR2_X1 port map( A1 => A(6), A2 => carry_6_port, ZN => carry_7_port);
   U39 : OR2_X1 port map( A1 => A(7), A2 => carry_7_port, ZN => carry_8_port);
   U40 : OR2_X1 port map( A1 => A(8), A2 => carry_8_port, ZN => carry_9_port);
   U41 : OR2_X1 port map( A1 => A(9), A2 => carry_9_port, ZN => carry_10_port);
   U42 : OR2_X1 port map( A1 => A(10), A2 => carry_10_port, ZN => carry_11_port
                           );
   U43 : OR2_X1 port map( A1 => A(11), A2 => carry_11_port, ZN => carry_12_port
                           );
   U44 : OR2_X1 port map( A1 => A(12), A2 => carry_12_port, ZN => carry_13_port
                           );
   U45 : OR2_X1 port map( A1 => A(13), A2 => carry_13_port, ZN => carry_14_port
                           );
   U46 : OR2_X1 port map( A1 => A(14), A2 => carry_14_port, ZN => carry_15_port
                           );
   U47 : OR2_X1 port map( A1 => A(15), A2 => carry_15_port, ZN => carry_16_port
                           );
   U48 : OR2_X1 port map( A1 => A(16), A2 => carry_16_port, ZN => carry_17_port
                           );
   U49 : OR2_X1 port map( A1 => A(17), A2 => carry_17_port, ZN => carry_18_port
                           );
   U50 : OR2_X1 port map( A1 => A(18), A2 => carry_18_port, ZN => carry_19_port
                           );
   U51 : OR2_X1 port map( A1 => A(19), A2 => carry_19_port, ZN => carry_20_port
                           );
   U52 : OR2_X1 port map( A1 => A(20), A2 => carry_20_port, ZN => carry_21_port
                           );
   U53 : OR2_X1 port map( A1 => A(21), A2 => carry_21_port, ZN => carry_22_port
                           );
   U54 : OR2_X1 port map( A1 => A(22), A2 => carry_22_port, ZN => carry_23_port
                           );
   U55 : OR2_X1 port map( A1 => A(23), A2 => carry_23_port, ZN => carry_24_port
                           );
   U56 : OR2_X1 port map( A1 => A(24), A2 => carry_24_port, ZN => carry_25_port
                           );
   U57 : OR2_X1 port map( A1 => A(25), A2 => carry_25_port, ZN => carry_26_port
                           );
   U58 : OR2_X1 port map( A1 => A(26), A2 => carry_26_port, ZN => carry_27_port
                           );
   U59 : OR2_X1 port map( A1 => A(27), A2 => carry_27_port, ZN => carry_28_port
                           );
   U60 : OR2_X1 port map( A1 => A(28), A2 => carry_28_port, ZN => carry_29_port
                           );
   U61 : OR2_X1 port map( A1 => A(29), A2 => carry_29_port, ZN => carry_30_port
                           );
   U62 : INV_X1 port map( A => B(2), ZN => n3);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity 
   stall_detection_unit_op_code_size6_func_size11_PC_reg_size32_reg_file_size32_DW01_sub_1 
   is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end 
   stall_detection_unit_op_code_size6_func_size11_PC_reg_size32_reg_file_size32_DW01_sub_1;

architecture SYN_rpl of 
   stall_detection_unit_op_code_size6_func_size11_PC_reg_size32_reg_file_size32_DW01_sub_1 
   is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal DIFF_31_port, DIFF_30_port, DIFF_29_port, DIFF_28_port, DIFF_27_port,
      DIFF_26_port, DIFF_25_port, DIFF_24_port, DIFF_23_port, DIFF_22_port, 
      DIFF_21_port, DIFF_20_port, DIFF_19_port, DIFF_18_port, DIFF_17_port, 
      DIFF_16_port, DIFF_15_port, DIFF_14_port, DIFF_13_port, DIFF_12_port, 
      DIFF_11_port, DIFF_10_port, DIFF_9_port, DIFF_8_port, DIFF_7_port, 
      DIFF_6_port, DIFF_5_port, DIFF_4_port, DIFF_3_port, DIFF_2_port, 
      carry_31_port, carry_30_port, carry_29_port, carry_28_port, carry_27_port
      , carry_26_port, carry_25_port, carry_24_port, carry_23_port, 
      carry_22_port, carry_21_port, carry_20_port, carry_19_port, carry_18_port
      , carry_17_port, carry_16_port, carry_15_port, carry_14_port, 
      carry_13_port, carry_12_port, carry_11_port, carry_10_port, carry_9_port,
      carry_8_port, carry_7_port, carry_6_port, carry_5_port, carry_4_port, 
      carry_3_port, n1, n2, n3 : std_logic;

begin
   DIFF <= ( DIFF_31_port, DIFF_30_port, DIFF_29_port, DIFF_28_port, 
      DIFF_27_port, DIFF_26_port, DIFF_25_port, DIFF_24_port, DIFF_23_port, 
      DIFF_22_port, DIFF_21_port, DIFF_20_port, DIFF_19_port, DIFF_18_port, 
      DIFF_17_port, DIFF_16_port, DIFF_15_port, DIFF_14_port, DIFF_13_port, 
      DIFF_12_port, DIFF_11_port, DIFF_10_port, DIFF_9_port, DIFF_8_port, 
      DIFF_7_port, DIFF_6_port, DIFF_5_port, DIFF_4_port, DIFF_3_port, 
      DIFF_2_port, A(1), A(0) );
   
   U1 : INV_X1 port map( A => B(2), ZN => n3);
   U2 : INV_X1 port map( A => carry_30_port, ZN => n2);
   U3 : XNOR2_X1 port map( A => A(8), B => carry_8_port, ZN => DIFF_8_port);
   U4 : XNOR2_X1 port map( A => A(9), B => carry_9_port, ZN => DIFF_9_port);
   U5 : XNOR2_X1 port map( A => A(10), B => carry_10_port, ZN => DIFF_10_port);
   U6 : XNOR2_X1 port map( A => A(11), B => carry_11_port, ZN => DIFF_11_port);
   U7 : XNOR2_X1 port map( A => A(12), B => carry_12_port, ZN => DIFF_12_port);
   U8 : XNOR2_X1 port map( A => A(13), B => carry_13_port, ZN => DIFF_13_port);
   U9 : XNOR2_X1 port map( A => A(14), B => carry_14_port, ZN => DIFF_14_port);
   U10 : XNOR2_X1 port map( A => A(15), B => carry_15_port, ZN => DIFF_15_port)
                           ;
   U11 : XNOR2_X1 port map( A => A(3), B => carry_3_port, ZN => DIFF_3_port);
   U12 : XNOR2_X1 port map( A => A(4), B => carry_4_port, ZN => DIFF_4_port);
   U13 : XNOR2_X1 port map( A => A(5), B => carry_5_port, ZN => DIFF_5_port);
   U14 : XNOR2_X1 port map( A => A(6), B => carry_6_port, ZN => DIFF_6_port);
   U15 : XNOR2_X1 port map( A => A(7), B => carry_7_port, ZN => DIFF_7_port);
   U16 : XNOR2_X1 port map( A => A(16), B => carry_16_port, ZN => DIFF_16_port)
                           ;
   U17 : XNOR2_X1 port map( A => A(17), B => carry_17_port, ZN => DIFF_17_port)
                           ;
   U18 : XNOR2_X1 port map( A => A(18), B => carry_18_port, ZN => DIFF_18_port)
                           ;
   U19 : XNOR2_X1 port map( A => A(19), B => carry_19_port, ZN => DIFF_19_port)
                           ;
   U20 : XNOR2_X1 port map( A => A(20), B => carry_20_port, ZN => DIFF_20_port)
                           ;
   U21 : XNOR2_X1 port map( A => A(21), B => carry_21_port, ZN => DIFF_21_port)
                           ;
   U22 : XNOR2_X1 port map( A => A(22), B => carry_22_port, ZN => DIFF_22_port)
                           ;
   U23 : XNOR2_X1 port map( A => A(23), B => carry_23_port, ZN => DIFF_23_port)
                           ;
   U24 : XNOR2_X1 port map( A => A(24), B => carry_24_port, ZN => DIFF_24_port)
                           ;
   U25 : XNOR2_X1 port map( A => A(25), B => carry_25_port, ZN => DIFF_25_port)
                           ;
   U26 : XNOR2_X1 port map( A => A(26), B => carry_26_port, ZN => DIFF_26_port)
                           ;
   U27 : XNOR2_X1 port map( A => A(27), B => carry_27_port, ZN => DIFF_27_port)
                           ;
   U28 : XNOR2_X1 port map( A => A(28), B => carry_28_port, ZN => DIFF_28_port)
                           ;
   U29 : XNOR2_X1 port map( A => A(29), B => carry_29_port, ZN => DIFF_29_port)
                           ;
   U30 : XNOR2_X1 port map( A => A(30), B => carry_30_port, ZN => DIFF_30_port)
                           ;
   U31 : XNOR2_X1 port map( A => n3, B => A(2), ZN => DIFF_2_port);
   U32 : XNOR2_X1 port map( A => A(31), B => carry_31_port, ZN => DIFF_31_port)
                           ;
   U33 : NAND2_X1 port map( A1 => n1, A2 => n2, ZN => carry_31_port);
   U34 : INV_X1 port map( A => A(30), ZN => n1);
   U35 : OR2_X1 port map( A1 => n3, A2 => A(2), ZN => carry_3_port);
   U36 : OR2_X1 port map( A1 => A(3), A2 => carry_3_port, ZN => carry_4_port);
   U37 : OR2_X1 port map( A1 => A(4), A2 => carry_4_port, ZN => carry_5_port);
   U38 : OR2_X1 port map( A1 => A(5), A2 => carry_5_port, ZN => carry_6_port);
   U39 : OR2_X1 port map( A1 => A(6), A2 => carry_6_port, ZN => carry_7_port);
   U40 : OR2_X1 port map( A1 => A(7), A2 => carry_7_port, ZN => carry_8_port);
   U41 : OR2_X1 port map( A1 => A(8), A2 => carry_8_port, ZN => carry_9_port);
   U42 : OR2_X1 port map( A1 => A(9), A2 => carry_9_port, ZN => carry_10_port);
   U43 : OR2_X1 port map( A1 => A(10), A2 => carry_10_port, ZN => carry_11_port
                           );
   U44 : OR2_X1 port map( A1 => A(11), A2 => carry_11_port, ZN => carry_12_port
                           );
   U45 : OR2_X1 port map( A1 => A(12), A2 => carry_12_port, ZN => carry_13_port
                           );
   U46 : OR2_X1 port map( A1 => A(13), A2 => carry_13_port, ZN => carry_14_port
                           );
   U47 : OR2_X1 port map( A1 => A(14), A2 => carry_14_port, ZN => carry_15_port
                           );
   U48 : OR2_X1 port map( A1 => A(15), A2 => carry_15_port, ZN => carry_16_port
                           );
   U49 : OR2_X1 port map( A1 => A(16), A2 => carry_16_port, ZN => carry_17_port
                           );
   U50 : OR2_X1 port map( A1 => A(17), A2 => carry_17_port, ZN => carry_18_port
                           );
   U51 : OR2_X1 port map( A1 => A(18), A2 => carry_18_port, ZN => carry_19_port
                           );
   U52 : OR2_X1 port map( A1 => A(19), A2 => carry_19_port, ZN => carry_20_port
                           );
   U53 : OR2_X1 port map( A1 => A(20), A2 => carry_20_port, ZN => carry_21_port
                           );
   U54 : OR2_X1 port map( A1 => A(21), A2 => carry_21_port, ZN => carry_22_port
                           );
   U55 : OR2_X1 port map( A1 => A(22), A2 => carry_22_port, ZN => carry_23_port
                           );
   U56 : OR2_X1 port map( A1 => A(23), A2 => carry_23_port, ZN => carry_24_port
                           );
   U57 : OR2_X1 port map( A1 => A(24), A2 => carry_24_port, ZN => carry_25_port
                           );
   U58 : OR2_X1 port map( A1 => A(25), A2 => carry_25_port, ZN => carry_26_port
                           );
   U59 : OR2_X1 port map( A1 => A(26), A2 => carry_26_port, ZN => carry_27_port
                           );
   U60 : OR2_X1 port map( A1 => A(27), A2 => carry_27_port, ZN => carry_28_port
                           );
   U61 : OR2_X1 port map( A1 => A(28), A2 => carry_28_port, ZN => carry_29_port
                           );
   U62 : OR2_X1 port map( A1 => A(29), A2 => carry_29_port, ZN => carry_30_port
                           );

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity 
   stall_detection_unit_op_code_size6_func_size11_PC_reg_size32_reg_file_size32_DW01_sub_0 
   is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end 
   stall_detection_unit_op_code_size6_func_size11_PC_reg_size32_reg_file_size32_DW01_sub_0;

architecture SYN_rpl of 
   stall_detection_unit_op_code_size6_func_size11_PC_reg_size32_reg_file_size32_DW01_sub_0 
   is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal DIFF_31_port, DIFF_30_port, DIFF_29_port, DIFF_28_port, DIFF_27_port,
      DIFF_26_port, DIFF_25_port, DIFF_24_port, DIFF_23_port, DIFF_22_port, 
      DIFF_21_port, DIFF_20_port, DIFF_19_port, DIFF_18_port, DIFF_17_port, 
      DIFF_16_port, DIFF_15_port, DIFF_14_port, DIFF_13_port, DIFF_12_port, 
      DIFF_11_port, DIFF_10_port, DIFF_9_port, DIFF_8_port, DIFF_7_port, 
      DIFF_6_port, DIFF_5_port, DIFF_4_port, DIFF_3_port, DIFF_2_port, 
      carry_31_port, carry_30_port, carry_29_port, carry_28_port, carry_27_port
      , carry_26_port, carry_25_port, carry_24_port, carry_23_port, 
      carry_22_port, carry_21_port, carry_20_port, carry_19_port, carry_18_port
      , carry_17_port, carry_16_port, carry_15_port, carry_14_port, 
      carry_13_port, carry_12_port, carry_11_port, carry_10_port, carry_9_port,
      carry_8_port, carry_7_port, carry_6_port, carry_5_port, carry_4_port, 
      carry_3_port, n1, n2, n3 : std_logic;

begin
   DIFF <= ( DIFF_31_port, DIFF_30_port, DIFF_29_port, DIFF_28_port, 
      DIFF_27_port, DIFF_26_port, DIFF_25_port, DIFF_24_port, DIFF_23_port, 
      DIFF_22_port, DIFF_21_port, DIFF_20_port, DIFF_19_port, DIFF_18_port, 
      DIFF_17_port, DIFF_16_port, DIFF_15_port, DIFF_14_port, DIFF_13_port, 
      DIFF_12_port, DIFF_11_port, DIFF_10_port, DIFF_9_port, DIFF_8_port, 
      DIFF_7_port, DIFF_6_port, DIFF_5_port, DIFF_4_port, DIFF_3_port, 
      DIFF_2_port, A(1), A(0) );
   
   U1 : XNOR2_X1 port map( A => A(10), B => carry_10_port, ZN => DIFF_10_port);
   U2 : XNOR2_X1 port map( A => A(11), B => carry_11_port, ZN => DIFF_11_port);
   U3 : XNOR2_X1 port map( A => A(13), B => carry_13_port, ZN => DIFF_13_port);
   U4 : XNOR2_X1 port map( A => A(15), B => carry_15_port, ZN => DIFF_15_port);
   U5 : XNOR2_X1 port map( A => A(16), B => carry_16_port, ZN => DIFF_16_port);
   U6 : XNOR2_X1 port map( A => A(17), B => carry_17_port, ZN => DIFF_17_port);
   U7 : XNOR2_X1 port map( A => A(18), B => carry_18_port, ZN => DIFF_18_port);
   U8 : XNOR2_X1 port map( A => A(19), B => carry_19_port, ZN => DIFF_19_port);
   U9 : XNOR2_X1 port map( A => A(5), B => carry_5_port, ZN => DIFF_5_port);
   U10 : XNOR2_X1 port map( A => A(8), B => carry_8_port, ZN => DIFF_8_port);
   U11 : XNOR2_X1 port map( A => A(9), B => carry_9_port, ZN => DIFF_9_port);
   U12 : XNOR2_X1 port map( A => A(20), B => carry_20_port, ZN => DIFF_20_port)
                           ;
   U13 : XNOR2_X1 port map( A => A(21), B => carry_21_port, ZN => DIFF_21_port)
                           ;
   U14 : XNOR2_X1 port map( A => A(22), B => carry_22_port, ZN => DIFF_22_port)
                           ;
   U15 : XNOR2_X1 port map( A => A(23), B => carry_23_port, ZN => DIFF_23_port)
                           ;
   U16 : XNOR2_X1 port map( A => A(24), B => carry_24_port, ZN => DIFF_24_port)
                           ;
   U17 : XNOR2_X1 port map( A => A(25), B => carry_25_port, ZN => DIFF_25_port)
                           ;
   U18 : XNOR2_X1 port map( A => A(26), B => carry_26_port, ZN => DIFF_26_port)
                           ;
   U19 : XNOR2_X1 port map( A => A(27), B => carry_27_port, ZN => DIFF_27_port)
                           ;
   U20 : XNOR2_X1 port map( A => A(28), B => carry_28_port, ZN => DIFF_28_port)
                           ;
   U21 : XNOR2_X1 port map( A => A(29), B => carry_29_port, ZN => DIFF_29_port)
                           ;
   U22 : XNOR2_X1 port map( A => A(30), B => carry_30_port, ZN => DIFF_30_port)
                           ;
   U23 : XNOR2_X1 port map( A => A(7), B => carry_7_port, ZN => DIFF_7_port);
   U24 : XNOR2_X1 port map( A => n3, B => A(2), ZN => DIFF_2_port);
   U25 : XNOR2_X1 port map( A => A(3), B => carry_3_port, ZN => DIFF_3_port);
   U26 : XNOR2_X1 port map( A => A(4), B => carry_4_port, ZN => DIFF_4_port);
   U27 : XNOR2_X1 port map( A => A(12), B => carry_12_port, ZN => DIFF_12_port)
                           ;
   U28 : XNOR2_X1 port map( A => A(14), B => carry_14_port, ZN => DIFF_14_port)
                           ;
   U29 : XNOR2_X1 port map( A => A(6), B => carry_6_port, ZN => DIFF_6_port);
   U30 : XNOR2_X1 port map( A => A(31), B => carry_31_port, ZN => DIFF_31_port)
                           ;
   U31 : NAND2_X1 port map( A1 => n1, A2 => n2, ZN => carry_31_port);
   U32 : INV_X1 port map( A => A(30), ZN => n1);
   U33 : INV_X1 port map( A => carry_30_port, ZN => n2);
   U34 : OR2_X1 port map( A1 => n3, A2 => A(2), ZN => carry_3_port);
   U35 : OR2_X1 port map( A1 => A(3), A2 => carry_3_port, ZN => carry_4_port);
   U36 : OR2_X1 port map( A1 => A(7), A2 => carry_7_port, ZN => carry_8_port);
   U37 : OR2_X1 port map( A1 => A(8), A2 => carry_8_port, ZN => carry_9_port);
   U38 : OR2_X1 port map( A1 => A(9), A2 => carry_9_port, ZN => carry_10_port);
   U39 : OR2_X1 port map( A1 => A(10), A2 => carry_10_port, ZN => carry_11_port
                           );
   U40 : OR2_X1 port map( A1 => A(11), A2 => carry_11_port, ZN => carry_12_port
                           );
   U41 : OR2_X1 port map( A1 => A(12), A2 => carry_12_port, ZN => carry_13_port
                           );
   U42 : OR2_X1 port map( A1 => A(13), A2 => carry_13_port, ZN => carry_14_port
                           );
   U43 : OR2_X1 port map( A1 => A(14), A2 => carry_14_port, ZN => carry_15_port
                           );
   U44 : OR2_X1 port map( A1 => A(15), A2 => carry_15_port, ZN => carry_16_port
                           );
   U45 : OR2_X1 port map( A1 => A(16), A2 => carry_16_port, ZN => carry_17_port
                           );
   U46 : OR2_X1 port map( A1 => A(22), A2 => carry_22_port, ZN => carry_23_port
                           );
   U47 : OR2_X1 port map( A1 => A(23), A2 => carry_23_port, ZN => carry_24_port
                           );
   U48 : OR2_X1 port map( A1 => A(24), A2 => carry_24_port, ZN => carry_25_port
                           );
   U49 : OR2_X1 port map( A1 => A(25), A2 => carry_25_port, ZN => carry_26_port
                           );
   U50 : OR2_X1 port map( A1 => A(26), A2 => carry_26_port, ZN => carry_27_port
                           );
   U51 : OR2_X1 port map( A1 => A(27), A2 => carry_27_port, ZN => carry_28_port
                           );
   U52 : OR2_X1 port map( A1 => A(28), A2 => carry_28_port, ZN => carry_29_port
                           );
   U53 : OR2_X1 port map( A1 => A(29), A2 => carry_29_port, ZN => carry_30_port
                           );
   U54 : OR2_X1 port map( A1 => A(4), A2 => carry_4_port, ZN => carry_5_port);
   U55 : OR2_X1 port map( A1 => A(5), A2 => carry_5_port, ZN => carry_6_port);
   U56 : OR2_X1 port map( A1 => A(6), A2 => carry_6_port, ZN => carry_7_port);
   U57 : INV_X1 port map( A => B(2), ZN => n3);
   U58 : OR2_X1 port map( A1 => A(17), A2 => carry_17_port, ZN => carry_18_port
                           );
   U59 : OR2_X1 port map( A1 => A(18), A2 => carry_18_port, ZN => carry_19_port
                           );
   U60 : OR2_X1 port map( A1 => A(19), A2 => carry_19_port, ZN => carry_20_port
                           );
   U61 : OR2_X1 port map( A1 => A(20), A2 => carry_20_port, ZN => carry_21_port
                           );
   U62 : OR2_X1 port map( A1 => A(21), A2 => carry_21_port, ZN => carry_22_port
                           );

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity negate_NBIT32_0_DW01_sub_0 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end negate_NBIT32_0_DW01_sub_0;

architecture SYN_rpl of negate_NBIT32_0_DW01_sub_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal DIFF_2_port, DIFF_3_port, DIFF_4_port, DIFF_1_port, n5, n6, n7, n8, 
      n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
      n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, DIFF_24_port, 
      DIFF_25_port, DIFF_26_port, DIFF_27_port, DIFF_28_port, DIFF_23_port, 
      DIFF_29_port, DIFF_30_port, DIFF_31_port, DIFF_12_port, DIFF_13_port, 
      DIFF_14_port, DIFF_15_port, DIFF_16_port, DIFF_17_port, DIFF_18_port, 
      DIFF_19_port, DIFF_20_port, DIFF_21_port, DIFF_22_port, DIFF_5_port, 
      DIFF_6_port, DIFF_7_port, DIFF_8_port, DIFF_9_port, DIFF_10_port, 
      DIFF_11_port, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
      n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87
      , n88, n89, n90, n91, n92 : std_logic;

begin
   DIFF <= ( DIFF_31_port, DIFF_30_port, DIFF_29_port, DIFF_28_port, 
      DIFF_27_port, DIFF_26_port, DIFF_25_port, DIFF_24_port, DIFF_23_port, 
      DIFF_22_port, DIFF_21_port, DIFF_20_port, DIFF_19_port, DIFF_18_port, 
      DIFF_17_port, DIFF_16_port, DIFF_15_port, DIFF_14_port, DIFF_13_port, 
      DIFF_12_port, DIFF_11_port, DIFF_10_port, DIFF_9_port, DIFF_8_port, 
      DIFF_7_port, DIFF_6_port, DIFF_5_port, DIFF_4_port, DIFF_3_port, 
      DIFF_2_port, DIFF_1_port, B(0) );
   
   U1 : XOR2_X1 port map( A => n63, B => n7, Z => DIFF_2_port);
   U2 : XOR2_X1 port map( A => n64, B => n8, Z => DIFF_3_port);
   U3 : XOR2_X1 port map( A => n65, B => n9, Z => DIFF_4_port);
   U4 : XOR2_X1 port map( A => n62, B => n92, Z => DIFF_1_port);
   U5 : AND2_X1 port map( A1 => n73, A2 => n22, ZN => n5);
   U6 : AND2_X1 port map( A1 => n74, A2 => n5, ZN => n6);
   U7 : AND2_X1 port map( A1 => n62, A2 => n92, ZN => n7);
   U8 : AND2_X1 port map( A1 => n63, A2 => n7, ZN => n8);
   U9 : AND2_X1 port map( A1 => n64, A2 => n8, ZN => n9);
   U10 : AND2_X1 port map( A1 => n65, A2 => n9, ZN => n10);
   U11 : AND2_X1 port map( A1 => n66, A2 => n10, ZN => n11);
   U12 : AND2_X1 port map( A1 => n67, A2 => n11, ZN => n12);
   U13 : AND2_X1 port map( A1 => n68, A2 => n12, ZN => n13);
   U14 : AND2_X1 port map( A1 => n85, A2 => n32, ZN => n14);
   U15 : AND2_X1 port map( A1 => n86, A2 => n14, ZN => n15);
   U16 : AND2_X1 port map( A1 => n87, A2 => n15, ZN => n16);
   U17 : AND2_X1 port map( A1 => n88, A2 => n16, ZN => n17);
   U18 : AND2_X1 port map( A1 => n89, A2 => n17, ZN => n18);
   U19 : AND2_X1 port map( A1 => n69, A2 => n13, ZN => n19);
   U20 : AND2_X1 port map( A1 => n70, A2 => n19, ZN => n20);
   U21 : AND2_X1 port map( A1 => n71, A2 => n20, ZN => n21);
   U22 : AND2_X1 port map( A1 => n72, A2 => n21, ZN => n22);
   U23 : AND2_X1 port map( A1 => n75, A2 => n6, ZN => n23);
   U24 : AND2_X1 port map( A1 => n76, A2 => n23, ZN => n24);
   U25 : AND2_X1 port map( A1 => n77, A2 => n24, ZN => n25);
   U26 : AND2_X1 port map( A1 => n78, A2 => n25, ZN => n26);
   U27 : AND2_X1 port map( A1 => n79, A2 => n26, ZN => n27);
   U28 : AND2_X1 port map( A1 => n80, A2 => n27, ZN => n28);
   U29 : AND2_X1 port map( A1 => n81, A2 => n28, ZN => n29);
   U30 : AND2_X1 port map( A1 => n82, A2 => n29, ZN => n30);
   U31 : AND2_X1 port map( A1 => n83, A2 => n30, ZN => n31);
   U32 : AND2_X1 port map( A1 => n84, A2 => n31, ZN => n32);
   U33 : AND2_X1 port map( A1 => n90, A2 => n18, ZN => n33);
   U34 : NAND2_X1 port map( A1 => n91, A2 => n33, ZN => n61);
   U35 : XOR2_X1 port map( A => n85, B => n32, Z => DIFF_24_port);
   U36 : XOR2_X1 port map( A => n86, B => n14, Z => DIFF_25_port);
   U37 : XOR2_X1 port map( A => n87, B => n15, Z => DIFF_26_port);
   U38 : XOR2_X1 port map( A => n88, B => n16, Z => DIFF_27_port);
   U39 : XOR2_X1 port map( A => n89, B => n17, Z => DIFF_28_port);
   U40 : XOR2_X1 port map( A => n84, B => n31, Z => DIFF_23_port);
   U41 : XOR2_X1 port map( A => n90, B => n18, Z => DIFF_29_port);
   U42 : XOR2_X1 port map( A => n91, B => n33, Z => DIFF_30_port);
   U43 : XOR2_X1 port map( A => B(31), B => n61, Z => DIFF_31_port);
   U44 : XOR2_X1 port map( A => n73, B => n22, Z => DIFF_12_port);
   U45 : XOR2_X1 port map( A => n74, B => n5, Z => DIFF_13_port);
   U46 : XOR2_X1 port map( A => n75, B => n6, Z => DIFF_14_port);
   U47 : XOR2_X1 port map( A => n76, B => n23, Z => DIFF_15_port);
   U48 : XOR2_X1 port map( A => n77, B => n24, Z => DIFF_16_port);
   U49 : XOR2_X1 port map( A => n78, B => n25, Z => DIFF_17_port);
   U50 : XOR2_X1 port map( A => n79, B => n26, Z => DIFF_18_port);
   U51 : XOR2_X1 port map( A => n80, B => n27, Z => DIFF_19_port);
   U52 : XOR2_X1 port map( A => n81, B => n28, Z => DIFF_20_port);
   U53 : XOR2_X1 port map( A => n82, B => n29, Z => DIFF_21_port);
   U54 : XOR2_X1 port map( A => n83, B => n30, Z => DIFF_22_port);
   U55 : XOR2_X1 port map( A => n66, B => n10, Z => DIFF_5_port);
   U56 : XOR2_X1 port map( A => n67, B => n11, Z => DIFF_6_port);
   U57 : XOR2_X1 port map( A => n68, B => n12, Z => DIFF_7_port);
   U58 : XOR2_X1 port map( A => n69, B => n13, Z => DIFF_8_port);
   U59 : XOR2_X1 port map( A => n70, B => n19, Z => DIFF_9_port);
   U60 : XOR2_X1 port map( A => n71, B => n20, Z => DIFF_10_port);
   U61 : XOR2_X1 port map( A => n72, B => n21, Z => DIFF_11_port);
   U62 : INV_X1 port map( A => B(0), ZN => n92);
   U63 : INV_X1 port map( A => B(1), ZN => n62);
   U64 : INV_X1 port map( A => B(2), ZN => n63);
   U65 : INV_X1 port map( A => B(3), ZN => n64);
   U66 : INV_X1 port map( A => B(4), ZN => n65);
   U67 : INV_X1 port map( A => B(5), ZN => n66);
   U68 : INV_X1 port map( A => B(6), ZN => n67);
   U69 : INV_X1 port map( A => B(7), ZN => n68);
   U70 : INV_X1 port map( A => B(8), ZN => n69);
   U71 : INV_X1 port map( A => B(9), ZN => n70);
   U72 : INV_X1 port map( A => B(10), ZN => n71);
   U73 : INV_X1 port map( A => B(11), ZN => n72);
   U74 : INV_X1 port map( A => B(12), ZN => n73);
   U75 : INV_X1 port map( A => B(13), ZN => n74);
   U76 : INV_X1 port map( A => B(14), ZN => n75);
   U77 : INV_X1 port map( A => B(15), ZN => n76);
   U78 : INV_X1 port map( A => B(16), ZN => n77);
   U79 : INV_X1 port map( A => B(17), ZN => n78);
   U80 : INV_X1 port map( A => B(18), ZN => n79);
   U81 : INV_X1 port map( A => B(19), ZN => n80);
   U82 : INV_X1 port map( A => B(20), ZN => n81);
   U83 : INV_X1 port map( A => B(24), ZN => n85);
   U84 : INV_X1 port map( A => B(25), ZN => n86);
   U85 : INV_X1 port map( A => B(26), ZN => n87);
   U86 : INV_X1 port map( A => B(27), ZN => n88);
   U87 : INV_X1 port map( A => B(28), ZN => n89);
   U88 : INV_X1 port map( A => B(21), ZN => n82);
   U89 : INV_X1 port map( A => B(22), ZN => n83);
   U90 : INV_X1 port map( A => B(23), ZN => n84);
   U91 : INV_X1 port map( A => B(29), ZN => n90);
   U92 : INV_X1 port map( A => B(30), ZN => n91);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity negate_NBIT32_7_DW01_sub_0 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end negate_NBIT32_7_DW01_sub_0;

architecture SYN_rpl of negate_NBIT32_7_DW01_sub_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal DIFF_31_port, DIFF_30_port, DIFF_23_port, DIFF_24_port, DIFF_29_port,
      DIFF_25_port, DIFF_26_port, DIFF_27_port, DIFF_28_port, DIFF_12_port, 
      DIFF_13_port, DIFF_14_port, DIFF_15_port, DIFF_16_port, DIFF_17_port, 
      DIFF_18_port, DIFF_19_port, DIFF_20_port, DIFF_21_port, DIFF_22_port, 
      DIFF_9_port, DIFF_10_port, DIFF_11_port, DIFF_8_port, DIFF_5_port, 
      DIFF_6_port, DIFF_7_port, n28, n29, n30, n31, n32, n33, n34, n35, n36, 
      n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51
      , n52, n53, n54, n55, DIFF_2_port, DIFF_3_port, DIFF_4_port, n59, 
      DIFF_1_port, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, 
      n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87
      , n88, n89, n90, n91, n92 : std_logic;

begin
   DIFF <= ( DIFF_31_port, DIFF_30_port, DIFF_29_port, DIFF_28_port, 
      DIFF_27_port, DIFF_26_port, DIFF_25_port, DIFF_24_port, DIFF_23_port, 
      DIFF_22_port, DIFF_21_port, DIFF_20_port, DIFF_19_port, DIFF_18_port, 
      DIFF_17_port, DIFF_16_port, DIFF_15_port, DIFF_14_port, DIFF_13_port, 
      DIFF_12_port, DIFF_11_port, DIFF_10_port, DIFF_9_port, DIFF_8_port, 
      DIFF_7_port, DIFF_6_port, DIFF_5_port, DIFF_4_port, DIFF_3_port, 
      DIFF_2_port, DIFF_1_port, B(0) );
   
   U1 : XOR2_X1 port map( A => B(31), B => n61, Z => DIFF_31_port);
   U2 : XOR2_X1 port map( A => n91, B => n41, Z => DIFF_30_port);
   U3 : XOR2_X1 port map( A => n84, B => n53, Z => DIFF_23_port);
   U4 : XOR2_X1 port map( A => n85, B => n54, Z => DIFF_24_port);
   U5 : XOR2_X1 port map( A => n90, B => n40, Z => DIFF_29_port);
   U6 : XOR2_X1 port map( A => n86, B => n55, Z => DIFF_25_port);
   U7 : XOR2_X1 port map( A => n87, B => n37, Z => DIFF_26_port);
   U8 : XOR2_X1 port map( A => n88, B => n38, Z => DIFF_27_port);
   U9 : XOR2_X1 port map( A => n89, B => n39, Z => DIFF_28_port);
   U10 : XOR2_X1 port map( A => n73, B => n44, Z => DIFF_12_port);
   U11 : XOR2_X1 port map( A => n74, B => n28, Z => DIFF_13_port);
   U12 : XOR2_X1 port map( A => n75, B => n29, Z => DIFF_14_port);
   U13 : XOR2_X1 port map( A => n76, B => n45, Z => DIFF_15_port);
   U14 : XOR2_X1 port map( A => n77, B => n46, Z => DIFF_16_port);
   U15 : XOR2_X1 port map( A => n78, B => n47, Z => DIFF_17_port);
   U16 : XOR2_X1 port map( A => n79, B => n48, Z => DIFF_18_port);
   U17 : XOR2_X1 port map( A => n80, B => n49, Z => DIFF_19_port);
   U18 : XOR2_X1 port map( A => n81, B => n50, Z => DIFF_20_port);
   U19 : XOR2_X1 port map( A => n82, B => n51, Z => DIFF_21_port);
   U20 : XOR2_X1 port map( A => n83, B => n52, Z => DIFF_22_port);
   U21 : XOR2_X1 port map( A => n70, B => n36, Z => DIFF_9_port);
   U22 : XOR2_X1 port map( A => n71, B => n42, Z => DIFF_10_port);
   U23 : XOR2_X1 port map( A => n72, B => n43, Z => DIFF_11_port);
   U24 : XOR2_X1 port map( A => n69, B => n35, Z => DIFF_8_port);
   U25 : XOR2_X1 port map( A => n66, B => n32, Z => DIFF_5_port);
   U26 : XOR2_X1 port map( A => n67, B => n33, Z => DIFF_6_port);
   U27 : XOR2_X1 port map( A => n68, B => n34, Z => DIFF_7_port);
   U28 : AND2_X1 port map( A1 => n73, A2 => n44, ZN => n28);
   U29 : AND2_X1 port map( A1 => n74, A2 => n28, ZN => n29);
   U30 : AND2_X1 port map( A1 => n63, A2 => n59, ZN => n30);
   U31 : AND2_X1 port map( A1 => n64, A2 => n30, ZN => n31);
   U32 : AND2_X1 port map( A1 => n65, A2 => n31, ZN => n32);
   U33 : AND2_X1 port map( A1 => n66, A2 => n32, ZN => n33);
   U34 : AND2_X1 port map( A1 => n67, A2 => n33, ZN => n34);
   U35 : AND2_X1 port map( A1 => n68, A2 => n34, ZN => n35);
   U36 : AND2_X1 port map( A1 => n69, A2 => n35, ZN => n36);
   U37 : AND2_X1 port map( A1 => n86, A2 => n55, ZN => n37);
   U38 : AND2_X1 port map( A1 => n87, A2 => n37, ZN => n38);
   U39 : AND2_X1 port map( A1 => n88, A2 => n38, ZN => n39);
   U40 : AND2_X1 port map( A1 => n89, A2 => n39, ZN => n40);
   U41 : AND2_X1 port map( A1 => n90, A2 => n40, ZN => n41);
   U42 : AND2_X1 port map( A1 => n70, A2 => n36, ZN => n42);
   U43 : AND2_X1 port map( A1 => n71, A2 => n42, ZN => n43);
   U44 : AND2_X1 port map( A1 => n72, A2 => n43, ZN => n44);
   U45 : AND2_X1 port map( A1 => n75, A2 => n29, ZN => n45);
   U46 : AND2_X1 port map( A1 => n76, A2 => n45, ZN => n46);
   U47 : AND2_X1 port map( A1 => n77, A2 => n46, ZN => n47);
   U48 : AND2_X1 port map( A1 => n78, A2 => n47, ZN => n48);
   U49 : AND2_X1 port map( A1 => n79, A2 => n48, ZN => n49);
   U50 : AND2_X1 port map( A1 => n80, A2 => n49, ZN => n50);
   U51 : AND2_X1 port map( A1 => n81, A2 => n50, ZN => n51);
   U52 : AND2_X1 port map( A1 => n82, A2 => n51, ZN => n52);
   U53 : AND2_X1 port map( A1 => n83, A2 => n52, ZN => n53);
   U54 : AND2_X1 port map( A1 => n84, A2 => n53, ZN => n54);
   U55 : AND2_X1 port map( A1 => n85, A2 => n54, ZN => n55);
   U56 : XOR2_X1 port map( A => n63, B => n59, Z => DIFF_2_port);
   U57 : XOR2_X1 port map( A => n64, B => n30, Z => DIFF_3_port);
   U58 : XOR2_X1 port map( A => n65, B => n31, Z => DIFF_4_port);
   U59 : INV_X1 port map( A => B(1), ZN => n92);
   U60 : INV_X1 port map( A => B(2), ZN => n63);
   U61 : INV_X1 port map( A => B(3), ZN => n64);
   U62 : INV_X1 port map( A => B(4), ZN => n65);
   U63 : INV_X1 port map( A => B(5), ZN => n66);
   U64 : INV_X1 port map( A => B(6), ZN => n67);
   U65 : INV_X1 port map( A => B(7), ZN => n68);
   U66 : INV_X1 port map( A => B(8), ZN => n69);
   U67 : INV_X1 port map( A => B(9), ZN => n70);
   U68 : NAND2_X1 port map( A1 => n91, A2 => n41, ZN => n61);
   U69 : AND2_X1 port map( A1 => n92, A2 => n62, ZN => n59);
   U70 : INV_X1 port map( A => B(10), ZN => n71);
   U71 : INV_X1 port map( A => B(11), ZN => n72);
   U72 : INV_X1 port map( A => B(12), ZN => n73);
   U73 : INV_X1 port map( A => B(13), ZN => n74);
   U74 : INV_X1 port map( A => B(14), ZN => n75);
   U75 : INV_X1 port map( A => B(15), ZN => n76);
   U76 : INV_X1 port map( A => B(16), ZN => n77);
   U77 : INV_X1 port map( A => B(17), ZN => n78);
   U78 : INV_X1 port map( A => B(18), ZN => n79);
   U79 : INV_X1 port map( A => B(19), ZN => n80);
   U80 : INV_X1 port map( A => B(25), ZN => n86);
   U81 : INV_X1 port map( A => B(26), ZN => n87);
   U82 : INV_X1 port map( A => B(27), ZN => n88);
   U83 : INV_X1 port map( A => B(28), ZN => n89);
   U84 : INV_X1 port map( A => B(29), ZN => n90);
   U85 : INV_X1 port map( A => B(20), ZN => n81);
   U86 : INV_X1 port map( A => B(21), ZN => n82);
   U87 : INV_X1 port map( A => B(22), ZN => n83);
   U88 : INV_X1 port map( A => B(23), ZN => n84);
   U89 : INV_X1 port map( A => B(24), ZN => n85);
   U90 : INV_X1 port map( A => B(30), ZN => n91);
   U91 : XOR2_X1 port map( A => n92, B => n62, Z => DIFF_1_port);
   U92 : INV_X1 port map( A => B(0), ZN => n62);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity negate_NBIT32_6_DW01_sub_0 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end negate_NBIT32_6_DW01_sub_0;

architecture SYN_rpl of negate_NBIT32_6_DW01_sub_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal DIFF_4_port, DIFF_5_port, DIFF_3_port, n4, n5, n6, n7, n8, n9, n10, 
      n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25
      , n26, n27, n28, n29, n30, n31, DIFF_26_port, DIFF_27_port, DIFF_28_port,
      DIFF_29_port, DIFF_30_port, DIFF_24_port, DIFF_25_port, DIFF_13_port, 
      DIFF_14_port, DIFF_15_port, DIFF_16_port, DIFF_17_port, DIFF_18_port, 
      DIFF_19_port, DIFF_20_port, DIFF_21_port, DIFF_22_port, DIFF_23_port, 
      DIFF_6_port, DIFF_7_port, DIFF_8_port, DIFF_9_port, DIFF_10_port, 
      DIFF_11_port, DIFF_12_port, DIFF_2_port, DIFF_31_port, n59, DIFF_1_port, 
      n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75
      , n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, 
      n90, n91, n92 : std_logic;

begin
   DIFF <= ( DIFF_31_port, DIFF_30_port, DIFF_29_port, DIFF_28_port, 
      DIFF_27_port, DIFF_26_port, DIFF_25_port, DIFF_24_port, DIFF_23_port, 
      DIFF_22_port, DIFF_21_port, DIFF_20_port, DIFF_19_port, DIFF_18_port, 
      DIFF_17_port, DIFF_16_port, DIFF_15_port, DIFF_14_port, DIFF_13_port, 
      DIFF_12_port, DIFF_11_port, DIFF_10_port, DIFF_9_port, DIFF_8_port, 
      DIFF_7_port, DIFF_6_port, DIFF_5_port, DIFF_4_port, DIFF_3_port, 
      DIFF_2_port, DIFF_1_port, B(0) );
   
   U1 : XOR2_X1 port map( A => n65, B => n8, Z => DIFF_4_port);
   U2 : XOR2_X1 port map( A => n66, B => n9, Z => DIFF_5_port);
   U3 : XOR2_X1 port map( A => n64, B => n7, Z => DIFF_3_port);
   U4 : NAND2_X1 port map( A1 => n91, A2 => n18, ZN => n61);
   U5 : AND2_X1 port map( A1 => n73, A2 => n20, ZN => n4);
   U6 : AND2_X1 port map( A1 => n74, A2 => n4, ZN => n5);
   U7 : AND2_X1 port map( A1 => n75, A2 => n5, ZN => n6);
   U8 : AND2_X1 port map( A1 => n92, A2 => n59, ZN => n7);
   U9 : AND2_X1 port map( A1 => n64, A2 => n7, ZN => n8);
   U10 : AND2_X1 port map( A1 => n65, A2 => n8, ZN => n9);
   U11 : AND2_X1 port map( A1 => n66, A2 => n9, ZN => n10);
   U12 : AND2_X1 port map( A1 => n67, A2 => n10, ZN => n11);
   U13 : AND2_X1 port map( A1 => n68, A2 => n11, ZN => n12);
   U14 : AND2_X1 port map( A1 => n69, A2 => n12, ZN => n13);
   U15 : AND2_X1 port map( A1 => n70, A2 => n13, ZN => n14);
   U16 : AND2_X1 port map( A1 => n87, A2 => n31, ZN => n15);
   U17 : AND2_X1 port map( A1 => n88, A2 => n15, ZN => n16);
   U18 : AND2_X1 port map( A1 => n89, A2 => n16, ZN => n17);
   U19 : AND2_X1 port map( A1 => n90, A2 => n17, ZN => n18);
   U20 : AND2_X1 port map( A1 => n71, A2 => n14, ZN => n19);
   U21 : AND2_X1 port map( A1 => n72, A2 => n19, ZN => n20);
   U22 : AND2_X1 port map( A1 => n76, A2 => n6, ZN => n21);
   U23 : AND2_X1 port map( A1 => n77, A2 => n21, ZN => n22);
   U24 : AND2_X1 port map( A1 => n78, A2 => n22, ZN => n23);
   U25 : AND2_X1 port map( A1 => n79, A2 => n23, ZN => n24);
   U26 : AND2_X1 port map( A1 => n80, A2 => n24, ZN => n25);
   U27 : AND2_X1 port map( A1 => n81, A2 => n25, ZN => n26);
   U28 : AND2_X1 port map( A1 => n82, A2 => n26, ZN => n27);
   U29 : AND2_X1 port map( A1 => n83, A2 => n27, ZN => n28);
   U30 : AND2_X1 port map( A1 => n84, A2 => n28, ZN => n29);
   U31 : AND2_X1 port map( A1 => n85, A2 => n29, ZN => n30);
   U32 : AND2_X1 port map( A1 => n86, A2 => n30, ZN => n31);
   U33 : XOR2_X1 port map( A => n87, B => n31, Z => DIFF_26_port);
   U34 : XOR2_X1 port map( A => n88, B => n15, Z => DIFF_27_port);
   U35 : XOR2_X1 port map( A => n89, B => n16, Z => DIFF_28_port);
   U36 : XOR2_X1 port map( A => n90, B => n17, Z => DIFF_29_port);
   U37 : XOR2_X1 port map( A => n91, B => n18, Z => DIFF_30_port);
   U38 : XOR2_X1 port map( A => n85, B => n29, Z => DIFF_24_port);
   U39 : XOR2_X1 port map( A => n86, B => n30, Z => DIFF_25_port);
   U40 : XOR2_X1 port map( A => n74, B => n4, Z => DIFF_13_port);
   U41 : XOR2_X1 port map( A => n75, B => n5, Z => DIFF_14_port);
   U42 : XOR2_X1 port map( A => n76, B => n6, Z => DIFF_15_port);
   U43 : XOR2_X1 port map( A => n77, B => n21, Z => DIFF_16_port);
   U44 : XOR2_X1 port map( A => n78, B => n22, Z => DIFF_17_port);
   U45 : XOR2_X1 port map( A => n79, B => n23, Z => DIFF_18_port);
   U46 : XOR2_X1 port map( A => n80, B => n24, Z => DIFF_19_port);
   U47 : XOR2_X1 port map( A => n81, B => n25, Z => DIFF_20_port);
   U48 : XOR2_X1 port map( A => n82, B => n26, Z => DIFF_21_port);
   U49 : XOR2_X1 port map( A => n83, B => n27, Z => DIFF_22_port);
   U50 : XOR2_X1 port map( A => n84, B => n28, Z => DIFF_23_port);
   U51 : XOR2_X1 port map( A => n67, B => n10, Z => DIFF_6_port);
   U52 : XOR2_X1 port map( A => n68, B => n11, Z => DIFF_7_port);
   U53 : XOR2_X1 port map( A => n69, B => n12, Z => DIFF_8_port);
   U54 : XOR2_X1 port map( A => n70, B => n13, Z => DIFF_9_port);
   U55 : XOR2_X1 port map( A => n71, B => n14, Z => DIFF_10_port);
   U56 : XOR2_X1 port map( A => n72, B => n19, Z => DIFF_11_port);
   U57 : XOR2_X1 port map( A => n73, B => n20, Z => DIFF_12_port);
   U58 : XOR2_X1 port map( A => n92, B => n59, Z => DIFF_2_port);
   U59 : INV_X1 port map( A => B(2), ZN => n92);
   U60 : INV_X1 port map( A => B(3), ZN => n64);
   U61 : INV_X1 port map( A => B(4), ZN => n65);
   U62 : INV_X1 port map( A => B(5), ZN => n66);
   U63 : INV_X1 port map( A => B(6), ZN => n67);
   U64 : INV_X1 port map( A => B(7), ZN => n68);
   U65 : INV_X1 port map( A => B(8), ZN => n69);
   U66 : INV_X1 port map( A => B(9), ZN => n70);
   U67 : XOR2_X1 port map( A => B(31), B => n61, Z => DIFF_31_port);
   U68 : INV_X1 port map( A => B(10), ZN => n71);
   U69 : INV_X1 port map( A => B(11), ZN => n72);
   U70 : INV_X1 port map( A => B(12), ZN => n73);
   U71 : INV_X1 port map( A => B(13), ZN => n74);
   U72 : INV_X1 port map( A => B(14), ZN => n75);
   U73 : INV_X1 port map( A => B(15), ZN => n76);
   U74 : INV_X1 port map( A => B(16), ZN => n77);
   U75 : INV_X1 port map( A => B(17), ZN => n78);
   U76 : INV_X1 port map( A => B(18), ZN => n79);
   U77 : INV_X1 port map( A => B(19), ZN => n80);
   U78 : INV_X1 port map( A => B(20), ZN => n81);
   U79 : INV_X1 port map( A => B(26), ZN => n87);
   U80 : INV_X1 port map( A => B(27), ZN => n88);
   U81 : INV_X1 port map( A => B(28), ZN => n89);
   U82 : INV_X1 port map( A => B(29), ZN => n90);
   U83 : INV_X1 port map( A => B(30), ZN => n91);
   U84 : INV_X1 port map( A => B(21), ZN => n82);
   U85 : INV_X1 port map( A => B(22), ZN => n83);
   U86 : INV_X1 port map( A => B(23), ZN => n84);
   U87 : INV_X1 port map( A => B(24), ZN => n85);
   U88 : INV_X1 port map( A => B(25), ZN => n86);
   U89 : AND2_X1 port map( A1 => n63, A2 => n62, ZN => n59);
   U90 : XOR2_X1 port map( A => n63, B => n62, Z => DIFF_1_port);
   U91 : INV_X1 port map( A => B(0), ZN => n62);
   U92 : INV_X1 port map( A => B(1), ZN => n63);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity negate_NBIT32_5_DW01_sub_0 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end negate_NBIT32_5_DW01_sub_0;

architecture SYN_rpl of negate_NBIT32_5_DW01_sub_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal DIFF_31_port, DIFF_25_port, DIFF_26_port, DIFF_30_port, DIFF_27_port,
      DIFF_28_port, DIFF_29_port, DIFF_24_port, DIFF_13_port, DIFF_14_port, 
      DIFF_15_port, DIFF_16_port, DIFF_17_port, DIFF_18_port, DIFF_19_port, 
      DIFF_20_port, DIFF_21_port, DIFF_22_port, DIFF_23_port, DIFF_11_port, 
      DIFF_12_port, DIFF_10_port, DIFF_6_port, DIFF_7_port, DIFF_8_port, 
      DIFF_9_port, DIFF_2_port, DIFF_1_port, n29, n30, n31, n32, n33, n34, n35,
      n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50
      , n51, n52, n53, n54, n55, DIFF_4_port, DIFF_5_port, DIFF_3_port, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92 : std_logic;

begin
   DIFF <= ( DIFF_31_port, DIFF_30_port, DIFF_29_port, DIFF_28_port, 
      DIFF_27_port, DIFF_26_port, DIFF_25_port, DIFF_24_port, DIFF_23_port, 
      DIFF_22_port, DIFF_21_port, DIFF_20_port, DIFF_19_port, DIFF_18_port, 
      DIFF_17_port, DIFF_16_port, DIFF_15_port, DIFF_14_port, DIFF_13_port, 
      DIFF_12_port, DIFF_11_port, DIFF_10_port, DIFF_9_port, DIFF_8_port, 
      DIFF_7_port, DIFF_6_port, DIFF_5_port, DIFF_4_port, DIFF_3_port, 
      DIFF_2_port, DIFF_1_port, B(0) );
   
   U1 : XOR2_X1 port map( A => B(31), B => n61, Z => DIFF_31_port);
   U2 : XOR2_X1 port map( A => n86, B => n53, Z => DIFF_25_port);
   U3 : XOR2_X1 port map( A => n87, B => n54, Z => DIFF_26_port);
   U4 : XOR2_X1 port map( A => n91, B => n43, Z => DIFF_30_port);
   U5 : XOR2_X1 port map( A => n88, B => n55, Z => DIFF_27_port);
   U6 : XOR2_X1 port map( A => n89, B => n41, Z => DIFF_28_port);
   U7 : XOR2_X1 port map( A => n90, B => n42, Z => DIFF_29_port);
   U8 : XOR2_X1 port map( A => n85, B => n52, Z => DIFF_24_port);
   U9 : XOR2_X1 port map( A => n74, B => n29, Z => DIFF_13_port);
   U10 : XOR2_X1 port map( A => n75, B => n30, Z => DIFF_14_port);
   U11 : XOR2_X1 port map( A => n76, B => n31, Z => DIFF_15_port);
   U12 : XOR2_X1 port map( A => n77, B => n32, Z => DIFF_16_port);
   U13 : XOR2_X1 port map( A => n78, B => n45, Z => DIFF_17_port);
   U14 : XOR2_X1 port map( A => n79, B => n46, Z => DIFF_18_port);
   U15 : XOR2_X1 port map( A => n80, B => n47, Z => DIFF_19_port);
   U16 : XOR2_X1 port map( A => n81, B => n48, Z => DIFF_20_port);
   U17 : XOR2_X1 port map( A => n82, B => n49, Z => DIFF_21_port);
   U18 : XOR2_X1 port map( A => n83, B => n50, Z => DIFF_22_port);
   U19 : XOR2_X1 port map( A => n84, B => n51, Z => DIFF_23_port);
   U20 : XOR2_X1 port map( A => n72, B => n40, Z => DIFF_11_port);
   U21 : XOR2_X1 port map( A => n73, B => n44, Z => DIFF_12_port);
   U22 : XOR2_X1 port map( A => n71, B => n39, Z => DIFF_10_port);
   U23 : XOR2_X1 port map( A => n67, B => n35, Z => DIFF_6_port);
   U24 : XOR2_X1 port map( A => n68, B => n36, Z => DIFF_7_port);
   U25 : XOR2_X1 port map( A => n69, B => n37, Z => DIFF_8_port);
   U26 : XOR2_X1 port map( A => n70, B => n38, Z => DIFF_9_port);
   U27 : XOR2_X1 port map( A => n64, B => n60, Z => DIFF_2_port);
   U28 : XOR2_X1 port map( A => n63, B => n62, Z => DIFF_1_port);
   U29 : AND2_X1 port map( A1 => n73, A2 => n44, ZN => n29);
   U30 : AND2_X1 port map( A1 => n74, A2 => n29, ZN => n30);
   U31 : AND2_X1 port map( A1 => n75, A2 => n30, ZN => n31);
   U32 : AND2_X1 port map( A1 => n76, A2 => n31, ZN => n32);
   U33 : AND2_X1 port map( A1 => n92, A2 => n59, ZN => n33);
   U34 : AND2_X1 port map( A1 => n65, A2 => n33, ZN => n34);
   U35 : AND2_X1 port map( A1 => n66, A2 => n34, ZN => n35);
   U36 : AND2_X1 port map( A1 => n67, A2 => n35, ZN => n36);
   U37 : AND2_X1 port map( A1 => n68, A2 => n36, ZN => n37);
   U38 : AND2_X1 port map( A1 => n69, A2 => n37, ZN => n38);
   U39 : AND2_X1 port map( A1 => n70, A2 => n38, ZN => n39);
   U40 : AND2_X1 port map( A1 => n71, A2 => n39, ZN => n40);
   U41 : AND2_X1 port map( A1 => n88, A2 => n55, ZN => n41);
   U42 : AND2_X1 port map( A1 => n89, A2 => n41, ZN => n42);
   U43 : AND2_X1 port map( A1 => n90, A2 => n42, ZN => n43);
   U44 : AND2_X1 port map( A1 => n72, A2 => n40, ZN => n44);
   U45 : AND2_X1 port map( A1 => n77, A2 => n32, ZN => n45);
   U46 : AND2_X1 port map( A1 => n78, A2 => n45, ZN => n46);
   U47 : AND2_X1 port map( A1 => n79, A2 => n46, ZN => n47);
   U48 : AND2_X1 port map( A1 => n80, A2 => n47, ZN => n48);
   U49 : AND2_X1 port map( A1 => n81, A2 => n48, ZN => n49);
   U50 : AND2_X1 port map( A1 => n82, A2 => n49, ZN => n50);
   U51 : AND2_X1 port map( A1 => n83, A2 => n50, ZN => n51);
   U52 : AND2_X1 port map( A1 => n84, A2 => n51, ZN => n52);
   U53 : AND2_X1 port map( A1 => n85, A2 => n52, ZN => n53);
   U54 : AND2_X1 port map( A1 => n86, A2 => n53, ZN => n54);
   U55 : AND2_X1 port map( A1 => n87, A2 => n54, ZN => n55);
   U56 : XOR2_X1 port map( A => n65, B => n33, Z => DIFF_4_port);
   U57 : XOR2_X1 port map( A => n66, B => n34, Z => DIFF_5_port);
   U58 : XOR2_X1 port map( A => n92, B => n59, Z => DIFF_3_port);
   U59 : INV_X1 port map( A => B(3), ZN => n92);
   U60 : INV_X1 port map( A => B(4), ZN => n65);
   U61 : INV_X1 port map( A => B(5), ZN => n66);
   U62 : INV_X1 port map( A => B(6), ZN => n67);
   U63 : INV_X1 port map( A => B(7), ZN => n68);
   U64 : INV_X1 port map( A => B(8), ZN => n69);
   U65 : INV_X1 port map( A => B(9), ZN => n70);
   U66 : NAND2_X1 port map( A1 => n91, A2 => n43, ZN => n61);
   U67 : INV_X1 port map( A => B(10), ZN => n71);
   U68 : INV_X1 port map( A => B(11), ZN => n72);
   U69 : INV_X1 port map( A => B(12), ZN => n73);
   U70 : INV_X1 port map( A => B(13), ZN => n74);
   U71 : INV_X1 port map( A => B(14), ZN => n75);
   U72 : INV_X1 port map( A => B(15), ZN => n76);
   U73 : INV_X1 port map( A => B(16), ZN => n77);
   U74 : INV_X1 port map( A => B(17), ZN => n78);
   U75 : INV_X1 port map( A => B(18), ZN => n79);
   U76 : INV_X1 port map( A => B(19), ZN => n80);
   U77 : INV_X1 port map( A => B(27), ZN => n88);
   U78 : INV_X1 port map( A => B(28), ZN => n89);
   U79 : INV_X1 port map( A => B(29), ZN => n90);
   U80 : INV_X1 port map( A => B(30), ZN => n91);
   U81 : INV_X1 port map( A => B(20), ZN => n81);
   U82 : INV_X1 port map( A => B(21), ZN => n82);
   U83 : INV_X1 port map( A => B(22), ZN => n83);
   U84 : INV_X1 port map( A => B(23), ZN => n84);
   U85 : INV_X1 port map( A => B(24), ZN => n85);
   U86 : INV_X1 port map( A => B(25), ZN => n86);
   U87 : INV_X1 port map( A => B(26), ZN => n87);
   U88 : AND2_X1 port map( A1 => n64, A2 => n60, ZN => n59);
   U89 : AND2_X1 port map( A1 => n63, A2 => n62, ZN => n60);
   U90 : INV_X1 port map( A => B(0), ZN => n62);
   U91 : INV_X1 port map( A => B(1), ZN => n63);
   U92 : INV_X1 port map( A => B(2), ZN => n64);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity negate_NBIT32_4_DW01_sub_0 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end negate_NBIT32_4_DW01_sub_0;

architecture SYN_rpl of negate_NBIT32_4_DW01_sub_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal DIFF_6_port, DIFF_5_port, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, 
      n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27
      , n28, DIFF_30_port, DIFF_29_port, DIFF_28_port, DIFF_27_port, 
      DIFF_26_port, DIFF_25_port, DIFF_24_port, DIFF_23_port, DIFF_22_port, 
      DIFF_21_port, DIFF_20_port, DIFF_19_port, DIFF_18_port, DIFF_17_port, 
      DIFF_16_port, DIFF_15_port, DIFF_14_port, DIFF_13_port, DIFF_12_port, 
      DIFF_11_port, DIFF_10_port, DIFF_9_port, DIFF_8_port, DIFF_7_port, 
      DIFF_4_port, n54, n55, n56, DIFF_3_port, DIFF_2_port, DIFF_1_port, 
      DIFF_31_port, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
      n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87
      , n88, n89, n90, n91, n92 : std_logic;

begin
   DIFF <= ( DIFF_31_port, DIFF_30_port, DIFF_29_port, DIFF_28_port, 
      DIFF_27_port, DIFF_26_port, DIFF_25_port, DIFF_24_port, DIFF_23_port, 
      DIFF_22_port, DIFF_21_port, DIFF_20_port, DIFF_19_port, DIFF_18_port, 
      DIFF_17_port, DIFF_16_port, DIFF_15_port, DIFF_14_port, DIFF_13_port, 
      DIFF_12_port, DIFF_11_port, DIFF_10_port, DIFF_9_port, DIFF_8_port, 
      DIFF_7_port, DIFF_6_port, DIFF_5_port, DIFF_4_port, DIFF_3_port, 
      DIFF_2_port, DIFF_1_port, B(0) );
   
   U1 : XOR2_X1 port map( A => n87, B => n4, Z => DIFF_6_port);
   U2 : XOR2_X1 port map( A => n88, B => n3, Z => DIFF_5_port);
   U3 : AND2_X1 port map( A1 => n89, A2 => n54, ZN => n3);
   U4 : AND2_X1 port map( A1 => n88, A2 => n3, ZN => n4);
   U5 : AND2_X1 port map( A1 => n87, A2 => n4, ZN => n5);
   U6 : AND2_X1 port map( A1 => n85, A2 => n28, ZN => n6);
   U7 : AND2_X1 port map( A1 => n84, A2 => n6, ZN => n7);
   U8 : AND2_X1 port map( A1 => n83, A2 => n7, ZN => n8);
   U9 : AND2_X1 port map( A1 => n82, A2 => n8, ZN => n9);
   U10 : AND2_X1 port map( A1 => n81, A2 => n9, ZN => n10);
   U11 : AND2_X1 port map( A1 => n80, A2 => n10, ZN => n11);
   U12 : AND2_X1 port map( A1 => n79, A2 => n11, ZN => n12);
   U13 : AND2_X1 port map( A1 => n78, A2 => n12, ZN => n13);
   U14 : AND2_X1 port map( A1 => n77, A2 => n13, ZN => n14);
   U15 : AND2_X1 port map( A1 => n76, A2 => n14, ZN => n15);
   U16 : AND2_X1 port map( A1 => n75, A2 => n15, ZN => n16);
   U17 : AND2_X1 port map( A1 => n74, A2 => n16, ZN => n17);
   U18 : AND2_X1 port map( A1 => n73, A2 => n17, ZN => n18);
   U19 : AND2_X1 port map( A1 => n72, A2 => n18, ZN => n19);
   U20 : AND2_X1 port map( A1 => n71, A2 => n19, ZN => n20);
   U21 : AND2_X1 port map( A1 => n70, A2 => n20, ZN => n21);
   U22 : AND2_X1 port map( A1 => n69, A2 => n21, ZN => n22);
   U23 : AND2_X1 port map( A1 => n68, A2 => n22, ZN => n23);
   U24 : AND2_X1 port map( A1 => n67, A2 => n23, ZN => n24);
   U25 : AND2_X1 port map( A1 => n66, A2 => n24, ZN => n25);
   U26 : AND2_X1 port map( A1 => n65, A2 => n25, ZN => n26);
   U27 : AND2_X1 port map( A1 => n64, A2 => n26, ZN => n27);
   U28 : AND2_X1 port map( A1 => n86, A2 => n5, ZN => n28);
   U29 : NAND2_X1 port map( A1 => n63, A2 => n27, ZN => n61);
   U30 : XOR2_X1 port map( A => n63, B => n27, Z => DIFF_30_port);
   U31 : XOR2_X1 port map( A => n64, B => n26, Z => DIFF_29_port);
   U32 : XOR2_X1 port map( A => n65, B => n25, Z => DIFF_28_port);
   U33 : XOR2_X1 port map( A => n66, B => n24, Z => DIFF_27_port);
   U34 : XOR2_X1 port map( A => n67, B => n23, Z => DIFF_26_port);
   U35 : XOR2_X1 port map( A => n68, B => n22, Z => DIFF_25_port);
   U36 : XOR2_X1 port map( A => n69, B => n21, Z => DIFF_24_port);
   U37 : XOR2_X1 port map( A => n70, B => n20, Z => DIFF_23_port);
   U38 : XOR2_X1 port map( A => n71, B => n19, Z => DIFF_22_port);
   U39 : XOR2_X1 port map( A => n72, B => n18, Z => DIFF_21_port);
   U40 : XOR2_X1 port map( A => n73, B => n17, Z => DIFF_20_port);
   U41 : XOR2_X1 port map( A => n74, B => n16, Z => DIFF_19_port);
   U42 : XOR2_X1 port map( A => n75, B => n15, Z => DIFF_18_port);
   U43 : XOR2_X1 port map( A => n76, B => n14, Z => DIFF_17_port);
   U44 : XOR2_X1 port map( A => n77, B => n13, Z => DIFF_16_port);
   U45 : XOR2_X1 port map( A => n78, B => n12, Z => DIFF_15_port);
   U46 : XOR2_X1 port map( A => n79, B => n11, Z => DIFF_14_port);
   U47 : XOR2_X1 port map( A => n80, B => n10, Z => DIFF_13_port);
   U48 : XOR2_X1 port map( A => n81, B => n9, Z => DIFF_12_port);
   U49 : XOR2_X1 port map( A => n82, B => n8, Z => DIFF_11_port);
   U50 : XOR2_X1 port map( A => n83, B => n7, Z => DIFF_10_port);
   U51 : XOR2_X1 port map( A => n84, B => n6, Z => DIFF_9_port);
   U52 : XOR2_X1 port map( A => n85, B => n28, Z => DIFF_8_port);
   U53 : XOR2_X1 port map( A => n86, B => n5, Z => DIFF_7_port);
   U54 : XOR2_X1 port map( A => n89, B => n54, Z => DIFF_4_port);
   U55 : AND2_X1 port map( A1 => n90, A2 => n55, ZN => n54);
   U56 : AND2_X1 port map( A1 => n91, A2 => n56, ZN => n55);
   U57 : AND2_X1 port map( A1 => n92, A2 => n62, ZN => n56);
   U58 : XOR2_X1 port map( A => n90, B => n55, Z => DIFF_3_port);
   U59 : XOR2_X1 port map( A => n91, B => n56, Z => DIFF_2_port);
   U60 : XOR2_X1 port map( A => n92, B => n62, Z => DIFF_1_port);
   U61 : INV_X1 port map( A => B(4), ZN => n89);
   U62 : INV_X1 port map( A => B(5), ZN => n88);
   U63 : INV_X1 port map( A => B(6), ZN => n87);
   U64 : INV_X1 port map( A => B(7), ZN => n86);
   U65 : INV_X1 port map( A => B(8), ZN => n85);
   U66 : INV_X1 port map( A => B(9), ZN => n84);
   U67 : INV_X1 port map( A => B(10), ZN => n83);
   U68 : INV_X1 port map( A => B(11), ZN => n82);
   U69 : INV_X1 port map( A => B(12), ZN => n81);
   U70 : INV_X1 port map( A => B(13), ZN => n80);
   U71 : XOR2_X1 port map( A => B(31), B => n61, Z => DIFF_31_port);
   U72 : INV_X1 port map( A => B(14), ZN => n79);
   U73 : INV_X1 port map( A => B(15), ZN => n78);
   U74 : INV_X1 port map( A => B(16), ZN => n77);
   U75 : INV_X1 port map( A => B(17), ZN => n76);
   U76 : INV_X1 port map( A => B(18), ZN => n75);
   U77 : INV_X1 port map( A => B(19), ZN => n74);
   U78 : INV_X1 port map( A => B(20), ZN => n73);
   U79 : INV_X1 port map( A => B(21), ZN => n72);
   U80 : INV_X1 port map( A => B(22), ZN => n71);
   U81 : INV_X1 port map( A => B(23), ZN => n70);
   U82 : INV_X1 port map( A => B(24), ZN => n69);
   U83 : INV_X1 port map( A => B(25), ZN => n68);
   U84 : INV_X1 port map( A => B(26), ZN => n67);
   U85 : INV_X1 port map( A => B(27), ZN => n66);
   U86 : INV_X1 port map( A => B(28), ZN => n65);
   U87 : INV_X1 port map( A => B(29), ZN => n64);
   U88 : INV_X1 port map( A => B(30), ZN => n63);
   U89 : INV_X1 port map( A => B(0), ZN => n62);
   U90 : INV_X1 port map( A => B(1), ZN => n92);
   U91 : INV_X1 port map( A => B(2), ZN => n91);
   U92 : INV_X1 port map( A => B(3), ZN => n90);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity negate_NBIT32_3_DW01_sub_0 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end negate_NBIT32_3_DW01_sub_0;

architecture SYN_rpl of negate_NBIT32_3_DW01_sub_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal DIFF_31_port, DIFF_30_port, DIFF_29_port, DIFF_28_port, DIFF_27_port,
      DIFF_26_port, DIFF_25_port, DIFF_24_port, DIFF_23_port, DIFF_22_port, 
      DIFF_21_port, DIFF_20_port, DIFF_19_port, DIFF_18_port, DIFF_17_port, 
      DIFF_16_port, DIFF_15_port, DIFF_14_port, DIFF_13_port, DIFF_12_port, 
      DIFF_11_port, DIFF_9_port, DIFF_8_port, DIFF_10_port, DIFF_7_port, 
      DIFF_4_port, DIFF_3_port, DIFF_2_port, DIFF_1_port, n30, n31, n32, n33, 
      n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48
      , n49, n50, n51, n52, n53, n54, DIFF_6_port, DIFF_5_port, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92 : std_logic;

begin
   DIFF <= ( DIFF_31_port, DIFF_30_port, DIFF_29_port, DIFF_28_port, 
      DIFF_27_port, DIFF_26_port, DIFF_25_port, DIFF_24_port, DIFF_23_port, 
      DIFF_22_port, DIFF_21_port, DIFF_20_port, DIFF_19_port, DIFF_18_port, 
      DIFF_17_port, DIFF_16_port, DIFF_15_port, DIFF_14_port, DIFF_13_port, 
      DIFF_12_port, DIFF_11_port, DIFF_10_port, DIFF_9_port, DIFF_8_port, 
      DIFF_7_port, DIFF_6_port, DIFF_5_port, DIFF_4_port, DIFF_3_port, 
      DIFF_2_port, DIFF_1_port, B(0) );
   
   U1 : XOR2_X1 port map( A => B(31), B => n61, Z => DIFF_31_port);
   U2 : XOR2_X1 port map( A => n64, B => n54, Z => DIFF_30_port);
   U3 : XOR2_X1 port map( A => n65, B => n53, Z => DIFF_29_port);
   U4 : XOR2_X1 port map( A => n66, B => n52, Z => DIFF_28_port);
   U5 : XOR2_X1 port map( A => n67, B => n51, Z => DIFF_27_port);
   U6 : XOR2_X1 port map( A => n68, B => n50, Z => DIFF_26_port);
   U7 : XOR2_X1 port map( A => n69, B => n49, Z => DIFF_25_port);
   U8 : XOR2_X1 port map( A => n70, B => n48, Z => DIFF_24_port);
   U9 : XOR2_X1 port map( A => n71, B => n47, Z => DIFF_23_port);
   U10 : XOR2_X1 port map( A => n72, B => n46, Z => DIFF_22_port);
   U11 : XOR2_X1 port map( A => n73, B => n45, Z => DIFF_21_port);
   U12 : XOR2_X1 port map( A => n74, B => n44, Z => DIFF_20_port);
   U13 : XOR2_X1 port map( A => n75, B => n43, Z => DIFF_19_port);
   U14 : XOR2_X1 port map( A => n76, B => n42, Z => DIFF_18_port);
   U15 : XOR2_X1 port map( A => n77, B => n41, Z => DIFF_17_port);
   U16 : XOR2_X1 port map( A => n78, B => n40, Z => DIFF_16_port);
   U17 : XOR2_X1 port map( A => n79, B => n39, Z => DIFF_15_port);
   U18 : XOR2_X1 port map( A => n80, B => n38, Z => DIFF_14_port);
   U19 : XOR2_X1 port map( A => n81, B => n37, Z => DIFF_13_port);
   U20 : XOR2_X1 port map( A => n82, B => n36, Z => DIFF_12_port);
   U21 : XOR2_X1 port map( A => n83, B => n35, Z => DIFF_11_port);
   U22 : XOR2_X1 port map( A => n85, B => n33, Z => DIFF_9_port);
   U23 : XOR2_X1 port map( A => n86, B => n32, Z => DIFF_8_port);
   U24 : XOR2_X1 port map( A => n84, B => n34, Z => DIFF_10_port);
   U25 : XOR2_X1 port map( A => n87, B => n31, Z => DIFF_7_port);
   U26 : XOR2_X1 port map( A => n90, B => n57, Z => DIFF_4_port);
   U27 : XOR2_X1 port map( A => n91, B => n59, Z => DIFF_3_port);
   U28 : XOR2_X1 port map( A => n92, B => n60, Z => DIFF_2_port);
   U29 : XOR2_X1 port map( A => n63, B => n62, Z => DIFF_1_port);
   U30 : AND2_X1 port map( A1 => n89, A2 => n58, ZN => n30);
   U31 : AND2_X1 port map( A1 => n88, A2 => n30, ZN => n31);
   U32 : AND2_X1 port map( A1 => n87, A2 => n31, ZN => n32);
   U33 : AND2_X1 port map( A1 => n86, A2 => n32, ZN => n33);
   U34 : AND2_X1 port map( A1 => n85, A2 => n33, ZN => n34);
   U35 : AND2_X1 port map( A1 => n84, A2 => n34, ZN => n35);
   U36 : AND2_X1 port map( A1 => n83, A2 => n35, ZN => n36);
   U37 : AND2_X1 port map( A1 => n82, A2 => n36, ZN => n37);
   U38 : AND2_X1 port map( A1 => n81, A2 => n37, ZN => n38);
   U39 : AND2_X1 port map( A1 => n80, A2 => n38, ZN => n39);
   U40 : AND2_X1 port map( A1 => n79, A2 => n39, ZN => n40);
   U41 : AND2_X1 port map( A1 => n78, A2 => n40, ZN => n41);
   U42 : AND2_X1 port map( A1 => n77, A2 => n41, ZN => n42);
   U43 : AND2_X1 port map( A1 => n76, A2 => n42, ZN => n43);
   U44 : AND2_X1 port map( A1 => n75, A2 => n43, ZN => n44);
   U45 : AND2_X1 port map( A1 => n74, A2 => n44, ZN => n45);
   U46 : AND2_X1 port map( A1 => n73, A2 => n45, ZN => n46);
   U47 : AND2_X1 port map( A1 => n72, A2 => n46, ZN => n47);
   U48 : AND2_X1 port map( A1 => n71, A2 => n47, ZN => n48);
   U49 : AND2_X1 port map( A1 => n70, A2 => n48, ZN => n49);
   U50 : AND2_X1 port map( A1 => n69, A2 => n49, ZN => n50);
   U51 : AND2_X1 port map( A1 => n68, A2 => n50, ZN => n51);
   U52 : AND2_X1 port map( A1 => n67, A2 => n51, ZN => n52);
   U53 : AND2_X1 port map( A1 => n66, A2 => n52, ZN => n53);
   U54 : AND2_X1 port map( A1 => n65, A2 => n53, ZN => n54);
   U55 : XOR2_X1 port map( A => n88, B => n30, Z => DIFF_6_port);
   U56 : XOR2_X1 port map( A => n89, B => n58, Z => DIFF_5_port);
   U57 : AND2_X1 port map( A1 => n91, A2 => n59, ZN => n57);
   U58 : AND2_X1 port map( A1 => n90, A2 => n57, ZN => n58);
   U59 : AND2_X1 port map( A1 => n92, A2 => n60, ZN => n59);
   U60 : AND2_X1 port map( A1 => n63, A2 => n62, ZN => n60);
   U61 : NAND2_X1 port map( A1 => n64, A2 => n54, ZN => n61);
   U62 : INV_X1 port map( A => B(5), ZN => n89);
   U63 : INV_X1 port map( A => B(6), ZN => n88);
   U64 : INV_X1 port map( A => B(7), ZN => n87);
   U65 : INV_X1 port map( A => B(8), ZN => n86);
   U66 : INV_X1 port map( A => B(9), ZN => n85);
   U67 : INV_X1 port map( A => B(10), ZN => n84);
   U68 : INV_X1 port map( A => B(11), ZN => n83);
   U69 : INV_X1 port map( A => B(12), ZN => n82);
   U70 : INV_X1 port map( A => B(13), ZN => n81);
   U71 : INV_X1 port map( A => B(14), ZN => n80);
   U72 : INV_X1 port map( A => B(15), ZN => n79);
   U73 : INV_X1 port map( A => B(16), ZN => n78);
   U74 : INV_X1 port map( A => B(17), ZN => n77);
   U75 : INV_X1 port map( A => B(18), ZN => n76);
   U76 : INV_X1 port map( A => B(19), ZN => n75);
   U77 : INV_X1 port map( A => B(20), ZN => n74);
   U78 : INV_X1 port map( A => B(21), ZN => n73);
   U79 : INV_X1 port map( A => B(22), ZN => n72);
   U80 : INV_X1 port map( A => B(23), ZN => n71);
   U81 : INV_X1 port map( A => B(24), ZN => n70);
   U82 : INV_X1 port map( A => B(25), ZN => n69);
   U83 : INV_X1 port map( A => B(26), ZN => n68);
   U84 : INV_X1 port map( A => B(27), ZN => n67);
   U85 : INV_X1 port map( A => B(28), ZN => n66);
   U86 : INV_X1 port map( A => B(29), ZN => n65);
   U87 : INV_X1 port map( A => B(30), ZN => n64);
   U88 : INV_X1 port map( A => B(0), ZN => n62);
   U89 : INV_X1 port map( A => B(1), ZN => n63);
   U90 : INV_X1 port map( A => B(2), ZN => n92);
   U91 : INV_X1 port map( A => B(3), ZN => n91);
   U92 : INV_X1 port map( A => B(4), ZN => n90);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity negate_NBIT32_2_DW01_sub_0 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end negate_NBIT32_2_DW01_sub_0;

architecture SYN_rpl of negate_NBIT32_2_DW01_sub_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal DIFF_5_port, DIFF_4_port, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, 
      n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27
      , n28, n29, DIFF_30_port, DIFF_29_port, DIFF_28_port, DIFF_27_port, 
      DIFF_26_port, DIFF_25_port, DIFF_24_port, DIFF_23_port, DIFF_22_port, 
      DIFF_21_port, DIFF_20_port, DIFF_19_port, DIFF_18_port, DIFF_17_port, 
      DIFF_16_port, DIFF_15_port, DIFF_14_port, DIFF_13_port, DIFF_12_port, 
      DIFF_11_port, DIFF_10_port, DIFF_9_port, DIFF_8_port, DIFF_7_port, 
      DIFF_6_port, DIFF_3_port, n56, n57, DIFF_2_port, DIFF_1_port, 
      DIFF_31_port, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
      n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87
      , n88, n89, n90, n91, n92 : std_logic;

begin
   DIFF <= ( DIFF_31_port, DIFF_30_port, DIFF_29_port, DIFF_28_port, 
      DIFF_27_port, DIFF_26_port, DIFF_25_port, DIFF_24_port, DIFF_23_port, 
      DIFF_22_port, DIFF_21_port, DIFF_20_port, DIFF_19_port, DIFF_18_port, 
      DIFF_17_port, DIFF_16_port, DIFF_15_port, DIFF_14_port, DIFF_13_port, 
      DIFF_12_port, DIFF_11_port, DIFF_10_port, DIFF_9_port, DIFF_8_port, 
      DIFF_7_port, DIFF_6_port, DIFF_5_port, DIFF_4_port, DIFF_3_port, 
      DIFF_2_port, DIFF_1_port, B(0) );
   
   U1 : XOR2_X1 port map( A => n88, B => n4, Z => DIFF_5_port);
   U2 : XOR2_X1 port map( A => n89, B => n3, Z => DIFF_4_port);
   U3 : AND2_X1 port map( A1 => n90, A2 => n56, ZN => n3);
   U4 : AND2_X1 port map( A1 => n89, A2 => n3, ZN => n4);
   U5 : AND2_X1 port map( A1 => n88, A2 => n4, ZN => n5);
   U6 : AND2_X1 port map( A1 => n87, A2 => n5, ZN => n6);
   U7 : AND2_X1 port map( A1 => n86, A2 => n6, ZN => n7);
   U8 : AND2_X1 port map( A1 => n85, A2 => n7, ZN => n8);
   U9 : AND2_X1 port map( A1 => n84, A2 => n8, ZN => n9);
   U10 : AND2_X1 port map( A1 => n83, A2 => n9, ZN => n10);
   U11 : AND2_X1 port map( A1 => n82, A2 => n10, ZN => n11);
   U12 : AND2_X1 port map( A1 => n81, A2 => n11, ZN => n12);
   U13 : AND2_X1 port map( A1 => n80, A2 => n12, ZN => n13);
   U14 : AND2_X1 port map( A1 => n79, A2 => n13, ZN => n14);
   U15 : AND2_X1 port map( A1 => n78, A2 => n14, ZN => n15);
   U16 : AND2_X1 port map( A1 => n77, A2 => n15, ZN => n16);
   U17 : AND2_X1 port map( A1 => n76, A2 => n16, ZN => n17);
   U18 : AND2_X1 port map( A1 => n75, A2 => n17, ZN => n18);
   U19 : AND2_X1 port map( A1 => n74, A2 => n18, ZN => n19);
   U20 : AND2_X1 port map( A1 => n73, A2 => n19, ZN => n20);
   U21 : AND2_X1 port map( A1 => n72, A2 => n20, ZN => n21);
   U22 : AND2_X1 port map( A1 => n71, A2 => n21, ZN => n22);
   U23 : AND2_X1 port map( A1 => n70, A2 => n22, ZN => n23);
   U24 : AND2_X1 port map( A1 => n69, A2 => n23, ZN => n24);
   U25 : AND2_X1 port map( A1 => n68, A2 => n24, ZN => n25);
   U26 : AND2_X1 port map( A1 => n67, A2 => n25, ZN => n26);
   U27 : AND2_X1 port map( A1 => n66, A2 => n26, ZN => n27);
   U28 : AND2_X1 port map( A1 => n65, A2 => n27, ZN => n28);
   U29 : AND2_X1 port map( A1 => n64, A2 => n28, ZN => n29);
   U30 : NAND2_X1 port map( A1 => n63, A2 => n29, ZN => n61);
   U31 : XOR2_X1 port map( A => n63, B => n29, Z => DIFF_30_port);
   U32 : XOR2_X1 port map( A => n64, B => n28, Z => DIFF_29_port);
   U33 : XOR2_X1 port map( A => n65, B => n27, Z => DIFF_28_port);
   U34 : XOR2_X1 port map( A => n66, B => n26, Z => DIFF_27_port);
   U35 : XOR2_X1 port map( A => n67, B => n25, Z => DIFF_26_port);
   U36 : XOR2_X1 port map( A => n68, B => n24, Z => DIFF_25_port);
   U37 : XOR2_X1 port map( A => n69, B => n23, Z => DIFF_24_port);
   U38 : XOR2_X1 port map( A => n70, B => n22, Z => DIFF_23_port);
   U39 : XOR2_X1 port map( A => n71, B => n21, Z => DIFF_22_port);
   U40 : XOR2_X1 port map( A => n72, B => n20, Z => DIFF_21_port);
   U41 : XOR2_X1 port map( A => n73, B => n19, Z => DIFF_20_port);
   U42 : XOR2_X1 port map( A => n74, B => n18, Z => DIFF_19_port);
   U43 : XOR2_X1 port map( A => n75, B => n17, Z => DIFF_18_port);
   U44 : XOR2_X1 port map( A => n76, B => n16, Z => DIFF_17_port);
   U45 : XOR2_X1 port map( A => n77, B => n15, Z => DIFF_16_port);
   U46 : XOR2_X1 port map( A => n78, B => n14, Z => DIFF_15_port);
   U47 : XOR2_X1 port map( A => n79, B => n13, Z => DIFF_14_port);
   U48 : XOR2_X1 port map( A => n80, B => n12, Z => DIFF_13_port);
   U49 : XOR2_X1 port map( A => n81, B => n11, Z => DIFF_12_port);
   U50 : XOR2_X1 port map( A => n82, B => n10, Z => DIFF_11_port);
   U51 : XOR2_X1 port map( A => n83, B => n9, Z => DIFF_10_port);
   U52 : XOR2_X1 port map( A => n84, B => n8, Z => DIFF_9_port);
   U53 : XOR2_X1 port map( A => n85, B => n7, Z => DIFF_8_port);
   U54 : XOR2_X1 port map( A => n86, B => n6, Z => DIFF_7_port);
   U55 : XOR2_X1 port map( A => n87, B => n5, Z => DIFF_6_port);
   U56 : XOR2_X1 port map( A => n90, B => n56, Z => DIFF_3_port);
   U57 : AND2_X1 port map( A1 => n91, A2 => n57, ZN => n56);
   U58 : AND2_X1 port map( A1 => n92, A2 => n62, ZN => n57);
   U59 : XOR2_X1 port map( A => n91, B => n57, Z => DIFF_2_port);
   U60 : XOR2_X1 port map( A => n92, B => n62, Z => DIFF_1_port);
   U61 : INV_X1 port map( A => B(3), ZN => n90);
   U62 : INV_X1 port map( A => B(4), ZN => n89);
   U63 : INV_X1 port map( A => B(5), ZN => n88);
   U64 : INV_X1 port map( A => B(6), ZN => n87);
   U65 : INV_X1 port map( A => B(7), ZN => n86);
   U66 : INV_X1 port map( A => B(8), ZN => n85);
   U67 : INV_X1 port map( A => B(9), ZN => n84);
   U68 : INV_X1 port map( A => B(10), ZN => n83);
   U69 : INV_X1 port map( A => B(11), ZN => n82);
   U70 : INV_X1 port map( A => B(12), ZN => n81);
   U71 : INV_X1 port map( A => B(13), ZN => n80);
   U72 : XOR2_X1 port map( A => B(31), B => n61, Z => DIFF_31_port);
   U73 : INV_X1 port map( A => B(14), ZN => n79);
   U74 : INV_X1 port map( A => B(15), ZN => n78);
   U75 : INV_X1 port map( A => B(16), ZN => n77);
   U76 : INV_X1 port map( A => B(17), ZN => n76);
   U77 : INV_X1 port map( A => B(18), ZN => n75);
   U78 : INV_X1 port map( A => B(19), ZN => n74);
   U79 : INV_X1 port map( A => B(20), ZN => n73);
   U80 : INV_X1 port map( A => B(21), ZN => n72);
   U81 : INV_X1 port map( A => B(22), ZN => n71);
   U82 : INV_X1 port map( A => B(23), ZN => n70);
   U83 : INV_X1 port map( A => B(24), ZN => n69);
   U84 : INV_X1 port map( A => B(25), ZN => n68);
   U85 : INV_X1 port map( A => B(26), ZN => n67);
   U86 : INV_X1 port map( A => B(27), ZN => n66);
   U87 : INV_X1 port map( A => B(28), ZN => n65);
   U88 : INV_X1 port map( A => B(29), ZN => n64);
   U89 : INV_X1 port map( A => B(30), ZN => n63);
   U90 : INV_X1 port map( A => B(0), ZN => n62);
   U91 : INV_X1 port map( A => B(1), ZN => n92);
   U92 : INV_X1 port map( A => B(2), ZN => n91);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity negate_NBIT32_1_DW01_sub_0 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  DIFF : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end negate_NBIT32_1_DW01_sub_0;

architecture SYN_rpl of negate_NBIT32_1_DW01_sub_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal DIFF_31_port, DIFF_30_port, DIFF_29_port, DIFF_28_port, DIFF_27_port,
      DIFF_26_port, DIFF_25_port, DIFF_24_port, DIFF_23_port, DIFF_22_port, 
      DIFF_21_port, DIFF_20_port, DIFF_19_port, DIFF_18_port, DIFF_17_port, 
      DIFF_16_port, DIFF_15_port, DIFF_14_port, DIFF_13_port, DIFF_12_port, 
      DIFF_11_port, DIFF_10_port, DIFF_9_port, DIFF_8_port, DIFF_7_port, 
      DIFF_6_port, DIFF_3_port, DIFF_2_port, DIFF_1_port, n30, n31, n32, n33, 
      n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48
      , n49, n50, n51, n52, n53, n54, n55, DIFF_5_port, DIFF_4_port, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92 : std_logic;

begin
   DIFF <= ( DIFF_31_port, DIFF_30_port, DIFF_29_port, DIFF_28_port, 
      DIFF_27_port, DIFF_26_port, DIFF_25_port, DIFF_24_port, DIFF_23_port, 
      DIFF_22_port, DIFF_21_port, DIFF_20_port, DIFF_19_port, DIFF_18_port, 
      DIFF_17_port, DIFF_16_port, DIFF_15_port, DIFF_14_port, DIFF_13_port, 
      DIFF_12_port, DIFF_11_port, DIFF_10_port, DIFF_9_port, DIFF_8_port, 
      DIFF_7_port, DIFF_6_port, DIFF_5_port, DIFF_4_port, DIFF_3_port, 
      DIFF_2_port, DIFF_1_port, B(0) );
   
   U1 : XOR2_X1 port map( A => B(31), B => n61, Z => DIFF_31_port);
   U2 : XOR2_X1 port map( A => n64, B => n55, Z => DIFF_30_port);
   U3 : XOR2_X1 port map( A => n65, B => n54, Z => DIFF_29_port);
   U4 : XOR2_X1 port map( A => n66, B => n53, Z => DIFF_28_port);
   U5 : XOR2_X1 port map( A => n67, B => n52, Z => DIFF_27_port);
   U6 : XOR2_X1 port map( A => n68, B => n51, Z => DIFF_26_port);
   U7 : XOR2_X1 port map( A => n69, B => n50, Z => DIFF_25_port);
   U8 : XOR2_X1 port map( A => n70, B => n49, Z => DIFF_24_port);
   U9 : XOR2_X1 port map( A => n71, B => n48, Z => DIFF_23_port);
   U10 : XOR2_X1 port map( A => n72, B => n47, Z => DIFF_22_port);
   U11 : XOR2_X1 port map( A => n73, B => n46, Z => DIFF_21_port);
   U12 : XOR2_X1 port map( A => n74, B => n45, Z => DIFF_20_port);
   U13 : XOR2_X1 port map( A => n75, B => n44, Z => DIFF_19_port);
   U14 : XOR2_X1 port map( A => n76, B => n43, Z => DIFF_18_port);
   U15 : XOR2_X1 port map( A => n77, B => n42, Z => DIFF_17_port);
   U16 : XOR2_X1 port map( A => n78, B => n41, Z => DIFF_16_port);
   U17 : XOR2_X1 port map( A => n79, B => n40, Z => DIFF_15_port);
   U18 : XOR2_X1 port map( A => n80, B => n39, Z => DIFF_14_port);
   U19 : XOR2_X1 port map( A => n81, B => n38, Z => DIFF_13_port);
   U20 : XOR2_X1 port map( A => n82, B => n37, Z => DIFF_12_port);
   U21 : XOR2_X1 port map( A => n83, B => n36, Z => DIFF_11_port);
   U22 : XOR2_X1 port map( A => n84, B => n35, Z => DIFF_10_port);
   U23 : XOR2_X1 port map( A => n85, B => n34, Z => DIFF_9_port);
   U24 : XOR2_X1 port map( A => n86, B => n33, Z => DIFF_8_port);
   U25 : XOR2_X1 port map( A => n87, B => n32, Z => DIFF_7_port);
   U26 : XOR2_X1 port map( A => n88, B => n31, Z => DIFF_6_port);
   U27 : XOR2_X1 port map( A => n91, B => n59, Z => DIFF_3_port);
   U28 : XOR2_X1 port map( A => n92, B => n60, Z => DIFF_2_port);
   U29 : XOR2_X1 port map( A => n63, B => n62, Z => DIFF_1_port);
   U30 : AND2_X1 port map( A1 => n90, A2 => n58, ZN => n30);
   U31 : AND2_X1 port map( A1 => n89, A2 => n30, ZN => n31);
   U32 : AND2_X1 port map( A1 => n88, A2 => n31, ZN => n32);
   U33 : AND2_X1 port map( A1 => n87, A2 => n32, ZN => n33);
   U34 : AND2_X1 port map( A1 => n86, A2 => n33, ZN => n34);
   U35 : AND2_X1 port map( A1 => n85, A2 => n34, ZN => n35);
   U36 : AND2_X1 port map( A1 => n84, A2 => n35, ZN => n36);
   U37 : AND2_X1 port map( A1 => n83, A2 => n36, ZN => n37);
   U38 : AND2_X1 port map( A1 => n82, A2 => n37, ZN => n38);
   U39 : AND2_X1 port map( A1 => n81, A2 => n38, ZN => n39);
   U40 : AND2_X1 port map( A1 => n80, A2 => n39, ZN => n40);
   U41 : AND2_X1 port map( A1 => n79, A2 => n40, ZN => n41);
   U42 : AND2_X1 port map( A1 => n78, A2 => n41, ZN => n42);
   U43 : AND2_X1 port map( A1 => n77, A2 => n42, ZN => n43);
   U44 : AND2_X1 port map( A1 => n76, A2 => n43, ZN => n44);
   U45 : AND2_X1 port map( A1 => n75, A2 => n44, ZN => n45);
   U46 : AND2_X1 port map( A1 => n74, A2 => n45, ZN => n46);
   U47 : AND2_X1 port map( A1 => n73, A2 => n46, ZN => n47);
   U48 : AND2_X1 port map( A1 => n72, A2 => n47, ZN => n48);
   U49 : AND2_X1 port map( A1 => n71, A2 => n48, ZN => n49);
   U50 : AND2_X1 port map( A1 => n70, A2 => n49, ZN => n50);
   U51 : AND2_X1 port map( A1 => n69, A2 => n50, ZN => n51);
   U52 : AND2_X1 port map( A1 => n68, A2 => n51, ZN => n52);
   U53 : AND2_X1 port map( A1 => n67, A2 => n52, ZN => n53);
   U54 : AND2_X1 port map( A1 => n66, A2 => n53, ZN => n54);
   U55 : AND2_X1 port map( A1 => n65, A2 => n54, ZN => n55);
   U56 : XOR2_X1 port map( A => n89, B => n30, Z => DIFF_5_port);
   U57 : XOR2_X1 port map( A => n90, B => n58, Z => DIFF_4_port);
   U58 : AND2_X1 port map( A1 => n91, A2 => n59, ZN => n58);
   U59 : AND2_X1 port map( A1 => n92, A2 => n60, ZN => n59);
   U60 : AND2_X1 port map( A1 => n63, A2 => n62, ZN => n60);
   U61 : NAND2_X1 port map( A1 => n64, A2 => n55, ZN => n61);
   U62 : INV_X1 port map( A => B(4), ZN => n90);
   U63 : INV_X1 port map( A => B(5), ZN => n89);
   U64 : INV_X1 port map( A => B(6), ZN => n88);
   U65 : INV_X1 port map( A => B(7), ZN => n87);
   U66 : INV_X1 port map( A => B(8), ZN => n86);
   U67 : INV_X1 port map( A => B(9), ZN => n85);
   U68 : INV_X1 port map( A => B(10), ZN => n84);
   U69 : INV_X1 port map( A => B(11), ZN => n83);
   U70 : INV_X1 port map( A => B(12), ZN => n82);
   U71 : INV_X1 port map( A => B(13), ZN => n81);
   U72 : INV_X1 port map( A => B(14), ZN => n80);
   U73 : INV_X1 port map( A => B(15), ZN => n79);
   U74 : INV_X1 port map( A => B(16), ZN => n78);
   U75 : INV_X1 port map( A => B(17), ZN => n77);
   U76 : INV_X1 port map( A => B(18), ZN => n76);
   U77 : INV_X1 port map( A => B(19), ZN => n75);
   U78 : INV_X1 port map( A => B(20), ZN => n74);
   U79 : INV_X1 port map( A => B(21), ZN => n73);
   U80 : INV_X1 port map( A => B(22), ZN => n72);
   U81 : INV_X1 port map( A => B(23), ZN => n71);
   U82 : INV_X1 port map( A => B(24), ZN => n70);
   U83 : INV_X1 port map( A => B(25), ZN => n69);
   U84 : INV_X1 port map( A => B(26), ZN => n68);
   U85 : INV_X1 port map( A => B(27), ZN => n67);
   U86 : INV_X1 port map( A => B(28), ZN => n66);
   U87 : INV_X1 port map( A => B(29), ZN => n65);
   U88 : INV_X1 port map( A => B(30), ZN => n64);
   U89 : INV_X1 port map( A => B(0), ZN => n62);
   U90 : INV_X1 port map( A => B(1), ZN => n63);
   U91 : INV_X1 port map( A => B(2), ZN => n92);
   U92 : INV_X1 port map( A => B(3), ZN => n91);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX81_31 is

   port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
         downto 0);  Y : out std_logic);

end MUX81_31;

architecture SYN_BEHAVIORAL_1 of MUX81_31 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n21, n22, n23, n24, n25, n26, n27, n28, n29, 
      n30, n31, n32, n33, n34, n35 : std_logic;

begin
   
   U20 : NAND3_X1 port map( A1 => S(1), A2 => n21, A3 => H, ZN => n23);
   U21 : NAND3_X1 port map( A1 => S(0), A2 => n2, A3 => F, ZN => n25);
   U1 : INV_X1 port map( A => n27, ZN => n6);
   U2 : NOR2_X1 port map( A1 => n1, A2 => n3, ZN => n27);
   U3 : INV_X1 port map( A => n22, ZN => n21);
   U4 : AOI22_X1 port map( A1 => n33, A2 => n5, B1 => B, B2 => n32, ZN => n35);
   U5 : INV_X1 port map( A => n32, ZN => n5);
   U6 : NOR3_X1 port map( A1 => S(1), A2 => n3, A3 => n1, ZN => n32);
   U7 : OAI21_X1 port map( B1 => n31, B2 => n30, A => n29, ZN => n33);
   U8 : NAND2_X1 port map( A1 => C, A2 => n30, ZN => n29);
   U9 : AOI22_X1 port map( A1 => n28, A2 => n6, B1 => D, B2 => n27, ZN => n31);
   U10 : NOR3_X1 port map( A1 => S(0), A2 => n3, A3 => n2, ZN => n30);
   U11 : NAND4_X1 port map( A1 => n26, A2 => n25, A3 => n24, A4 => n23, ZN => 
                           n28);
   U12 : NAND4_X1 port map( A1 => E, A2 => n3, A3 => n1, A4 => n2, ZN => n26);
   U13 : NAND2_X1 port map( A1 => G, A2 => n22, ZN => n24);
   U14 : NAND2_X1 port map( A1 => n35, A2 => n34, ZN => Y);
   U15 : NOR2_X1 port map( A1 => n2, A2 => S(0), ZN => n22);
   U16 : NAND4_X1 port map( A1 => A, A2 => n1, A3 => n2, A4 => n4, ZN => n34);
   U17 : INV_X1 port map( A => S(0), ZN => n1);
   U18 : INV_X1 port map( A => S(1), ZN => n2);
   U19 : INV_X1 port map( A => n4, ZN => n3);
   U22 : INV_X1 port map( A => S(2), ZN => n4);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX81_30 is

   port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
         downto 0);  Y : out std_logic);

end MUX81_30;

architecture SYN_BEHAVIORAL_1 of MUX81_30 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n21, n22, n23, n24, n25, n26, n27, n28, n29, 
      n30, n31, n32, n33, n34, n35 : std_logic;

begin
   
   U20 : NAND3_X1 port map( A1 => S(1), A2 => n21, A3 => H, ZN => n23);
   U21 : NAND3_X1 port map( A1 => S(0), A2 => n2, A3 => F, ZN => n25);
   U1 : INV_X1 port map( A => n27, ZN => n6);
   U2 : NOR2_X1 port map( A1 => n1, A2 => n3, ZN => n27);
   U3 : NAND4_X1 port map( A1 => A, A2 => n1, A3 => n2, A4 => n4, ZN => n34);
   U4 : INV_X1 port map( A => n22, ZN => n21);
   U5 : AOI22_X1 port map( A1 => n33, A2 => n5, B1 => B, B2 => n32, ZN => n35);
   U6 : INV_X1 port map( A => n32, ZN => n5);
   U7 : NOR3_X1 port map( A1 => S(1), A2 => n3, A3 => n1, ZN => n32);
   U8 : OAI21_X1 port map( B1 => n31, B2 => n30, A => n29, ZN => n33);
   U9 : NAND2_X1 port map( A1 => C, A2 => n30, ZN => n29);
   U10 : AOI22_X1 port map( A1 => n28, A2 => n6, B1 => D, B2 => n27, ZN => n31)
                           ;
   U11 : NOR3_X1 port map( A1 => S(0), A2 => n3, A3 => n2, ZN => n30);
   U12 : NAND4_X1 port map( A1 => n26, A2 => n25, A3 => n24, A4 => n23, ZN => 
                           n28);
   U13 : NAND4_X1 port map( A1 => E, A2 => n3, A3 => n1, A4 => n2, ZN => n26);
   U14 : NAND2_X1 port map( A1 => G, A2 => n22, ZN => n24);
   U15 : NAND2_X1 port map( A1 => n35, A2 => n34, ZN => Y);
   U16 : NOR2_X1 port map( A1 => n2, A2 => S(0), ZN => n22);
   U17 : INV_X1 port map( A => S(0), ZN => n1);
   U18 : INV_X1 port map( A => S(1), ZN => n2);
   U19 : INV_X1 port map( A => n4, ZN => n3);
   U22 : INV_X1 port map( A => S(2), ZN => n4);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX81_29 is

   port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
         downto 0);  Y : out std_logic);

end MUX81_29;

architecture SYN_BEHAVIORAL_1 of MUX81_29 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n21, n22, n23, n24, n25, n26, n27, n28, n29, 
      n30, n31, n32, n33, n34, n35 : std_logic;

begin
   
   U20 : NAND3_X1 port map( A1 => S(1), A2 => n21, A3 => H, ZN => n23);
   U21 : NAND3_X1 port map( A1 => S(0), A2 => n2, A3 => F, ZN => n25);
   U1 : INV_X1 port map( A => n27, ZN => n6);
   U2 : NOR2_X1 port map( A1 => n1, A2 => n3, ZN => n27);
   U3 : NAND4_X1 port map( A1 => A, A2 => n1, A3 => n2, A4 => n4, ZN => n34);
   U4 : INV_X1 port map( A => n22, ZN => n21);
   U5 : AOI22_X1 port map( A1 => n33, A2 => n5, B1 => B, B2 => n32, ZN => n35);
   U6 : INV_X1 port map( A => n32, ZN => n5);
   U7 : NOR3_X1 port map( A1 => S(1), A2 => n3, A3 => n1, ZN => n32);
   U8 : OAI21_X1 port map( B1 => n31, B2 => n30, A => n29, ZN => n33);
   U9 : NAND2_X1 port map( A1 => C, A2 => n30, ZN => n29);
   U10 : AOI22_X1 port map( A1 => n28, A2 => n6, B1 => D, B2 => n27, ZN => n31)
                           ;
   U11 : NOR3_X1 port map( A1 => S(0), A2 => n3, A3 => n2, ZN => n30);
   U12 : NAND4_X1 port map( A1 => n26, A2 => n25, A3 => n24, A4 => n23, ZN => 
                           n28);
   U13 : NAND4_X1 port map( A1 => E, A2 => n3, A3 => n1, A4 => n2, ZN => n26);
   U14 : NAND2_X1 port map( A1 => G, A2 => n22, ZN => n24);
   U15 : NAND2_X1 port map( A1 => n35, A2 => n34, ZN => Y);
   U16 : NOR2_X1 port map( A1 => n2, A2 => S(0), ZN => n22);
   U17 : INV_X1 port map( A => S(0), ZN => n1);
   U18 : INV_X1 port map( A => S(1), ZN => n2);
   U19 : INV_X1 port map( A => n4, ZN => n3);
   U22 : INV_X1 port map( A => S(2), ZN => n4);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX81_28 is

   port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
         downto 0);  Y : out std_logic);

end MUX81_28;

architecture SYN_BEHAVIORAL_1 of MUX81_28 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n21, n22, n23, n24, n25, n26, n27, n28, n29, 
      n30, n31, n32, n33, n34, n35 : std_logic;

begin
   
   U20 : NAND3_X1 port map( A1 => S(1), A2 => n21, A3 => H, ZN => n23);
   U21 : NAND3_X1 port map( A1 => S(0), A2 => n2, A3 => F, ZN => n25);
   U1 : INV_X1 port map( A => n27, ZN => n6);
   U2 : NOR2_X1 port map( A1 => n1, A2 => n3, ZN => n27);
   U3 : NAND4_X1 port map( A1 => A, A2 => n1, A3 => n2, A4 => n4, ZN => n34);
   U4 : INV_X1 port map( A => n22, ZN => n21);
   U5 : AOI22_X1 port map( A1 => n33, A2 => n5, B1 => B, B2 => n32, ZN => n35);
   U6 : INV_X1 port map( A => n32, ZN => n5);
   U7 : NOR3_X1 port map( A1 => S(1), A2 => n3, A3 => n1, ZN => n32);
   U8 : OAI21_X1 port map( B1 => n31, B2 => n30, A => n29, ZN => n33);
   U9 : NAND2_X1 port map( A1 => C, A2 => n30, ZN => n29);
   U10 : AOI22_X1 port map( A1 => n28, A2 => n6, B1 => D, B2 => n27, ZN => n31)
                           ;
   U11 : NOR3_X1 port map( A1 => S(0), A2 => n3, A3 => n2, ZN => n30);
   U12 : NAND4_X1 port map( A1 => n26, A2 => n25, A3 => n24, A4 => n23, ZN => 
                           n28);
   U13 : NAND4_X1 port map( A1 => E, A2 => n3, A3 => n1, A4 => n2, ZN => n26);
   U14 : NAND2_X1 port map( A1 => G, A2 => n22, ZN => n24);
   U15 : NOR2_X1 port map( A1 => n2, A2 => S(0), ZN => n22);
   U16 : NAND2_X1 port map( A1 => n35, A2 => n34, ZN => Y);
   U17 : INV_X1 port map( A => S(0), ZN => n1);
   U18 : INV_X1 port map( A => S(1), ZN => n2);
   U19 : INV_X1 port map( A => n4, ZN => n3);
   U22 : INV_X1 port map( A => S(2), ZN => n4);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX81_27 is

   port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
         downto 0);  Y : out std_logic);

end MUX81_27;

architecture SYN_BEHAVIORAL_1 of MUX81_27 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n21, n22, n23, n24, n25, n26, n27, n28, n29, 
      n30, n31, n32, n33, n34, n35 : std_logic;

begin
   
   U20 : NAND3_X1 port map( A1 => S(1), A2 => n21, A3 => H, ZN => n23);
   U21 : NAND3_X1 port map( A1 => S(0), A2 => n2, A3 => F, ZN => n25);
   U1 : INV_X1 port map( A => n27, ZN => n6);
   U2 : NOR2_X1 port map( A1 => n1, A2 => n3, ZN => n27);
   U3 : NAND4_X1 port map( A1 => A, A2 => n1, A3 => n2, A4 => n4, ZN => n34);
   U4 : INV_X1 port map( A => n22, ZN => n21);
   U5 : AOI22_X1 port map( A1 => n33, A2 => n5, B1 => B, B2 => n32, ZN => n35);
   U6 : INV_X1 port map( A => n32, ZN => n5);
   U7 : NOR3_X1 port map( A1 => S(1), A2 => n3, A3 => n1, ZN => n32);
   U8 : OAI21_X1 port map( B1 => n31, B2 => n30, A => n29, ZN => n33);
   U9 : NAND2_X1 port map( A1 => C, A2 => n30, ZN => n29);
   U10 : AOI22_X1 port map( A1 => n28, A2 => n6, B1 => D, B2 => n27, ZN => n31)
                           ;
   U11 : NOR3_X1 port map( A1 => S(0), A2 => n3, A3 => n2, ZN => n30);
   U12 : NAND4_X1 port map( A1 => n26, A2 => n25, A3 => n24, A4 => n23, ZN => 
                           n28);
   U13 : NAND4_X1 port map( A1 => E, A2 => n3, A3 => n1, A4 => n2, ZN => n26);
   U14 : NAND2_X1 port map( A1 => G, A2 => n22, ZN => n24);
   U15 : NAND2_X1 port map( A1 => n35, A2 => n34, ZN => Y);
   U16 : NOR2_X1 port map( A1 => n2, A2 => S(0), ZN => n22);
   U17 : INV_X1 port map( A => S(0), ZN => n1);
   U18 : INV_X1 port map( A => S(1), ZN => n2);
   U19 : INV_X1 port map( A => n4, ZN => n3);
   U22 : INV_X1 port map( A => S(2), ZN => n4);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX81_26 is

   port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
         downto 0);  Y : out std_logic);

end MUX81_26;

architecture SYN_BEHAVIORAL_1 of MUX81_26 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n21, n22, n23, n24, n25, n26, n27, n28, n29, 
      n30, n31, n32, n33, n34, n35 : std_logic;

begin
   
   U20 : NAND3_X1 port map( A1 => S(1), A2 => n21, A3 => H, ZN => n23);
   U21 : NAND3_X1 port map( A1 => S(0), A2 => n2, A3 => F, ZN => n25);
   U1 : INV_X1 port map( A => n27, ZN => n6);
   U2 : NAND2_X1 port map( A1 => G, A2 => n22, ZN => n24);
   U3 : NOR2_X1 port map( A1 => n1, A2 => n3, ZN => n27);
   U4 : NAND4_X1 port map( A1 => A, A2 => n1, A3 => n2, A4 => n4, ZN => n34);
   U5 : INV_X1 port map( A => n22, ZN => n21);
   U6 : AOI22_X1 port map( A1 => n33, A2 => n5, B1 => B, B2 => n32, ZN => n35);
   U7 : INV_X1 port map( A => n32, ZN => n5);
   U8 : NOR3_X1 port map( A1 => S(1), A2 => n3, A3 => n1, ZN => n32);
   U9 : OAI21_X1 port map( B1 => n31, B2 => n30, A => n29, ZN => n33);
   U10 : NAND2_X1 port map( A1 => C, A2 => n30, ZN => n29);
   U11 : AOI22_X1 port map( A1 => n28, A2 => n6, B1 => D, B2 => n27, ZN => n31)
                           ;
   U12 : NOR3_X1 port map( A1 => S(0), A2 => n3, A3 => n2, ZN => n30);
   U13 : NAND4_X1 port map( A1 => n26, A2 => n25, A3 => n24, A4 => n23, ZN => 
                           n28);
   U14 : NAND4_X1 port map( A1 => E, A2 => n3, A3 => n1, A4 => n2, ZN => n26);
   U15 : NAND2_X1 port map( A1 => n35, A2 => n34, ZN => Y);
   U16 : NOR2_X1 port map( A1 => n2, A2 => S(0), ZN => n22);
   U17 : INV_X1 port map( A => S(0), ZN => n1);
   U18 : INV_X1 port map( A => S(1), ZN => n2);
   U19 : INV_X1 port map( A => n4, ZN => n3);
   U22 : INV_X1 port map( A => S(2), ZN => n4);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX81_25 is

   port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
         downto 0);  Y : out std_logic);

end MUX81_25;

architecture SYN_BEHAVIORAL_1 of MUX81_25 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n21, n22, n23, n24, n25, n26, n27, n28, n29, 
      n30, n31, n32, n33, n34, n35 : std_logic;

begin
   
   U20 : NAND3_X1 port map( A1 => S(1), A2 => n21, A3 => H, ZN => n23);
   U21 : NAND3_X1 port map( A1 => S(0), A2 => n2, A3 => F, ZN => n25);
   U1 : INV_X1 port map( A => n27, ZN => n6);
   U2 : NOR2_X1 port map( A1 => n1, A2 => n3, ZN => n27);
   U3 : NAND4_X1 port map( A1 => A, A2 => n1, A3 => n2, A4 => n4, ZN => n34);
   U4 : INV_X1 port map( A => n22, ZN => n21);
   U5 : AOI22_X1 port map( A1 => n33, A2 => n5, B1 => B, B2 => n32, ZN => n35);
   U6 : INV_X1 port map( A => n32, ZN => n5);
   U7 : NOR3_X1 port map( A1 => S(1), A2 => n3, A3 => n1, ZN => n32);
   U8 : OAI21_X1 port map( B1 => n31, B2 => n30, A => n29, ZN => n33);
   U9 : NAND2_X1 port map( A1 => C, A2 => n30, ZN => n29);
   U10 : AOI22_X1 port map( A1 => n28, A2 => n6, B1 => D, B2 => n27, ZN => n31)
                           ;
   U11 : NOR3_X1 port map( A1 => S(0), A2 => n3, A3 => n2, ZN => n30);
   U12 : NAND4_X1 port map( A1 => n26, A2 => n25, A3 => n24, A4 => n23, ZN => 
                           n28);
   U13 : NAND4_X1 port map( A1 => E, A2 => n3, A3 => n1, A4 => n2, ZN => n26);
   U14 : NAND2_X1 port map( A1 => G, A2 => n22, ZN => n24);
   U15 : NAND2_X1 port map( A1 => n35, A2 => n34, ZN => Y);
   U16 : NOR2_X1 port map( A1 => n2, A2 => S(0), ZN => n22);
   U17 : INV_X1 port map( A => S(0), ZN => n1);
   U18 : INV_X1 port map( A => S(1), ZN => n2);
   U19 : INV_X1 port map( A => n4, ZN => n3);
   U22 : INV_X1 port map( A => S(2), ZN => n4);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX81_24 is

   port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
         downto 0);  Y : out std_logic);

end MUX81_24;

architecture SYN_BEHAVIORAL_1 of MUX81_24 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n21, n22, n23, n24, n25, n26, n27, n28, n29, 
      n30, n31, n32, n33, n34, n35 : std_logic;

begin
   
   U20 : NAND3_X1 port map( A1 => S(1), A2 => n21, A3 => H, ZN => n23);
   U21 : NAND3_X1 port map( A1 => S(0), A2 => n2, A3 => F, ZN => n25);
   U1 : INV_X1 port map( A => n27, ZN => n6);
   U2 : NOR2_X1 port map( A1 => n1, A2 => n3, ZN => n27);
   U3 : NAND4_X1 port map( A1 => A, A2 => n1, A3 => n2, A4 => n4, ZN => n34);
   U4 : INV_X1 port map( A => n22, ZN => n21);
   U5 : AOI22_X1 port map( A1 => n33, A2 => n5, B1 => B, B2 => n32, ZN => n35);
   U6 : INV_X1 port map( A => n32, ZN => n5);
   U7 : NOR3_X1 port map( A1 => S(1), A2 => n3, A3 => n1, ZN => n32);
   U8 : OAI21_X1 port map( B1 => n31, B2 => n30, A => n29, ZN => n33);
   U9 : NAND2_X1 port map( A1 => C, A2 => n30, ZN => n29);
   U10 : AOI22_X1 port map( A1 => n28, A2 => n6, B1 => D, B2 => n27, ZN => n31)
                           ;
   U11 : NOR3_X1 port map( A1 => S(0), A2 => n3, A3 => n2, ZN => n30);
   U12 : NAND4_X1 port map( A1 => n26, A2 => n25, A3 => n24, A4 => n23, ZN => 
                           n28);
   U13 : NAND4_X1 port map( A1 => E, A2 => n3, A3 => n1, A4 => n2, ZN => n26);
   U14 : NAND2_X1 port map( A1 => G, A2 => n22, ZN => n24);
   U15 : NOR2_X1 port map( A1 => n2, A2 => S(0), ZN => n22);
   U16 : NAND2_X1 port map( A1 => n35, A2 => n34, ZN => Y);
   U17 : INV_X1 port map( A => S(0), ZN => n1);
   U18 : INV_X1 port map( A => S(1), ZN => n2);
   U19 : INV_X1 port map( A => n4, ZN => n3);
   U22 : INV_X1 port map( A => S(2), ZN => n4);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX81_23 is

   port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
         downto 0);  Y : out std_logic);

end MUX81_23;

architecture SYN_BEHAVIORAL_1 of MUX81_23 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n21, n22, n23, n24, n25, n26, n27, n28, n29, 
      n30, n31, n32, n33, n34 : std_logic;

begin
   
   U20 : NAND3_X1 port map( A1 => S(1), A2 => n6, A3 => H, ZN => n22);
   U21 : NAND3_X1 port map( A1 => S(0), A2 => n2, A3 => F, ZN => n24);
   U1 : INV_X1 port map( A => n26, ZN => n5);
   U2 : NAND2_X1 port map( A1 => G, A2 => n21, ZN => n23);
   U3 : NOR2_X1 port map( A1 => n1, A2 => S(2), ZN => n26);
   U4 : NAND4_X1 port map( A1 => A, A2 => n1, A3 => n2, A4 => n3, ZN => n33);
   U5 : INV_X1 port map( A => n21, ZN => n6);
   U6 : AOI22_X1 port map( A1 => n32, A2 => n4, B1 => B, B2 => n31, ZN => n34);
   U7 : INV_X1 port map( A => n31, ZN => n4);
   U8 : NOR3_X1 port map( A1 => S(1), A2 => S(2), A3 => n1, ZN => n31);
   U9 : OAI21_X1 port map( B1 => n30, B2 => n29, A => n28, ZN => n32);
   U10 : NAND2_X1 port map( A1 => C, A2 => n29, ZN => n28);
   U11 : AOI22_X1 port map( A1 => n27, A2 => n5, B1 => D, B2 => n26, ZN => n30)
                           ;
   U12 : NOR3_X1 port map( A1 => S(0), A2 => S(2), A3 => n2, ZN => n29);
   U13 : NAND4_X1 port map( A1 => n25, A2 => n24, A3 => n23, A4 => n22, ZN => 
                           n27);
   U14 : NAND4_X1 port map( A1 => E, A2 => S(2), A3 => n1, A4 => n2, ZN => n25)
                           ;
   U15 : NAND2_X1 port map( A1 => n34, A2 => n33, ZN => Y);
   U16 : NOR2_X1 port map( A1 => n2, A2 => S(0), ZN => n21);
   U17 : INV_X1 port map( A => S(0), ZN => n1);
   U18 : INV_X1 port map( A => S(1), ZN => n2);
   U19 : INV_X1 port map( A => S(2), ZN => n3);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX81_22 is

   port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
         downto 0);  Y : out std_logic);

end MUX81_22;

architecture SYN_BEHAVIORAL_1 of MUX81_22 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n21, n22, n23, n24, n25, n26, n27, n28, n29, 
      n30, n31, n32, n33, n34 : std_logic;

begin
   
   U20 : NAND3_X1 port map( A1 => S(1), A2 => n6, A3 => H, ZN => n22);
   U21 : NAND3_X1 port map( A1 => S(0), A2 => n2, A3 => F, ZN => n24);
   U1 : INV_X1 port map( A => n26, ZN => n5);
   U2 : NAND2_X1 port map( A1 => G, A2 => n21, ZN => n23);
   U3 : NOR2_X1 port map( A1 => n1, A2 => S(2), ZN => n26);
   U4 : NAND4_X1 port map( A1 => A, A2 => n1, A3 => n2, A4 => n3, ZN => n33);
   U5 : INV_X1 port map( A => n21, ZN => n6);
   U6 : NAND2_X1 port map( A1 => n34, A2 => n33, ZN => Y);
   U7 : AOI22_X1 port map( A1 => n32, A2 => n4, B1 => B, B2 => n31, ZN => n34);
   U8 : INV_X1 port map( A => n31, ZN => n4);
   U9 : NOR3_X1 port map( A1 => S(1), A2 => S(2), A3 => n1, ZN => n31);
   U10 : OAI21_X1 port map( B1 => n30, B2 => n29, A => n28, ZN => n32);
   U11 : NAND2_X1 port map( A1 => C, A2 => n29, ZN => n28);
   U12 : AOI22_X1 port map( A1 => n27, A2 => n5, B1 => D, B2 => n26, ZN => n30)
                           ;
   U13 : NOR3_X1 port map( A1 => S(0), A2 => S(2), A3 => n2, ZN => n29);
   U14 : NAND4_X1 port map( A1 => n25, A2 => n24, A3 => n23, A4 => n22, ZN => 
                           n27);
   U15 : NAND4_X1 port map( A1 => E, A2 => S(2), A3 => n1, A4 => n2, ZN => n25)
                           ;
   U16 : NOR2_X1 port map( A1 => n2, A2 => S(0), ZN => n21);
   U17 : INV_X1 port map( A => S(0), ZN => n1);
   U18 : INV_X1 port map( A => S(1), ZN => n2);
   U19 : INV_X1 port map( A => S(2), ZN => n3);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX81_21 is

   port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
         downto 0);  Y : out std_logic);

end MUX81_21;

architecture SYN_BEHAVIORAL_1 of MUX81_21 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n21, n22, n23, n24, n25, n26, n27, n28, n29, 
      n30, n31, n32, n33, n34 : std_logic;

begin
   
   U20 : NAND3_X1 port map( A1 => S(1), A2 => n6, A3 => H, ZN => n22);
   U21 : NAND3_X1 port map( A1 => S(0), A2 => n2, A3 => F, ZN => n24);
   U1 : INV_X1 port map( A => n26, ZN => n5);
   U2 : NOR2_X1 port map( A1 => n1, A2 => S(2), ZN => n26);
   U3 : NAND4_X1 port map( A1 => A, A2 => n1, A3 => n2, A4 => n3, ZN => n33);
   U4 : NAND2_X1 port map( A1 => n34, A2 => n33, ZN => Y);
   U5 : INV_X1 port map( A => n21, ZN => n6);
   U6 : AOI22_X1 port map( A1 => n32, A2 => n4, B1 => B, B2 => n31, ZN => n34);
   U7 : INV_X1 port map( A => n31, ZN => n4);
   U8 : NOR3_X1 port map( A1 => S(1), A2 => S(2), A3 => n1, ZN => n31);
   U9 : OAI21_X1 port map( B1 => n30, B2 => n29, A => n28, ZN => n32);
   U10 : NAND2_X1 port map( A1 => C, A2 => n29, ZN => n28);
   U11 : AOI22_X1 port map( A1 => n27, A2 => n5, B1 => D, B2 => n26, ZN => n30)
                           ;
   U12 : NOR3_X1 port map( A1 => S(0), A2 => S(2), A3 => n2, ZN => n29);
   U13 : NAND4_X1 port map( A1 => n25, A2 => n24, A3 => n23, A4 => n22, ZN => 
                           n27);
   U14 : NAND4_X1 port map( A1 => E, A2 => S(2), A3 => n1, A4 => n2, ZN => n25)
                           ;
   U15 : NAND2_X1 port map( A1 => G, A2 => n21, ZN => n23);
   U16 : NOR2_X1 port map( A1 => n2, A2 => S(0), ZN => n21);
   U17 : INV_X1 port map( A => S(0), ZN => n1);
   U18 : INV_X1 port map( A => S(1), ZN => n2);
   U19 : INV_X1 port map( A => S(2), ZN => n3);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX81_20 is

   port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
         downto 0);  Y : out std_logic);

end MUX81_20;

architecture SYN_BEHAVIORAL_1 of MUX81_20 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n21, n22, n23, n24, n25, n26, n27, n28, n29, 
      n30, n31, n32, n33, n34, n35 : std_logic;

begin
   
   U20 : NAND3_X1 port map( A1 => S(1), A2 => n21, A3 => H, ZN => n23);
   U21 : NAND3_X1 port map( A1 => S(0), A2 => n2, A3 => F, ZN => n25);
   U1 : INV_X1 port map( A => n27, ZN => n6);
   U2 : NOR2_X1 port map( A1 => n1, A2 => n3, ZN => n27);
   U3 : NAND4_X1 port map( A1 => A, A2 => n1, A3 => n2, A4 => n4, ZN => n34);
   U4 : INV_X1 port map( A => n22, ZN => n21);
   U5 : AOI22_X1 port map( A1 => n33, A2 => n5, B1 => B, B2 => n32, ZN => n35);
   U6 : INV_X1 port map( A => n32, ZN => n5);
   U7 : NOR3_X1 port map( A1 => S(1), A2 => n3, A3 => n1, ZN => n32);
   U8 : OAI21_X1 port map( B1 => n31, B2 => n30, A => n29, ZN => n33);
   U9 : NAND2_X1 port map( A1 => C, A2 => n30, ZN => n29);
   U10 : AOI22_X1 port map( A1 => n28, A2 => n6, B1 => D, B2 => n27, ZN => n31)
                           ;
   U11 : NOR3_X1 port map( A1 => S(0), A2 => n3, A3 => n2, ZN => n30);
   U12 : NAND4_X1 port map( A1 => n26, A2 => n25, A3 => n24, A4 => n23, ZN => 
                           n28);
   U13 : NAND4_X1 port map( A1 => E, A2 => n3, A3 => n1, A4 => n2, ZN => n26);
   U14 : NAND2_X1 port map( A1 => G, A2 => n22, ZN => n24);
   U15 : NOR2_X1 port map( A1 => n2, A2 => S(0), ZN => n22);
   U16 : NAND2_X1 port map( A1 => n35, A2 => n34, ZN => Y);
   U17 : INV_X1 port map( A => S(0), ZN => n1);
   U18 : INV_X1 port map( A => S(1), ZN => n2);
   U19 : INV_X1 port map( A => n4, ZN => n3);
   U22 : INV_X1 port map( A => S(2), ZN => n4);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX81_19 is

   port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
         downto 0);  Y : out std_logic);

end MUX81_19;

architecture SYN_BEHAVIORAL_1 of MUX81_19 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n21, n22, n23, n24, n25, n26, n27, n28, n29, 
      n30, n31, n32, n33, n34, n35 : std_logic;

begin
   
   U20 : NAND3_X1 port map( A1 => S(1), A2 => n21, A3 => H, ZN => n23);
   U21 : NAND3_X1 port map( A1 => S(0), A2 => n2, A3 => F, ZN => n25);
   U1 : INV_X1 port map( A => n27, ZN => n6);
   U2 : NOR2_X1 port map( A1 => n1, A2 => n3, ZN => n27);
   U3 : NAND4_X1 port map( A1 => A, A2 => n1, A3 => n2, A4 => n4, ZN => n34);
   U4 : NAND2_X1 port map( A1 => n35, A2 => n34, ZN => Y);
   U5 : INV_X1 port map( A => n22, ZN => n21);
   U6 : AOI22_X1 port map( A1 => n33, A2 => n5, B1 => B, B2 => n32, ZN => n35);
   U7 : INV_X1 port map( A => n32, ZN => n5);
   U8 : NOR3_X1 port map( A1 => S(1), A2 => n3, A3 => n1, ZN => n32);
   U9 : OAI21_X1 port map( B1 => n31, B2 => n30, A => n29, ZN => n33);
   U10 : NAND2_X1 port map( A1 => C, A2 => n30, ZN => n29);
   U11 : AOI22_X1 port map( A1 => n28, A2 => n6, B1 => D, B2 => n27, ZN => n31)
                           ;
   U12 : NOR3_X1 port map( A1 => S(0), A2 => n3, A3 => n2, ZN => n30);
   U13 : NAND4_X1 port map( A1 => n26, A2 => n25, A3 => n24, A4 => n23, ZN => 
                           n28);
   U14 : NAND4_X1 port map( A1 => E, A2 => n3, A3 => n1, A4 => n2, ZN => n26);
   U15 : NAND2_X1 port map( A1 => G, A2 => n22, ZN => n24);
   U16 : NOR2_X1 port map( A1 => n2, A2 => S(0), ZN => n22);
   U17 : INV_X1 port map( A => S(0), ZN => n1);
   U18 : INV_X1 port map( A => S(1), ZN => n2);
   U19 : INV_X1 port map( A => n4, ZN => n3);
   U22 : INV_X1 port map( A => S(2), ZN => n4);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX81_18 is

   port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
         downto 0);  Y : out std_logic);

end MUX81_18;

architecture SYN_BEHAVIORAL_1 of MUX81_18 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n21, n22, n23, n24, n25, n26, n27, n28, n29, 
      n30, n31, n32, n33, n34, n35 : std_logic;

begin
   
   U20 : NAND3_X1 port map( A1 => S(1), A2 => n21, A3 => H, ZN => n23);
   U21 : NAND3_X1 port map( A1 => S(0), A2 => n2, A3 => F, ZN => n25);
   U1 : INV_X1 port map( A => n27, ZN => n6);
   U2 : NOR2_X1 port map( A1 => n1, A2 => n3, ZN => n27);
   U3 : NAND4_X1 port map( A1 => A, A2 => n1, A3 => n2, A4 => n4, ZN => n34);
   U4 : NAND2_X1 port map( A1 => n35, A2 => n34, ZN => Y);
   U5 : INV_X1 port map( A => n22, ZN => n21);
   U6 : AOI22_X1 port map( A1 => n33, A2 => n5, B1 => B, B2 => n32, ZN => n35);
   U7 : INV_X1 port map( A => n32, ZN => n5);
   U8 : NOR3_X1 port map( A1 => S(1), A2 => n3, A3 => n1, ZN => n32);
   U9 : OAI21_X1 port map( B1 => n31, B2 => n30, A => n29, ZN => n33);
   U10 : NAND2_X1 port map( A1 => C, A2 => n30, ZN => n29);
   U11 : AOI22_X1 port map( A1 => n28, A2 => n6, B1 => D, B2 => n27, ZN => n31)
                           ;
   U12 : NOR3_X1 port map( A1 => S(0), A2 => n3, A3 => n2, ZN => n30);
   U13 : NAND4_X1 port map( A1 => n26, A2 => n25, A3 => n24, A4 => n23, ZN => 
                           n28);
   U14 : NAND4_X1 port map( A1 => E, A2 => n3, A3 => n1, A4 => n2, ZN => n26);
   U15 : NAND2_X1 port map( A1 => G, A2 => n22, ZN => n24);
   U16 : NOR2_X1 port map( A1 => n2, A2 => S(0), ZN => n22);
   U17 : INV_X1 port map( A => S(0), ZN => n1);
   U18 : INV_X1 port map( A => S(1), ZN => n2);
   U19 : INV_X1 port map( A => n4, ZN => n3);
   U22 : INV_X1 port map( A => S(2), ZN => n4);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX81_17 is

   port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
         downto 0);  Y : out std_logic);

end MUX81_17;

architecture SYN_BEHAVIORAL_1 of MUX81_17 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n21, n22, n23, n24, n25, n26, n27, n28, n29, 
      n30, n31, n32, n33, n34, n35 : std_logic;

begin
   
   U20 : NAND3_X1 port map( A1 => S(1), A2 => n21, A3 => H, ZN => n23);
   U21 : NAND3_X1 port map( A1 => S(0), A2 => n2, A3 => F, ZN => n25);
   U1 : INV_X1 port map( A => n27, ZN => n6);
   U2 : NOR2_X1 port map( A1 => n1, A2 => n3, ZN => n27);
   U3 : NAND4_X1 port map( A1 => A, A2 => n1, A3 => n2, A4 => n4, ZN => n34);
   U4 : NAND2_X1 port map( A1 => n35, A2 => n34, ZN => Y);
   U5 : INV_X1 port map( A => n22, ZN => n21);
   U6 : AOI22_X1 port map( A1 => n33, A2 => n5, B1 => B, B2 => n32, ZN => n35);
   U7 : INV_X1 port map( A => n32, ZN => n5);
   U8 : NOR3_X1 port map( A1 => S(1), A2 => n3, A3 => n1, ZN => n32);
   U9 : OAI21_X1 port map( B1 => n31, B2 => n30, A => n29, ZN => n33);
   U10 : NAND2_X1 port map( A1 => C, A2 => n30, ZN => n29);
   U11 : AOI22_X1 port map( A1 => n28, A2 => n6, B1 => D, B2 => n27, ZN => n31)
                           ;
   U12 : NOR3_X1 port map( A1 => S(0), A2 => n3, A3 => n2, ZN => n30);
   U13 : NAND4_X1 port map( A1 => n26, A2 => n25, A3 => n24, A4 => n23, ZN => 
                           n28);
   U14 : NAND4_X1 port map( A1 => E, A2 => n3, A3 => n1, A4 => n2, ZN => n26);
   U15 : NAND2_X1 port map( A1 => G, A2 => n22, ZN => n24);
   U16 : NOR2_X1 port map( A1 => n2, A2 => S(0), ZN => n22);
   U17 : INV_X1 port map( A => S(0), ZN => n1);
   U18 : INV_X1 port map( A => S(1), ZN => n2);
   U19 : INV_X1 port map( A => n4, ZN => n3);
   U22 : INV_X1 port map( A => S(2), ZN => n4);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX81_16 is

   port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
         downto 0);  Y : out std_logic);

end MUX81_16;

architecture SYN_BEHAVIORAL_1 of MUX81_16 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n21, n22, n23, n24, n25, n26, n27, n28, n29, 
      n30, n31, n32, n33, n34, n35 : std_logic;

begin
   
   U20 : NAND3_X1 port map( A1 => S(1), A2 => n21, A3 => H, ZN => n23);
   U21 : NAND3_X1 port map( A1 => S(0), A2 => n2, A3 => F, ZN => n25);
   U1 : INV_X1 port map( A => n27, ZN => n6);
   U2 : NOR2_X1 port map( A1 => n1, A2 => n3, ZN => n27);
   U3 : NAND4_X1 port map( A1 => A, A2 => n1, A3 => n2, A4 => n4, ZN => n34);
   U4 : INV_X1 port map( A => n22, ZN => n21);
   U5 : AOI22_X1 port map( A1 => n33, A2 => n5, B1 => B, B2 => n32, ZN => n35);
   U6 : INV_X1 port map( A => n32, ZN => n5);
   U7 : NOR3_X1 port map( A1 => S(1), A2 => n3, A3 => n1, ZN => n32);
   U8 : OAI21_X1 port map( B1 => n31, B2 => n30, A => n29, ZN => n33);
   U9 : NAND2_X1 port map( A1 => C, A2 => n30, ZN => n29);
   U10 : AOI22_X1 port map( A1 => n28, A2 => n6, B1 => D, B2 => n27, ZN => n31)
                           ;
   U11 : NOR3_X1 port map( A1 => S(0), A2 => n3, A3 => n2, ZN => n30);
   U12 : NAND4_X1 port map( A1 => n26, A2 => n25, A3 => n24, A4 => n23, ZN => 
                           n28);
   U13 : NAND4_X1 port map( A1 => E, A2 => n3, A3 => n1, A4 => n2, ZN => n26);
   U14 : NAND2_X1 port map( A1 => G, A2 => n22, ZN => n24);
   U15 : NOR2_X1 port map( A1 => n2, A2 => S(0), ZN => n22);
   U16 : NAND2_X1 port map( A1 => n35, A2 => n34, ZN => Y);
   U17 : INV_X1 port map( A => S(0), ZN => n1);
   U18 : INV_X1 port map( A => S(1), ZN => n2);
   U19 : INV_X1 port map( A => n4, ZN => n3);
   U22 : INV_X1 port map( A => S(2), ZN => n4);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX81_15 is

   port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
         downto 0);  Y : out std_logic);

end MUX81_15;

architecture SYN_BEHAVIORAL_1 of MUX81_15 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n21, n22, n23, n24, n25, n26, n27, n28, n29, 
      n30, n31, n32, n33, n34, n35 : std_logic;

begin
   
   U20 : NAND3_X1 port map( A1 => S(1), A2 => n21, A3 => H, ZN => n23);
   U21 : NAND3_X1 port map( A1 => S(0), A2 => n2, A3 => F, ZN => n25);
   U1 : INV_X1 port map( A => n27, ZN => n6);
   U2 : NOR2_X1 port map( A1 => n1, A2 => n3, ZN => n27);
   U3 : NAND4_X1 port map( A1 => A, A2 => n1, A3 => n2, A4 => n4, ZN => n34);
   U4 : INV_X1 port map( A => n22, ZN => n21);
   U5 : AOI22_X1 port map( A1 => n33, A2 => n5, B1 => B, B2 => n32, ZN => n35);
   U6 : INV_X1 port map( A => n32, ZN => n5);
   U7 : NOR3_X1 port map( A1 => S(1), A2 => n3, A3 => n1, ZN => n32);
   U8 : OAI21_X1 port map( B1 => n31, B2 => n30, A => n29, ZN => n33);
   U9 : NAND2_X1 port map( A1 => C, A2 => n30, ZN => n29);
   U10 : AOI22_X1 port map( A1 => n28, A2 => n6, B1 => D, B2 => n27, ZN => n31)
                           ;
   U11 : NOR3_X1 port map( A1 => S(0), A2 => n3, A3 => n2, ZN => n30);
   U12 : NAND4_X1 port map( A1 => n26, A2 => n25, A3 => n24, A4 => n23, ZN => 
                           n28);
   U13 : NAND4_X1 port map( A1 => E, A2 => n3, A3 => n1, A4 => n2, ZN => n26);
   U14 : NAND2_X1 port map( A1 => G, A2 => n22, ZN => n24);
   U15 : NAND2_X1 port map( A1 => n35, A2 => n34, ZN => Y);
   U16 : NOR2_X1 port map( A1 => n2, A2 => S(0), ZN => n22);
   U17 : INV_X1 port map( A => S(0), ZN => n1);
   U18 : INV_X1 port map( A => S(1), ZN => n2);
   U19 : INV_X1 port map( A => n4, ZN => n3);
   U22 : INV_X1 port map( A => S(2), ZN => n4);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX81_14 is

   port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
         downto 0);  Y : out std_logic);

end MUX81_14;

architecture SYN_BEHAVIORAL_1 of MUX81_14 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n21, n22, n23, n24, n25, n26, n27, n28, n29, 
      n30, n31, n32, n33, n34, n35 : std_logic;

begin
   
   U20 : NAND3_X1 port map( A1 => S(1), A2 => n21, A3 => H, ZN => n23);
   U21 : NAND3_X1 port map( A1 => S(0), A2 => n2, A3 => F, ZN => n25);
   U1 : INV_X1 port map( A => n27, ZN => n6);
   U2 : NAND2_X1 port map( A1 => G, A2 => n22, ZN => n24);
   U3 : NOR2_X1 port map( A1 => n1, A2 => n3, ZN => n27);
   U4 : NAND4_X1 port map( A1 => A, A2 => n1, A3 => n2, A4 => n4, ZN => n34);
   U5 : INV_X1 port map( A => n22, ZN => n21);
   U6 : AOI22_X1 port map( A1 => n33, A2 => n5, B1 => B, B2 => n32, ZN => n35);
   U7 : INV_X1 port map( A => n32, ZN => n5);
   U8 : NOR3_X1 port map( A1 => S(1), A2 => n3, A3 => n1, ZN => n32);
   U9 : OAI21_X1 port map( B1 => n31, B2 => n30, A => n29, ZN => n33);
   U10 : NAND2_X1 port map( A1 => C, A2 => n30, ZN => n29);
   U11 : AOI22_X1 port map( A1 => n28, A2 => n6, B1 => D, B2 => n27, ZN => n31)
                           ;
   U12 : NOR3_X1 port map( A1 => S(0), A2 => n3, A3 => n2, ZN => n30);
   U13 : NAND4_X1 port map( A1 => n26, A2 => n25, A3 => n24, A4 => n23, ZN => 
                           n28);
   U14 : NAND4_X1 port map( A1 => E, A2 => n3, A3 => n1, A4 => n2, ZN => n26);
   U15 : NAND2_X1 port map( A1 => n35, A2 => n34, ZN => Y);
   U16 : NOR2_X1 port map( A1 => n2, A2 => S(0), ZN => n22);
   U17 : INV_X1 port map( A => S(0), ZN => n1);
   U18 : INV_X1 port map( A => S(1), ZN => n2);
   U19 : INV_X1 port map( A => n4, ZN => n3);
   U22 : INV_X1 port map( A => S(2), ZN => n4);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX81_13 is

   port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
         downto 0);  Y : out std_logic);

end MUX81_13;

architecture SYN_BEHAVIORAL_1 of MUX81_13 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n21, n22, n23, n24, n25, n26, n27, n28, n29, 
      n30, n31, n32, n33, n34, n35 : std_logic;

begin
   
   U20 : NAND3_X1 port map( A1 => S(1), A2 => n21, A3 => H, ZN => n23);
   U21 : NAND3_X1 port map( A1 => S(0), A2 => n2, A3 => F, ZN => n25);
   U1 : INV_X1 port map( A => n27, ZN => n6);
   U2 : NAND2_X1 port map( A1 => G, A2 => n22, ZN => n24);
   U3 : NOR2_X1 port map( A1 => n1, A2 => n3, ZN => n27);
   U4 : NAND4_X1 port map( A1 => A, A2 => n1, A3 => n2, A4 => n4, ZN => n34);
   U5 : INV_X1 port map( A => n22, ZN => n21);
   U6 : NAND2_X1 port map( A1 => n35, A2 => n34, ZN => Y);
   U7 : AOI22_X1 port map( A1 => n33, A2 => n5, B1 => B, B2 => n32, ZN => n35);
   U8 : INV_X1 port map( A => n32, ZN => n5);
   U9 : NOR3_X1 port map( A1 => S(1), A2 => n3, A3 => n1, ZN => n32);
   U10 : OAI21_X1 port map( B1 => n31, B2 => n30, A => n29, ZN => n33);
   U11 : NAND2_X1 port map( A1 => C, A2 => n30, ZN => n29);
   U12 : AOI22_X1 port map( A1 => n28, A2 => n6, B1 => D, B2 => n27, ZN => n31)
                           ;
   U13 : NOR3_X1 port map( A1 => S(0), A2 => n3, A3 => n2, ZN => n30);
   U14 : NAND4_X1 port map( A1 => n26, A2 => n25, A3 => n24, A4 => n23, ZN => 
                           n28);
   U15 : NAND4_X1 port map( A1 => E, A2 => n3, A3 => n1, A4 => n2, ZN => n26);
   U16 : NOR2_X1 port map( A1 => n2, A2 => S(0), ZN => n22);
   U17 : INV_X1 port map( A => S(0), ZN => n1);
   U18 : INV_X1 port map( A => S(1), ZN => n2);
   U19 : INV_X1 port map( A => n4, ZN => n3);
   U22 : INV_X1 port map( A => S(2), ZN => n4);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX81_12 is

   port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
         downto 0);  Y : out std_logic);

end MUX81_12;

architecture SYN_BEHAVIORAL_1 of MUX81_12 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n21, n22, n23, n24, n25, n26, n27, n28, n29, 
      n30, n31, n32, n33, n34 : std_logic;

begin
   
   U20 : NAND3_X1 port map( A1 => S(1), A2 => n6, A3 => H, ZN => n22);
   U21 : NAND3_X1 port map( A1 => S(0), A2 => n2, A3 => F, ZN => n24);
   U1 : INV_X1 port map( A => n26, ZN => n5);
   U2 : NAND2_X1 port map( A1 => G, A2 => n21, ZN => n23);
   U3 : NOR2_X1 port map( A1 => n1, A2 => S(2), ZN => n26);
   U4 : NAND4_X1 port map( A1 => A, A2 => n1, A3 => n2, A4 => n3, ZN => n33);
   U5 : INV_X1 port map( A => n21, ZN => n6);
   U6 : AOI22_X1 port map( A1 => n32, A2 => n4, B1 => B, B2 => n31, ZN => n34);
   U7 : INV_X1 port map( A => n31, ZN => n4);
   U8 : NOR3_X1 port map( A1 => S(1), A2 => S(2), A3 => n1, ZN => n31);
   U9 : OAI21_X1 port map( B1 => n30, B2 => n29, A => n28, ZN => n32);
   U10 : NAND2_X1 port map( A1 => C, A2 => n29, ZN => n28);
   U11 : AOI22_X1 port map( A1 => n27, A2 => n5, B1 => D, B2 => n26, ZN => n30)
                           ;
   U12 : NOR3_X1 port map( A1 => S(0), A2 => S(2), A3 => n2, ZN => n29);
   U13 : NAND4_X1 port map( A1 => n25, A2 => n24, A3 => n23, A4 => n22, ZN => 
                           n27);
   U14 : NAND4_X1 port map( A1 => E, A2 => S(2), A3 => n1, A4 => n2, ZN => n25)
                           ;
   U15 : NOR2_X1 port map( A1 => n2, A2 => S(0), ZN => n21);
   U16 : NAND2_X1 port map( A1 => n34, A2 => n33, ZN => Y);
   U17 : INV_X1 port map( A => S(0), ZN => n1);
   U18 : INV_X1 port map( A => S(1), ZN => n2);
   U19 : INV_X1 port map( A => S(2), ZN => n3);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX81_11 is

   port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
         downto 0);  Y : out std_logic);

end MUX81_11;

architecture SYN_BEHAVIORAL_1 of MUX81_11 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n21, n22, n23, n24, n25, n26, n27, n28, n29, 
      n30, n31, n32, n33, n34 : std_logic;

begin
   
   U20 : NAND3_X1 port map( A1 => S(1), A2 => n6, A3 => H, ZN => n22);
   U21 : NAND3_X1 port map( A1 => S(0), A2 => n2, A3 => F, ZN => n24);
   U1 : INV_X1 port map( A => n26, ZN => n5);
   U2 : NAND2_X1 port map( A1 => G, A2 => n21, ZN => n23);
   U3 : NOR2_X1 port map( A1 => n1, A2 => S(2), ZN => n26);
   U4 : NAND4_X1 port map( A1 => A, A2 => n1, A3 => n2, A4 => n3, ZN => n33);
   U5 : INV_X1 port map( A => n21, ZN => n6);
   U6 : NAND2_X1 port map( A1 => n34, A2 => n33, ZN => Y);
   U7 : AOI22_X1 port map( A1 => n32, A2 => n4, B1 => B, B2 => n31, ZN => n34);
   U8 : INV_X1 port map( A => n31, ZN => n4);
   U9 : NOR3_X1 port map( A1 => S(1), A2 => S(2), A3 => n1, ZN => n31);
   U10 : OAI21_X1 port map( B1 => n30, B2 => n29, A => n28, ZN => n32);
   U11 : NAND2_X1 port map( A1 => C, A2 => n29, ZN => n28);
   U12 : AOI22_X1 port map( A1 => n27, A2 => n5, B1 => D, B2 => n26, ZN => n30)
                           ;
   U13 : NOR3_X1 port map( A1 => S(0), A2 => S(2), A3 => n2, ZN => n29);
   U14 : NAND4_X1 port map( A1 => n25, A2 => n24, A3 => n23, A4 => n22, ZN => 
                           n27);
   U15 : NAND4_X1 port map( A1 => E, A2 => S(2), A3 => n1, A4 => n2, ZN => n25)
                           ;
   U16 : NOR2_X1 port map( A1 => n2, A2 => S(0), ZN => n21);
   U17 : INV_X1 port map( A => S(0), ZN => n1);
   U18 : INV_X1 port map( A => S(1), ZN => n2);
   U19 : INV_X1 port map( A => S(2), ZN => n3);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX81_10 is

   port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
         downto 0);  Y : out std_logic);

end MUX81_10;

architecture SYN_BEHAVIORAL_1 of MUX81_10 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n21, n22, n23, n24, n25, n26, n27, n28, n29, 
      n30, n31, n32, n33, n34 : std_logic;

begin
   
   U20 : NAND3_X1 port map( A1 => S(1), A2 => n6, A3 => H, ZN => n22);
   U21 : NAND3_X1 port map( A1 => S(0), A2 => n2, A3 => F, ZN => n24);
   U1 : INV_X1 port map( A => n26, ZN => n5);
   U2 : NAND2_X1 port map( A1 => G, A2 => n21, ZN => n23);
   U3 : NOR2_X1 port map( A1 => n1, A2 => S(2), ZN => n26);
   U4 : NAND4_X1 port map( A1 => A, A2 => n1, A3 => n2, A4 => n3, ZN => n33);
   U5 : INV_X1 port map( A => n21, ZN => n6);
   U6 : NAND2_X1 port map( A1 => n34, A2 => n33, ZN => Y);
   U7 : AOI22_X1 port map( A1 => n32, A2 => n4, B1 => B, B2 => n31, ZN => n34);
   U8 : INV_X1 port map( A => n31, ZN => n4);
   U9 : NOR3_X1 port map( A1 => S(1), A2 => S(2), A3 => n1, ZN => n31);
   U10 : OAI21_X1 port map( B1 => n30, B2 => n29, A => n28, ZN => n32);
   U11 : NAND2_X1 port map( A1 => C, A2 => n29, ZN => n28);
   U12 : AOI22_X1 port map( A1 => n27, A2 => n5, B1 => D, B2 => n26, ZN => n30)
                           ;
   U13 : NOR3_X1 port map( A1 => S(0), A2 => S(2), A3 => n2, ZN => n29);
   U14 : NAND4_X1 port map( A1 => n25, A2 => n24, A3 => n23, A4 => n22, ZN => 
                           n27);
   U15 : NAND4_X1 port map( A1 => E, A2 => S(2), A3 => n1, A4 => n2, ZN => n25)
                           ;
   U16 : NOR2_X1 port map( A1 => n2, A2 => S(0), ZN => n21);
   U17 : INV_X1 port map( A => S(0), ZN => n1);
   U18 : INV_X1 port map( A => S(1), ZN => n2);
   U19 : INV_X1 port map( A => S(2), ZN => n3);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX81_9 is

   port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
         downto 0);  Y : out std_logic);

end MUX81_9;

architecture SYN_BEHAVIORAL_1 of MUX81_9 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n21, n22, n23, n24, n25, n26, n27, n28, n29, 
      n30, n31, n32, n33, n34, n35 : std_logic;

begin
   
   U20 : NAND3_X1 port map( A1 => S(1), A2 => n21, A3 => H, ZN => n23);
   U21 : NAND3_X1 port map( A1 => S(0), A2 => n2, A3 => F, ZN => n25);
   U1 : INV_X1 port map( A => n27, ZN => n6);
   U2 : NOR2_X1 port map( A1 => n1, A2 => n3, ZN => n27);
   U3 : NAND4_X1 port map( A1 => A, A2 => n1, A3 => n2, A4 => n4, ZN => n34);
   U4 : INV_X1 port map( A => n22, ZN => n21);
   U5 : AOI22_X1 port map( A1 => n33, A2 => n5, B1 => B, B2 => n32, ZN => n35);
   U6 : INV_X1 port map( A => n32, ZN => n5);
   U7 : NOR3_X1 port map( A1 => S(1), A2 => n3, A3 => n1, ZN => n32);
   U8 : OAI21_X1 port map( B1 => n31, B2 => n30, A => n29, ZN => n33);
   U9 : NAND2_X1 port map( A1 => C, A2 => n30, ZN => n29);
   U10 : AOI22_X1 port map( A1 => n28, A2 => n6, B1 => D, B2 => n27, ZN => n31)
                           ;
   U11 : NOR3_X1 port map( A1 => S(0), A2 => n3, A3 => n2, ZN => n30);
   U12 : NAND4_X1 port map( A1 => n26, A2 => n25, A3 => n24, A4 => n23, ZN => 
                           n28);
   U13 : NAND4_X1 port map( A1 => E, A2 => n3, A3 => n1, A4 => n2, ZN => n26);
   U14 : NAND2_X1 port map( A1 => G, A2 => n22, ZN => n24);
   U15 : NAND2_X1 port map( A1 => n35, A2 => n34, ZN => Y);
   U16 : NOR2_X1 port map( A1 => n2, A2 => S(0), ZN => n22);
   U17 : INV_X1 port map( A => S(0), ZN => n1);
   U18 : INV_X1 port map( A => S(1), ZN => n2);
   U19 : INV_X1 port map( A => n4, ZN => n3);
   U22 : INV_X1 port map( A => S(2), ZN => n4);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX81_8 is

   port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
         downto 0);  Y : out std_logic);

end MUX81_8;

architecture SYN_BEHAVIORAL_1 of MUX81_8 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n21, n22, n23, n24, n25, n26, n27, n28, n29, 
      n30, n31, n32, n33, n34, n35 : std_logic;

begin
   
   U20 : NAND3_X1 port map( A1 => S(1), A2 => n21, A3 => H, ZN => n23);
   U21 : NAND3_X1 port map( A1 => S(0), A2 => n2, A3 => F, ZN => n25);
   U1 : INV_X1 port map( A => n27, ZN => n6);
   U2 : NOR2_X1 port map( A1 => n1, A2 => n3, ZN => n27);
   U3 : NAND4_X1 port map( A1 => A, A2 => n1, A3 => n2, A4 => n4, ZN => n34);
   U4 : INV_X1 port map( A => n22, ZN => n21);
   U5 : AOI22_X1 port map( A1 => n33, A2 => n5, B1 => B, B2 => n32, ZN => n35);
   U6 : INV_X1 port map( A => n32, ZN => n5);
   U7 : NOR3_X1 port map( A1 => S(1), A2 => n3, A3 => n1, ZN => n32);
   U8 : OAI21_X1 port map( B1 => n31, B2 => n30, A => n29, ZN => n33);
   U9 : NAND2_X1 port map( A1 => C, A2 => n30, ZN => n29);
   U10 : AOI22_X1 port map( A1 => n28, A2 => n6, B1 => D, B2 => n27, ZN => n31)
                           ;
   U11 : NOR3_X1 port map( A1 => S(0), A2 => n3, A3 => n2, ZN => n30);
   U12 : NAND4_X1 port map( A1 => n26, A2 => n25, A3 => n24, A4 => n23, ZN => 
                           n28);
   U13 : NAND4_X1 port map( A1 => E, A2 => n3, A3 => n1, A4 => n2, ZN => n26);
   U14 : NAND2_X1 port map( A1 => G, A2 => n22, ZN => n24);
   U15 : NOR2_X1 port map( A1 => n2, A2 => S(0), ZN => n22);
   U16 : NAND2_X1 port map( A1 => n35, A2 => n34, ZN => Y);
   U17 : INV_X1 port map( A => S(0), ZN => n1);
   U18 : INV_X1 port map( A => S(1), ZN => n2);
   U19 : INV_X1 port map( A => n4, ZN => n3);
   U22 : INV_X1 port map( A => S(2), ZN => n4);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX81_7 is

   port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
         downto 0);  Y : out std_logic);

end MUX81_7;

architecture SYN_BEHAVIORAL_1 of MUX81_7 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n21, n22, n23, n24, n25, n26, n27, n28, n29, 
      n30, n31, n32, n33, n34, n35 : std_logic;

begin
   
   U20 : NAND3_X1 port map( A1 => S(1), A2 => n21, A3 => H, ZN => n23);
   U21 : NAND3_X1 port map( A1 => S(0), A2 => n2, A3 => F, ZN => n25);
   U1 : INV_X1 port map( A => n27, ZN => n6);
   U2 : NAND2_X1 port map( A1 => G, A2 => n22, ZN => n24);
   U3 : NOR2_X1 port map( A1 => n1, A2 => n3, ZN => n27);
   U4 : NAND4_X1 port map( A1 => A, A2 => n1, A3 => n2, A4 => n4, ZN => n34);
   U5 : INV_X1 port map( A => n22, ZN => n21);
   U6 : AOI22_X1 port map( A1 => n33, A2 => n5, B1 => B, B2 => n32, ZN => n35);
   U7 : INV_X1 port map( A => n32, ZN => n5);
   U8 : NOR3_X1 port map( A1 => S(1), A2 => n3, A3 => n1, ZN => n32);
   U9 : OAI21_X1 port map( B1 => n31, B2 => n30, A => n29, ZN => n33);
   U10 : NAND2_X1 port map( A1 => C, A2 => n30, ZN => n29);
   U11 : AOI22_X1 port map( A1 => n28, A2 => n6, B1 => D, B2 => n27, ZN => n31)
                           ;
   U12 : NOR3_X1 port map( A1 => S(0), A2 => n3, A3 => n2, ZN => n30);
   U13 : NAND4_X1 port map( A1 => n26, A2 => n25, A3 => n24, A4 => n23, ZN => 
                           n28);
   U14 : NAND4_X1 port map( A1 => E, A2 => n3, A3 => n1, A4 => n2, ZN => n26);
   U15 : NAND2_X1 port map( A1 => n35, A2 => n34, ZN => Y);
   U16 : NOR2_X1 port map( A1 => n2, A2 => S(0), ZN => n22);
   U17 : INV_X1 port map( A => S(0), ZN => n1);
   U18 : INV_X1 port map( A => S(1), ZN => n2);
   U19 : INV_X1 port map( A => n4, ZN => n3);
   U22 : INV_X1 port map( A => S(2), ZN => n4);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX81_6 is

   port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
         downto 0);  Y : out std_logic);

end MUX81_6;

architecture SYN_BEHAVIORAL_1 of MUX81_6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n21, n22, n23, n24, n25, n26, n27, n28, n29, 
      n30, n31, n32, n33, n34, n35 : std_logic;

begin
   
   U20 : NAND3_X1 port map( A1 => S(1), A2 => n21, A3 => H, ZN => n23);
   U21 : NAND3_X1 port map( A1 => S(0), A2 => n2, A3 => F, ZN => n25);
   U1 : INV_X1 port map( A => n27, ZN => n6);
   U2 : NOR2_X1 port map( A1 => n1, A2 => n3, ZN => n27);
   U3 : NAND4_X1 port map( A1 => A, A2 => n1, A3 => n2, A4 => n4, ZN => n34);
   U4 : INV_X1 port map( A => n22, ZN => n21);
   U5 : AOI22_X1 port map( A1 => n33, A2 => n5, B1 => B, B2 => n32, ZN => n35);
   U6 : INV_X1 port map( A => n32, ZN => n5);
   U7 : NOR3_X1 port map( A1 => S(1), A2 => n3, A3 => n1, ZN => n32);
   U8 : OAI21_X1 port map( B1 => n31, B2 => n30, A => n29, ZN => n33);
   U9 : NAND2_X1 port map( A1 => C, A2 => n30, ZN => n29);
   U10 : AOI22_X1 port map( A1 => n28, A2 => n6, B1 => D, B2 => n27, ZN => n31)
                           ;
   U11 : NOR3_X1 port map( A1 => S(0), A2 => n3, A3 => n2, ZN => n30);
   U12 : NAND4_X1 port map( A1 => n26, A2 => n25, A3 => n24, A4 => n23, ZN => 
                           n28);
   U13 : NAND4_X1 port map( A1 => E, A2 => n3, A3 => n1, A4 => n2, ZN => n26);
   U14 : NAND2_X1 port map( A1 => G, A2 => n22, ZN => n24);
   U15 : NAND2_X1 port map( A1 => n35, A2 => n34, ZN => Y);
   U16 : NOR2_X1 port map( A1 => n2, A2 => S(0), ZN => n22);
   U17 : INV_X1 port map( A => S(0), ZN => n1);
   U18 : INV_X1 port map( A => S(1), ZN => n2);
   U19 : INV_X1 port map( A => n4, ZN => n3);
   U22 : INV_X1 port map( A => S(2), ZN => n4);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX81_5 is

   port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
         downto 0);  Y : out std_logic);

end MUX81_5;

architecture SYN_BEHAVIORAL_1 of MUX81_5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n21, n22, n23, n24, n25, n26, n27, n28, n29, 
      n30, n31, n32, n33, n34, n35 : std_logic;

begin
   
   U20 : NAND3_X1 port map( A1 => S(1), A2 => n21, A3 => H, ZN => n23);
   U21 : NAND3_X1 port map( A1 => S(0), A2 => n2, A3 => F, ZN => n25);
   U1 : INV_X1 port map( A => n27, ZN => n6);
   U2 : NOR2_X1 port map( A1 => n1, A2 => n3, ZN => n27);
   U3 : NAND4_X1 port map( A1 => A, A2 => n1, A3 => n2, A4 => n4, ZN => n34);
   U4 : INV_X1 port map( A => n22, ZN => n21);
   U5 : AOI22_X1 port map( A1 => n33, A2 => n5, B1 => B, B2 => n32, ZN => n35);
   U6 : INV_X1 port map( A => n32, ZN => n5);
   U7 : NOR3_X1 port map( A1 => S(1), A2 => n3, A3 => n1, ZN => n32);
   U8 : OAI21_X1 port map( B1 => n31, B2 => n30, A => n29, ZN => n33);
   U9 : NAND2_X1 port map( A1 => C, A2 => n30, ZN => n29);
   U10 : AOI22_X1 port map( A1 => n28, A2 => n6, B1 => D, B2 => n27, ZN => n31)
                           ;
   U11 : NOR3_X1 port map( A1 => S(0), A2 => n3, A3 => n2, ZN => n30);
   U12 : NAND4_X1 port map( A1 => n26, A2 => n25, A3 => n24, A4 => n23, ZN => 
                           n28);
   U13 : NAND4_X1 port map( A1 => E, A2 => n3, A3 => n1, A4 => n2, ZN => n26);
   U14 : NAND2_X1 port map( A1 => G, A2 => n22, ZN => n24);
   U15 : NAND2_X1 port map( A1 => n35, A2 => n34, ZN => Y);
   U16 : NOR2_X1 port map( A1 => n2, A2 => S(0), ZN => n22);
   U17 : INV_X1 port map( A => S(0), ZN => n1);
   U18 : INV_X1 port map( A => S(1), ZN => n2);
   U19 : INV_X1 port map( A => n4, ZN => n3);
   U22 : INV_X1 port map( A => S(2), ZN => n4);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX81_4 is

   port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
         downto 0);  Y : out std_logic);

end MUX81_4;

architecture SYN_BEHAVIORAL_1 of MUX81_4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n21, n22, n23, n24, n25, n26, n27, n28, n29, 
      n30, n31, n32, n33, n34, n35 : std_logic;

begin
   
   U20 : NAND3_X1 port map( A1 => S(1), A2 => n21, A3 => H, ZN => n23);
   U21 : NAND3_X1 port map( A1 => S(0), A2 => n2, A3 => F, ZN => n25);
   U1 : INV_X1 port map( A => n27, ZN => n6);
   U2 : NOR2_X1 port map( A1 => n1, A2 => n3, ZN => n27);
   U3 : NAND4_X1 port map( A1 => A, A2 => n1, A3 => n2, A4 => n4, ZN => n34);
   U4 : INV_X1 port map( A => n22, ZN => n21);
   U5 : AOI22_X1 port map( A1 => n33, A2 => n5, B1 => B, B2 => n32, ZN => n35);
   U6 : INV_X1 port map( A => n32, ZN => n5);
   U7 : NOR3_X1 port map( A1 => S(1), A2 => n3, A3 => n1, ZN => n32);
   U8 : OAI21_X1 port map( B1 => n31, B2 => n30, A => n29, ZN => n33);
   U9 : NAND2_X1 port map( A1 => C, A2 => n30, ZN => n29);
   U10 : AOI22_X1 port map( A1 => n28, A2 => n6, B1 => D, B2 => n27, ZN => n31)
                           ;
   U11 : NOR3_X1 port map( A1 => S(0), A2 => n3, A3 => n2, ZN => n30);
   U12 : NAND4_X1 port map( A1 => n26, A2 => n25, A3 => n24, A4 => n23, ZN => 
                           n28);
   U13 : NAND4_X1 port map( A1 => E, A2 => n3, A3 => n1, A4 => n2, ZN => n26);
   U14 : NAND2_X1 port map( A1 => G, A2 => n22, ZN => n24);
   U15 : NOR2_X1 port map( A1 => n2, A2 => S(0), ZN => n22);
   U16 : NAND2_X1 port map( A1 => n35, A2 => n34, ZN => Y);
   U17 : INV_X1 port map( A => S(0), ZN => n1);
   U18 : INV_X1 port map( A => S(1), ZN => n2);
   U19 : INV_X1 port map( A => n4, ZN => n3);
   U22 : INV_X1 port map( A => S(2), ZN => n4);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX81_3 is

   port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
         downto 0);  Y : out std_logic);

end MUX81_3;

architecture SYN_BEHAVIORAL_1 of MUX81_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n21, n22, n23, n24, n25, n26, n27, n28, n29, 
      n30, n31, n32, n33, n34, n35 : std_logic;

begin
   
   U20 : NAND3_X1 port map( A1 => S(1), A2 => n21, A3 => H, ZN => n23);
   U21 : NAND3_X1 port map( A1 => S(0), A2 => n2, A3 => F, ZN => n25);
   U1 : INV_X1 port map( A => n27, ZN => n6);
   U2 : NOR2_X1 port map( A1 => n1, A2 => n3, ZN => n27);
   U3 : NAND4_X1 port map( A1 => A, A2 => n1, A3 => n2, A4 => n4, ZN => n34);
   U4 : INV_X1 port map( A => n22, ZN => n21);
   U5 : AOI22_X1 port map( A1 => n33, A2 => n5, B1 => B, B2 => n32, ZN => n35);
   U6 : INV_X1 port map( A => n32, ZN => n5);
   U7 : NOR3_X1 port map( A1 => S(1), A2 => n3, A3 => n1, ZN => n32);
   U8 : OAI21_X1 port map( B1 => n31, B2 => n30, A => n29, ZN => n33);
   U9 : NAND2_X1 port map( A1 => C, A2 => n30, ZN => n29);
   U10 : AOI22_X1 port map( A1 => n28, A2 => n6, B1 => D, B2 => n27, ZN => n31)
                           ;
   U11 : NOR3_X1 port map( A1 => S(0), A2 => n3, A3 => n2, ZN => n30);
   U12 : NAND4_X1 port map( A1 => n26, A2 => n25, A3 => n24, A4 => n23, ZN => 
                           n28);
   U13 : NAND4_X1 port map( A1 => E, A2 => n3, A3 => n1, A4 => n2, ZN => n26);
   U14 : NAND2_X1 port map( A1 => G, A2 => n22, ZN => n24);
   U15 : NAND2_X1 port map( A1 => n35, A2 => n34, ZN => Y);
   U16 : NOR2_X1 port map( A1 => n2, A2 => S(0), ZN => n22);
   U17 : INV_X1 port map( A => S(0), ZN => n1);
   U18 : INV_X1 port map( A => S(1), ZN => n2);
   U19 : INV_X1 port map( A => n4, ZN => n3);
   U22 : INV_X1 port map( A => S(2), ZN => n4);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX81_2 is

   port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
         downto 0);  Y : out std_logic);

end MUX81_2;

architecture SYN_BEHAVIORAL_1 of MUX81_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n21, n22, n23, n24, n25, n26, n27, n28, n29, 
      n30, n31, n32, n33, n34 : std_logic;

begin
   
   U20 : NAND3_X1 port map( A1 => S(1), A2 => n6, A3 => H, ZN => n22);
   U21 : NAND3_X1 port map( A1 => S(0), A2 => n2, A3 => F, ZN => n24);
   U1 : INV_X1 port map( A => n26, ZN => n5);
   U2 : NOR2_X1 port map( A1 => n1, A2 => S(2), ZN => n26);
   U3 : NAND4_X1 port map( A1 => A, A2 => n1, A3 => n2, A4 => n3, ZN => n33);
   U4 : INV_X1 port map( A => n21, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n32, A2 => n4, B1 => B, B2 => n31, ZN => n34);
   U6 : INV_X1 port map( A => n31, ZN => n4);
   U7 : NOR3_X1 port map( A1 => S(1), A2 => S(2), A3 => n1, ZN => n31);
   U8 : OAI21_X1 port map( B1 => n30, B2 => n29, A => n28, ZN => n32);
   U9 : NAND2_X1 port map( A1 => C, A2 => n29, ZN => n28);
   U10 : AOI22_X1 port map( A1 => n27, A2 => n5, B1 => D, B2 => n26, ZN => n30)
                           ;
   U11 : NOR3_X1 port map( A1 => S(0), A2 => S(2), A3 => n2, ZN => n29);
   U12 : NAND4_X1 port map( A1 => n25, A2 => n24, A3 => n23, A4 => n22, ZN => 
                           n27);
   U13 : NAND4_X1 port map( A1 => E, A2 => S(2), A3 => n1, A4 => n2, ZN => n25)
                           ;
   U14 : NAND2_X1 port map( A1 => G, A2 => n21, ZN => n23);
   U15 : NAND2_X1 port map( A1 => n34, A2 => n33, ZN => Y);
   U16 : NOR2_X1 port map( A1 => n2, A2 => S(0), ZN => n21);
   U17 : INV_X1 port map( A => S(0), ZN => n1);
   U18 : INV_X1 port map( A => S(1), ZN => n2);
   U19 : INV_X1 port map( A => S(2), ZN => n3);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX81_1 is

   port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
         downto 0);  Y : out std_logic);

end MUX81_1;

architecture SYN_BEHAVIORAL_1 of MUX81_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n21, n22, n23, n24, n25, n26, n27, n28, n29, 
      n30, n31, n32, n33, n34 : std_logic;

begin
   
   U20 : NAND3_X1 port map( A1 => S(1), A2 => n6, A3 => H, ZN => n22);
   U21 : NAND3_X1 port map( A1 => S(0), A2 => n2, A3 => F, ZN => n24);
   U1 : INV_X1 port map( A => n26, ZN => n5);
   U2 : NOR2_X1 port map( A1 => n1, A2 => S(2), ZN => n26);
   U3 : NAND4_X1 port map( A1 => A, A2 => n1, A3 => n2, A4 => n3, ZN => n33);
   U4 : INV_X1 port map( A => n21, ZN => n6);
   U5 : AOI22_X1 port map( A1 => n32, A2 => n4, B1 => B, B2 => n31, ZN => n34);
   U6 : INV_X1 port map( A => n31, ZN => n4);
   U7 : NOR3_X1 port map( A1 => S(1), A2 => S(2), A3 => n1, ZN => n31);
   U8 : OAI21_X1 port map( B1 => n30, B2 => n29, A => n28, ZN => n32);
   U9 : NAND2_X1 port map( A1 => C, A2 => n29, ZN => n28);
   U10 : AOI22_X1 port map( A1 => n27, A2 => n5, B1 => D, B2 => n26, ZN => n30)
                           ;
   U11 : NOR3_X1 port map( A1 => S(0), A2 => S(2), A3 => n2, ZN => n29);
   U12 : NAND4_X1 port map( A1 => n25, A2 => n24, A3 => n23, A4 => n22, ZN => 
                           n27);
   U13 : NAND4_X1 port map( A1 => E, A2 => S(2), A3 => n1, A4 => n2, ZN => n25)
                           ;
   U14 : NAND2_X1 port map( A1 => G, A2 => n21, ZN => n23);
   U15 : NAND2_X1 port map( A1 => n34, A2 => n33, ZN => Y);
   U16 : NOR2_X1 port map( A1 => n2, A2 => S(0), ZN => n21);
   U17 : INV_X1 port map( A => S(0), ZN => n1);
   U18 : INV_X1 port map( A => S(1), ZN => n2);
   U19 : INV_X1 port map( A => S(2), ZN => n3);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_GENERIC_NBIT8_3 is

   port( A, B, C, D : in std_logic_vector (7 downto 0);  SEL : in 
         std_logic_vector (1 downto 0);  Y : out std_logic_vector (7 downto 0)
         );

end MUX41_GENERIC_NBIT8_3;

architecture SYN_structural of MUX41_GENERIC_NBIT8_3 is

   component MUX41_17
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_18
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_19
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_20
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_21
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_22
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_23
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_24
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX41_24 port map( A => A(0), B => B(0), C => C(0), D => D(0), 
                           S(1) => SEL(1), S(0) => SEL(0), Y => Y(0));
   MUXES_1 : MUX41_23 port map( A => A(1), B => B(1), C => C(1), D => D(1), 
                           S(1) => SEL(1), S(0) => SEL(0), Y => Y(1));
   MUXES_2 : MUX41_22 port map( A => A(2), B => B(2), C => C(2), D => D(2), 
                           S(1) => SEL(1), S(0) => SEL(0), Y => Y(2));
   MUXES_3 : MUX41_21 port map( A => A(3), B => B(3), C => C(3), D => D(3), 
                           S(1) => SEL(1), S(0) => SEL(0), Y => Y(3));
   MUXES_4 : MUX41_20 port map( A => A(4), B => B(4), C => C(4), D => D(4), 
                           S(1) => SEL(1), S(0) => SEL(0), Y => Y(4));
   MUXES_5 : MUX41_19 port map( A => A(5), B => B(5), C => C(5), D => D(5), 
                           S(1) => SEL(1), S(0) => SEL(0), Y => Y(5));
   MUXES_6 : MUX41_18 port map( A => A(6), B => B(6), C => C(6), D => D(6), 
                           S(1) => SEL(1), S(0) => SEL(0), Y => Y(6));
   MUXES_7 : MUX41_17 port map( A => A(7), B => B(7), C => C(7), D => D(7), 
                           S(1) => SEL(1), S(0) => SEL(0), Y => Y(7));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_GENERIC_NBIT8_2 is

   port( A, B, C, D : in std_logic_vector (7 downto 0);  SEL : in 
         std_logic_vector (1 downto 0);  Y : out std_logic_vector (7 downto 0)
         );

end MUX41_GENERIC_NBIT8_2;

architecture SYN_structural of MUX41_GENERIC_NBIT8_2 is

   component MUX41_9
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_10
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_11
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_12
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_13
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_14
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_15
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_16
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX41_16 port map( A => A(0), B => B(0), C => C(0), D => D(0), 
                           S(1) => SEL(1), S(0) => SEL(0), Y => Y(0));
   MUXES_1 : MUX41_15 port map( A => A(1), B => B(1), C => C(1), D => D(1), 
                           S(1) => SEL(1), S(0) => SEL(0), Y => Y(1));
   MUXES_2 : MUX41_14 port map( A => A(2), B => B(2), C => C(2), D => D(2), 
                           S(1) => SEL(1), S(0) => SEL(0), Y => Y(2));
   MUXES_3 : MUX41_13 port map( A => A(3), B => B(3), C => C(3), D => D(3), 
                           S(1) => SEL(1), S(0) => SEL(0), Y => Y(3));
   MUXES_4 : MUX41_12 port map( A => A(4), B => B(4), C => C(4), D => D(4), 
                           S(1) => SEL(1), S(0) => SEL(0), Y => Y(4));
   MUXES_5 : MUX41_11 port map( A => A(5), B => B(5), C => C(5), D => D(5), 
                           S(1) => SEL(1), S(0) => SEL(0), Y => Y(5));
   MUXES_6 : MUX41_10 port map( A => A(6), B => B(6), C => C(6), D => D(6), 
                           S(1) => SEL(1), S(0) => SEL(0), Y => Y(6));
   MUXES_7 : MUX41_9 port map( A => A(7), B => B(7), C => C(7), D => D(7), S(1)
                           => SEL(1), S(0) => SEL(0), Y => Y(7));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_GENERIC_NBIT8_1 is

   port( A, B, C, D : in std_logic_vector (7 downto 0);  SEL : in 
         std_logic_vector (1 downto 0);  Y : out std_logic_vector (7 downto 0)
         );

end MUX41_GENERIC_NBIT8_1;

architecture SYN_structural of MUX41_GENERIC_NBIT8_1 is

   component MUX41_1
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_2
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_3
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_4
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_5
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_6
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_7
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_8
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX41_8 port map( A => A(0), B => B(0), C => C(0), D => D(0), S(1)
                           => SEL(1), S(0) => SEL(0), Y => Y(0));
   MUXES_1 : MUX41_7 port map( A => A(1), B => B(1), C => C(1), D => D(1), S(1)
                           => SEL(1), S(0) => SEL(0), Y => Y(1));
   MUXES_2 : MUX41_6 port map( A => A(2), B => B(2), C => C(2), D => D(2), S(1)
                           => SEL(1), S(0) => SEL(0), Y => Y(2));
   MUXES_3 : MUX41_5 port map( A => A(3), B => B(3), C => C(3), D => D(3), S(1)
                           => SEL(1), S(0) => SEL(0), Y => Y(3));
   MUXES_4 : MUX41_4 port map( A => A(4), B => B(4), C => C(4), D => D(4), S(1)
                           => SEL(1), S(0) => SEL(0), Y => Y(4));
   MUXES_5 : MUX41_3 port map( A => A(5), B => B(5), C => C(5), D => D(5), S(1)
                           => SEL(1), S(0) => SEL(0), Y => Y(5));
   MUXES_6 : MUX41_2 port map( A => A(6), B => B(6), C => C(6), D => D(6), S(1)
                           => SEL(1), S(0) => SEL(0), Y => Y(6));
   MUXES_7 : MUX41_1 port map( A => A(7), B => B(7), C => C(7), D => D(7), S(1)
                           => SEL(1), S(0) => SEL(0), Y => Y(7));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT8_16 is

   port( A, B : in std_logic_vector (7 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (7 downto 0));

end MUX21_GENERIC_NBIT8_16;

architecture SYN_structural of MUX21_GENERIC_NBIT8_16 is

   component MUX21_345
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_346
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_347
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_348
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_349
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_350
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_351
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_352
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_352 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_351 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_350 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_349 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));
   MUXES_4 : MUX21_348 port map( A => A(4), B => B(4), S => SEL, Y => Y(4));
   MUXES_5 : MUX21_347 port map( A => A(5), B => B(5), S => SEL, Y => Y(5));
   MUXES_6 : MUX21_346 port map( A => A(6), B => B(6), S => SEL, Y => Y(6));
   MUXES_7 : MUX21_345 port map( A => A(7), B => B(7), S => SEL, Y => Y(7));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT8_15 is

   port( A, B : in std_logic_vector (7 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (7 downto 0));

end MUX21_GENERIC_NBIT8_15;

architecture SYN_structural of MUX21_GENERIC_NBIT8_15 is

   component MUX21_337
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_338
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_339
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_340
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_341
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_342
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_343
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_344
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_344 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_343 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_342 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_341 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));
   MUXES_4 : MUX21_340 port map( A => A(4), B => B(4), S => SEL, Y => Y(4));
   MUXES_5 : MUX21_339 port map( A => A(5), B => B(5), S => SEL, Y => Y(5));
   MUXES_6 : MUX21_338 port map( A => A(6), B => B(6), S => SEL, Y => Y(6));
   MUXES_7 : MUX21_337 port map( A => A(7), B => B(7), S => SEL, Y => Y(7));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT8_14 is

   port( A, B : in std_logic_vector (7 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (7 downto 0));

end MUX21_GENERIC_NBIT8_14;

architecture SYN_structural of MUX21_GENERIC_NBIT8_14 is

   component MUX21_329
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_330
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_331
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_332
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_333
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_334
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_335
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_336
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_336 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_335 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_334 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_333 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));
   MUXES_4 : MUX21_332 port map( A => A(4), B => B(4), S => SEL, Y => Y(4));
   MUXES_5 : MUX21_331 port map( A => A(5), B => B(5), S => SEL, Y => Y(5));
   MUXES_6 : MUX21_330 port map( A => A(6), B => B(6), S => SEL, Y => Y(6));
   MUXES_7 : MUX21_329 port map( A => A(7), B => B(7), S => SEL, Y => Y(7));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT8_13 is

   port( A, B : in std_logic_vector (7 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (7 downto 0));

end MUX21_GENERIC_NBIT8_13;

architecture SYN_structural of MUX21_GENERIC_NBIT8_13 is

   component MUX21_321
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_322
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_323
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_324
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_325
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_326
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_327
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_328
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_328 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_327 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_326 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_325 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));
   MUXES_4 : MUX21_324 port map( A => A(4), B => B(4), S => SEL, Y => Y(4));
   MUXES_5 : MUX21_323 port map( A => A(5), B => B(5), S => SEL, Y => Y(5));
   MUXES_6 : MUX21_322 port map( A => A(6), B => B(6), S => SEL, Y => Y(6));
   MUXES_7 : MUX21_321 port map( A => A(7), B => B(7), S => SEL, Y => Y(7));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT8_12 is

   port( A, B : in std_logic_vector (7 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (7 downto 0));

end MUX21_GENERIC_NBIT8_12;

architecture SYN_structural of MUX21_GENERIC_NBIT8_12 is

   component MUX21_313
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_314
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_315
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_316
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_317
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_318
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_319
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_320
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_320 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_319 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_318 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_317 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));
   MUXES_4 : MUX21_316 port map( A => A(4), B => B(4), S => SEL, Y => Y(4));
   MUXES_5 : MUX21_315 port map( A => A(5), B => B(5), S => SEL, Y => Y(5));
   MUXES_6 : MUX21_314 port map( A => A(6), B => B(6), S => SEL, Y => Y(6));
   MUXES_7 : MUX21_313 port map( A => A(7), B => B(7), S => SEL, Y => Y(7));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT8_11 is

   port( A, B : in std_logic_vector (7 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (7 downto 0));

end MUX21_GENERIC_NBIT8_11;

architecture SYN_structural of MUX21_GENERIC_NBIT8_11 is

   component MUX21_305
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_306
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_307
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_308
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_309
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_310
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_311
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_312
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_312 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_311 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_310 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_309 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));
   MUXES_4 : MUX21_308 port map( A => A(4), B => B(4), S => SEL, Y => Y(4));
   MUXES_5 : MUX21_307 port map( A => A(5), B => B(5), S => SEL, Y => Y(5));
   MUXES_6 : MUX21_306 port map( A => A(6), B => B(6), S => SEL, Y => Y(6));
   MUXES_7 : MUX21_305 port map( A => A(7), B => B(7), S => SEL, Y => Y(7));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT8_10 is

   port( A, B : in std_logic_vector (7 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (7 downto 0));

end MUX21_GENERIC_NBIT8_10;

architecture SYN_structural of MUX21_GENERIC_NBIT8_10 is

   component MUX21_297
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_298
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_299
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_300
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_301
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_302
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_303
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_304
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_304 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_303 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_302 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_301 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));
   MUXES_4 : MUX21_300 port map( A => A(4), B => B(4), S => SEL, Y => Y(4));
   MUXES_5 : MUX21_299 port map( A => A(5), B => B(5), S => SEL, Y => Y(5));
   MUXES_6 : MUX21_298 port map( A => A(6), B => B(6), S => SEL, Y => Y(6));
   MUXES_7 : MUX21_297 port map( A => A(7), B => B(7), S => SEL, Y => Y(7));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT8_9 is

   port( A, B : in std_logic_vector (7 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (7 downto 0));

end MUX21_GENERIC_NBIT8_9;

architecture SYN_structural of MUX21_GENERIC_NBIT8_9 is

   component MUX21_289
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_290
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_291
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_292
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_293
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_294
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_295
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_296
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_296 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_295 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_294 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_293 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));
   MUXES_4 : MUX21_292 port map( A => A(4), B => B(4), S => SEL, Y => Y(4));
   MUXES_5 : MUX21_291 port map( A => A(5), B => B(5), S => SEL, Y => Y(5));
   MUXES_6 : MUX21_290 port map( A => A(6), B => B(6), S => SEL, Y => Y(6));
   MUXES_7 : MUX21_289 port map( A => A(7), B => B(7), S => SEL, Y => Y(7));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT8_8 is

   port( A, B : in std_logic_vector (7 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (7 downto 0));

end MUX21_GENERIC_NBIT8_8;

architecture SYN_structural of MUX21_GENERIC_NBIT8_8 is

   component MUX21_281
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_282
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_283
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_284
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_285
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_286
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_287
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_288
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_288 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_287 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_286 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_285 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));
   MUXES_4 : MUX21_284 port map( A => A(4), B => B(4), S => SEL, Y => Y(4));
   MUXES_5 : MUX21_283 port map( A => A(5), B => B(5), S => SEL, Y => Y(5));
   MUXES_6 : MUX21_282 port map( A => A(6), B => B(6), S => SEL, Y => Y(6));
   MUXES_7 : MUX21_281 port map( A => A(7), B => B(7), S => SEL, Y => Y(7));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT8_7 is

   port( A, B : in std_logic_vector (7 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (7 downto 0));

end MUX21_GENERIC_NBIT8_7;

architecture SYN_structural of MUX21_GENERIC_NBIT8_7 is

   component MUX21_273
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_274
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_275
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_276
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_277
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_278
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_279
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_280
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_280 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_279 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_278 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_277 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));
   MUXES_4 : MUX21_276 port map( A => A(4), B => B(4), S => SEL, Y => Y(4));
   MUXES_5 : MUX21_275 port map( A => A(5), B => B(5), S => SEL, Y => Y(5));
   MUXES_6 : MUX21_274 port map( A => A(6), B => B(6), S => SEL, Y => Y(6));
   MUXES_7 : MUX21_273 port map( A => A(7), B => B(7), S => SEL, Y => Y(7));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT8_6 is

   port( A, B : in std_logic_vector (7 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (7 downto 0));

end MUX21_GENERIC_NBIT8_6;

architecture SYN_structural of MUX21_GENERIC_NBIT8_6 is

   component MUX21_265
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_266
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_267
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_268
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_269
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_270
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_271
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_272
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_272 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_271 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_270 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_269 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));
   MUXES_4 : MUX21_268 port map( A => A(4), B => B(4), S => SEL, Y => Y(4));
   MUXES_5 : MUX21_267 port map( A => A(5), B => B(5), S => SEL, Y => Y(5));
   MUXES_6 : MUX21_266 port map( A => A(6), B => B(6), S => SEL, Y => Y(6));
   MUXES_7 : MUX21_265 port map( A => A(7), B => B(7), S => SEL, Y => Y(7));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT8_5 is

   port( A, B : in std_logic_vector (7 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (7 downto 0));

end MUX21_GENERIC_NBIT8_5;

architecture SYN_structural of MUX21_GENERIC_NBIT8_5 is

   component MUX21_257
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_258
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_259
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_260
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_261
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_262
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_263
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_264
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_264 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_263 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_262 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_261 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));
   MUXES_4 : MUX21_260 port map( A => A(4), B => B(4), S => SEL, Y => Y(4));
   MUXES_5 : MUX21_259 port map( A => A(5), B => B(5), S => SEL, Y => Y(5));
   MUXES_6 : MUX21_258 port map( A => A(6), B => B(6), S => SEL, Y => Y(6));
   MUXES_7 : MUX21_257 port map( A => A(7), B => B(7), S => SEL, Y => Y(7));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT8_4 is

   port( A, B : in std_logic_vector (7 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (7 downto 0));

end MUX21_GENERIC_NBIT8_4;

architecture SYN_structural of MUX21_GENERIC_NBIT8_4 is

   component MUX21_249
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_250
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_251
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_252
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_253
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_254
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_255
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_256
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_256 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_255 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_254 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_253 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));
   MUXES_4 : MUX21_252 port map( A => A(4), B => B(4), S => SEL, Y => Y(4));
   MUXES_5 : MUX21_251 port map( A => A(5), B => B(5), S => SEL, Y => Y(5));
   MUXES_6 : MUX21_250 port map( A => A(6), B => B(6), S => SEL, Y => Y(6));
   MUXES_7 : MUX21_249 port map( A => A(7), B => B(7), S => SEL, Y => Y(7));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT8_3 is

   port( A, B : in std_logic_vector (7 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (7 downto 0));

end MUX21_GENERIC_NBIT8_3;

architecture SYN_structural of MUX21_GENERIC_NBIT8_3 is

   component MUX21_241
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_242
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_243
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_244
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_245
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_246
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_247
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_248
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_248 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_247 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_246 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_245 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));
   MUXES_4 : MUX21_244 port map( A => A(4), B => B(4), S => SEL, Y => Y(4));
   MUXES_5 : MUX21_243 port map( A => A(5), B => B(5), S => SEL, Y => Y(5));
   MUXES_6 : MUX21_242 port map( A => A(6), B => B(6), S => SEL, Y => Y(6));
   MUXES_7 : MUX21_241 port map( A => A(7), B => B(7), S => SEL, Y => Y(7));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT8_2 is

   port( A, B : in std_logic_vector (7 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (7 downto 0));

end MUX21_GENERIC_NBIT8_2;

architecture SYN_structural of MUX21_GENERIC_NBIT8_2 is

   component MUX21_233
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_234
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_235
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_236
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_237
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_238
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_239
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_240
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_240 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_239 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_238 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_237 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));
   MUXES_4 : MUX21_236 port map( A => A(4), B => B(4), S => SEL, Y => Y(4));
   MUXES_5 : MUX21_235 port map( A => A(5), B => B(5), S => SEL, Y => Y(5));
   MUXES_6 : MUX21_234 port map( A => A(6), B => B(6), S => SEL, Y => Y(6));
   MUXES_7 : MUX21_233 port map( A => A(7), B => B(7), S => SEL, Y => Y(7));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT8_1 is

   port( A, B : in std_logic_vector (7 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (7 downto 0));

end MUX21_GENERIC_NBIT8_1;

architecture SYN_structural of MUX21_GENERIC_NBIT8_1 is

   component MUX21_225
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_226
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_227
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_228
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_229
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_230
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_231
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_232
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_232 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_231 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_230 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_229 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));
   MUXES_4 : MUX21_228 port map( A => A(4), B => B(4), S => SEL, Y => Y(4));
   MUXES_5 : MUX21_227 port map( A => A(5), B => B(5), S => SEL, Y => Y(5));
   MUXES_6 : MUX21_226 port map( A => A(6), B => B(6), S => SEL, Y => Y(6));
   MUXES_7 : MUX21_225 port map( A => A(7), B => B(7), S => SEL, Y => Y(7));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_511 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_511;

architecture SYN_BEHAVIORAL of FA_511 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_510 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_510;

architecture SYN_BEHAVIORAL of FA_510 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_509 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_509;

architecture SYN_BEHAVIORAL of FA_509 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_508 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_508;

architecture SYN_BEHAVIORAL of FA_508 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_507 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_507;

architecture SYN_BEHAVIORAL of FA_507 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_506 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_506;

architecture SYN_BEHAVIORAL of FA_506 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_505 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_505;

architecture SYN_BEHAVIORAL of FA_505 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_504 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_504;

architecture SYN_BEHAVIORAL of FA_504 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_503 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_503;

architecture SYN_BEHAVIORAL of FA_503 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_502 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_502;

architecture SYN_BEHAVIORAL of FA_502 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_501 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_501;

architecture SYN_BEHAVIORAL of FA_501 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_500 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_500;

architecture SYN_BEHAVIORAL of FA_500 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_499 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_499;

architecture SYN_BEHAVIORAL of FA_499 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_498 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_498;

architecture SYN_BEHAVIORAL of FA_498 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_497 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_497;

architecture SYN_BEHAVIORAL of FA_497 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_496 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_496;

architecture SYN_BEHAVIORAL of FA_496 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_495 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_495;

architecture SYN_BEHAVIORAL of FA_495 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_494 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_494;

architecture SYN_BEHAVIORAL of FA_494 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_493 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_493;

architecture SYN_BEHAVIORAL of FA_493 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_492 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_492;

architecture SYN_BEHAVIORAL of FA_492 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_491 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_491;

architecture SYN_BEHAVIORAL of FA_491 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_490 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_490;

architecture SYN_BEHAVIORAL of FA_490 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_489 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_489;

architecture SYN_BEHAVIORAL of FA_489 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_488 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_488;

architecture SYN_BEHAVIORAL of FA_488 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_487 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_487;

architecture SYN_BEHAVIORAL of FA_487 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_486 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_486;

architecture SYN_BEHAVIORAL of FA_486 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_485 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_485;

architecture SYN_BEHAVIORAL of FA_485 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_484 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_484;

architecture SYN_BEHAVIORAL of FA_484 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_483 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_483;

architecture SYN_BEHAVIORAL of FA_483 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_482 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_482;

architecture SYN_BEHAVIORAL of FA_482 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_481 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_481;

architecture SYN_BEHAVIORAL of FA_481 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_480 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_480;

architecture SYN_BEHAVIORAL of FA_480 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_479 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_479;

architecture SYN_BEHAVIORAL of FA_479 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_478 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_478;

architecture SYN_BEHAVIORAL of FA_478 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_477 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_477;

architecture SYN_BEHAVIORAL of FA_477 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_476 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_476;

architecture SYN_BEHAVIORAL of FA_476 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_475 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_475;

architecture SYN_BEHAVIORAL of FA_475 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_474 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_474;

architecture SYN_BEHAVIORAL of FA_474 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_473 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_473;

architecture SYN_BEHAVIORAL of FA_473 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_472 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_472;

architecture SYN_BEHAVIORAL of FA_472 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_471 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_471;

architecture SYN_BEHAVIORAL of FA_471 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_470 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_470;

architecture SYN_BEHAVIORAL of FA_470 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_469 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_469;

architecture SYN_BEHAVIORAL of FA_469 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_468 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_468;

architecture SYN_BEHAVIORAL of FA_468 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_467 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_467;

architecture SYN_BEHAVIORAL of FA_467 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_466 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_466;

architecture SYN_BEHAVIORAL of FA_466 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_465 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_465;

architecture SYN_BEHAVIORAL of FA_465 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_464 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_464;

architecture SYN_BEHAVIORAL of FA_464 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_463 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_463;

architecture SYN_BEHAVIORAL of FA_463 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_462 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_462;

architecture SYN_BEHAVIORAL of FA_462 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_461 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_461;

architecture SYN_BEHAVIORAL of FA_461 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_460 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_460;

architecture SYN_BEHAVIORAL of FA_460 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_459 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_459;

architecture SYN_BEHAVIORAL of FA_459 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_458 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_458;

architecture SYN_BEHAVIORAL of FA_458 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_457 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_457;

architecture SYN_BEHAVIORAL of FA_457 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_456 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_456;

architecture SYN_BEHAVIORAL of FA_456 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_455 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_455;

architecture SYN_BEHAVIORAL of FA_455 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_454 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_454;

architecture SYN_BEHAVIORAL of FA_454 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_453 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_453;

architecture SYN_BEHAVIORAL of FA_453 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_452 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_452;

architecture SYN_BEHAVIORAL of FA_452 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_451 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_451;

architecture SYN_BEHAVIORAL of FA_451 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_450 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_450;

architecture SYN_BEHAVIORAL of FA_450 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_449 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_449;

architecture SYN_BEHAVIORAL of FA_449 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_448 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_448;

architecture SYN_BEHAVIORAL of FA_448 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_447 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_447;

architecture SYN_BEHAVIORAL of FA_447 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_446 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_446;

architecture SYN_BEHAVIORAL of FA_446 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_445 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_445;

architecture SYN_BEHAVIORAL of FA_445 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_444 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_444;

architecture SYN_BEHAVIORAL of FA_444 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_443 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_443;

architecture SYN_BEHAVIORAL of FA_443 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_442 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_442;

architecture SYN_BEHAVIORAL of FA_442 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_441 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_441;

architecture SYN_BEHAVIORAL of FA_441 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_440 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_440;

architecture SYN_BEHAVIORAL of FA_440 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_439 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_439;

architecture SYN_BEHAVIORAL of FA_439 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_438 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_438;

architecture SYN_BEHAVIORAL of FA_438 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_437 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_437;

architecture SYN_BEHAVIORAL of FA_437 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_436 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_436;

architecture SYN_BEHAVIORAL of FA_436 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_435 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_435;

architecture SYN_BEHAVIORAL of FA_435 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_434 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_434;

architecture SYN_BEHAVIORAL of FA_434 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_433 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_433;

architecture SYN_BEHAVIORAL of FA_433 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_432 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_432;

architecture SYN_BEHAVIORAL of FA_432 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_431 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_431;

architecture SYN_BEHAVIORAL of FA_431 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_430 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_430;

architecture SYN_BEHAVIORAL of FA_430 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_429 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_429;

architecture SYN_BEHAVIORAL of FA_429 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_428 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_428;

architecture SYN_BEHAVIORAL of FA_428 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_427 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_427;

architecture SYN_BEHAVIORAL of FA_427 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_426 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_426;

architecture SYN_BEHAVIORAL of FA_426 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_425 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_425;

architecture SYN_BEHAVIORAL of FA_425 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_424 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_424;

architecture SYN_BEHAVIORAL of FA_424 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_423 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_423;

architecture SYN_BEHAVIORAL of FA_423 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_422 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_422;

architecture SYN_BEHAVIORAL of FA_422 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_421 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_421;

architecture SYN_BEHAVIORAL of FA_421 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_420 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_420;

architecture SYN_BEHAVIORAL of FA_420 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_419 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_419;

architecture SYN_BEHAVIORAL of FA_419 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_418 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_418;

architecture SYN_BEHAVIORAL of FA_418 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_417 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_417;

architecture SYN_BEHAVIORAL of FA_417 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_416 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_416;

architecture SYN_BEHAVIORAL of FA_416 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_415 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_415;

architecture SYN_BEHAVIORAL of FA_415 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_414 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_414;

architecture SYN_BEHAVIORAL of FA_414 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_413 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_413;

architecture SYN_BEHAVIORAL of FA_413 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_412 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_412;

architecture SYN_BEHAVIORAL of FA_412 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_411 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_411;

architecture SYN_BEHAVIORAL of FA_411 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_410 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_410;

architecture SYN_BEHAVIORAL of FA_410 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_409 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_409;

architecture SYN_BEHAVIORAL of FA_409 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_408 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_408;

architecture SYN_BEHAVIORAL of FA_408 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_407 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_407;

architecture SYN_BEHAVIORAL of FA_407 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_406 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_406;

architecture SYN_BEHAVIORAL of FA_406 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_405 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_405;

architecture SYN_BEHAVIORAL of FA_405 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_404 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_404;

architecture SYN_BEHAVIORAL of FA_404 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_403 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_403;

architecture SYN_BEHAVIORAL of FA_403 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_402 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_402;

architecture SYN_BEHAVIORAL of FA_402 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_401 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_401;

architecture SYN_BEHAVIORAL of FA_401 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_400 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_400;

architecture SYN_BEHAVIORAL of FA_400 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_399 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_399;

architecture SYN_BEHAVIORAL of FA_399 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_398 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_398;

architecture SYN_BEHAVIORAL of FA_398 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_397 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_397;

architecture SYN_BEHAVIORAL of FA_397 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_396 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_396;

architecture SYN_BEHAVIORAL of FA_396 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_395 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_395;

architecture SYN_BEHAVIORAL of FA_395 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_394 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_394;

architecture SYN_BEHAVIORAL of FA_394 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_393 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_393;

architecture SYN_BEHAVIORAL of FA_393 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_392 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_392;

architecture SYN_BEHAVIORAL of FA_392 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_391 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_391;

architecture SYN_BEHAVIORAL of FA_391 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_390 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_390;

architecture SYN_BEHAVIORAL of FA_390 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_389 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_389;

architecture SYN_BEHAVIORAL of FA_389 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_388 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_388;

architecture SYN_BEHAVIORAL of FA_388 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_387 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_387;

architecture SYN_BEHAVIORAL of FA_387 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_386 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_386;

architecture SYN_BEHAVIORAL of FA_386 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_385 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_385;

architecture SYN_BEHAVIORAL of FA_385 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_384 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_384;

architecture SYN_BEHAVIORAL of FA_384 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_383 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_383;

architecture SYN_BEHAVIORAL of FA_383 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_382 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_382;

architecture SYN_BEHAVIORAL of FA_382 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_381 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_381;

architecture SYN_BEHAVIORAL of FA_381 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_380 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_380;

architecture SYN_BEHAVIORAL of FA_380 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_379 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_379;

architecture SYN_BEHAVIORAL of FA_379 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_378 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_378;

architecture SYN_BEHAVIORAL of FA_378 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_377 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_377;

architecture SYN_BEHAVIORAL of FA_377 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_376 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_376;

architecture SYN_BEHAVIORAL of FA_376 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_375 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_375;

architecture SYN_BEHAVIORAL of FA_375 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_374 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_374;

architecture SYN_BEHAVIORAL of FA_374 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_373 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_373;

architecture SYN_BEHAVIORAL of FA_373 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_372 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_372;

architecture SYN_BEHAVIORAL of FA_372 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_371 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_371;

architecture SYN_BEHAVIORAL of FA_371 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_370 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_370;

architecture SYN_BEHAVIORAL of FA_370 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_369 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_369;

architecture SYN_BEHAVIORAL of FA_369 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_368 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_368;

architecture SYN_BEHAVIORAL of FA_368 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_367 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_367;

architecture SYN_BEHAVIORAL of FA_367 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_366 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_366;

architecture SYN_BEHAVIORAL of FA_366 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_365 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_365;

architecture SYN_BEHAVIORAL of FA_365 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_364 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_364;

architecture SYN_BEHAVIORAL of FA_364 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_363 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_363;

architecture SYN_BEHAVIORAL of FA_363 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_362 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_362;

architecture SYN_BEHAVIORAL of FA_362 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_361 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_361;

architecture SYN_BEHAVIORAL of FA_361 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_360 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_360;

architecture SYN_BEHAVIORAL of FA_360 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_359 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_359;

architecture SYN_BEHAVIORAL of FA_359 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_358 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_358;

architecture SYN_BEHAVIORAL of FA_358 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_357 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_357;

architecture SYN_BEHAVIORAL of FA_357 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_356 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_356;

architecture SYN_BEHAVIORAL of FA_356 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_355 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_355;

architecture SYN_BEHAVIORAL of FA_355 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_354 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_354;

architecture SYN_BEHAVIORAL of FA_354 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_353 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_353;

architecture SYN_BEHAVIORAL of FA_353 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_352 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_352;

architecture SYN_BEHAVIORAL of FA_352 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_351 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_351;

architecture SYN_BEHAVIORAL of FA_351 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_350 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_350;

architecture SYN_BEHAVIORAL of FA_350 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_349 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_349;

architecture SYN_BEHAVIORAL of FA_349 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_348 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_348;

architecture SYN_BEHAVIORAL of FA_348 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_347 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_347;

architecture SYN_BEHAVIORAL of FA_347 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_346 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_346;

architecture SYN_BEHAVIORAL of FA_346 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_345 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_345;

architecture SYN_BEHAVIORAL of FA_345 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_344 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_344;

architecture SYN_BEHAVIORAL of FA_344 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_343 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_343;

architecture SYN_BEHAVIORAL of FA_343 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_342 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_342;

architecture SYN_BEHAVIORAL of FA_342 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_341 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_341;

architecture SYN_BEHAVIORAL of FA_341 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_340 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_340;

architecture SYN_BEHAVIORAL of FA_340 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_339 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_339;

architecture SYN_BEHAVIORAL of FA_339 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_338 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_338;

architecture SYN_BEHAVIORAL of FA_338 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_337 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_337;

architecture SYN_BEHAVIORAL of FA_337 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_336 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_336;

architecture SYN_BEHAVIORAL of FA_336 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_335 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_335;

architecture SYN_BEHAVIORAL of FA_335 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_334 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_334;

architecture SYN_BEHAVIORAL of FA_334 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_333 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_333;

architecture SYN_BEHAVIORAL of FA_333 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_332 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_332;

architecture SYN_BEHAVIORAL of FA_332 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_331 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_331;

architecture SYN_BEHAVIORAL of FA_331 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_330 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_330;

architecture SYN_BEHAVIORAL of FA_330 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_329 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_329;

architecture SYN_BEHAVIORAL of FA_329 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_328 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_328;

architecture SYN_BEHAVIORAL of FA_328 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_327 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_327;

architecture SYN_BEHAVIORAL of FA_327 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_326 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_326;

architecture SYN_BEHAVIORAL of FA_326 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_325 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_325;

architecture SYN_BEHAVIORAL of FA_325 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_324 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_324;

architecture SYN_BEHAVIORAL of FA_324 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_323 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_323;

architecture SYN_BEHAVIORAL of FA_323 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_322 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_322;

architecture SYN_BEHAVIORAL of FA_322 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_321 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_321;

architecture SYN_BEHAVIORAL of FA_321 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_320 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_320;

architecture SYN_BEHAVIORAL of FA_320 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_319 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_319;

architecture SYN_BEHAVIORAL of FA_319 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_318 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_318;

architecture SYN_BEHAVIORAL of FA_318 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_317 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_317;

architecture SYN_BEHAVIORAL of FA_317 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_316 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_316;

architecture SYN_BEHAVIORAL of FA_316 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_315 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_315;

architecture SYN_BEHAVIORAL of FA_315 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_314 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_314;

architecture SYN_BEHAVIORAL of FA_314 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_313 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_313;

architecture SYN_BEHAVIORAL of FA_313 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_312 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_312;

architecture SYN_BEHAVIORAL of FA_312 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_311 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_311;

architecture SYN_BEHAVIORAL of FA_311 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_310 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_310;

architecture SYN_BEHAVIORAL of FA_310 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_309 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_309;

architecture SYN_BEHAVIORAL of FA_309 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_308 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_308;

architecture SYN_BEHAVIORAL of FA_308 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_307 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_307;

architecture SYN_BEHAVIORAL of FA_307 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_306 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_306;

architecture SYN_BEHAVIORAL of FA_306 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_305 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_305;

architecture SYN_BEHAVIORAL of FA_305 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_304 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_304;

architecture SYN_BEHAVIORAL of FA_304 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_303 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_303;

architecture SYN_BEHAVIORAL of FA_303 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_302 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_302;

architecture SYN_BEHAVIORAL of FA_302 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_301 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_301;

architecture SYN_BEHAVIORAL of FA_301 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_300 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_300;

architecture SYN_BEHAVIORAL of FA_300 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_299 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_299;

architecture SYN_BEHAVIORAL of FA_299 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_298 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_298;

architecture SYN_BEHAVIORAL of FA_298 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_297 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_297;

architecture SYN_BEHAVIORAL of FA_297 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_296 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_296;

architecture SYN_BEHAVIORAL of FA_296 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_295 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_295;

architecture SYN_BEHAVIORAL of FA_295 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_294 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_294;

architecture SYN_BEHAVIORAL of FA_294 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_293 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_293;

architecture SYN_BEHAVIORAL of FA_293 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_292 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_292;

architecture SYN_BEHAVIORAL of FA_292 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_291 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_291;

architecture SYN_BEHAVIORAL of FA_291 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_290 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_290;

architecture SYN_BEHAVIORAL of FA_290 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_289 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_289;

architecture SYN_BEHAVIORAL of FA_289 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_288 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_288;

architecture SYN_BEHAVIORAL of FA_288 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_287 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_287;

architecture SYN_BEHAVIORAL of FA_287 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_286 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_286;

architecture SYN_BEHAVIORAL of FA_286 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_285 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_285;

architecture SYN_BEHAVIORAL of FA_285 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_284 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_284;

architecture SYN_BEHAVIORAL of FA_284 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_283 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_283;

architecture SYN_BEHAVIORAL of FA_283 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_282 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_282;

architecture SYN_BEHAVIORAL of FA_282 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_281 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_281;

architecture SYN_BEHAVIORAL of FA_281 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_280 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_280;

architecture SYN_BEHAVIORAL of FA_280 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_279 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_279;

architecture SYN_BEHAVIORAL of FA_279 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_278 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_278;

architecture SYN_BEHAVIORAL of FA_278 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_277 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_277;

architecture SYN_BEHAVIORAL of FA_277 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_276 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_276;

architecture SYN_BEHAVIORAL of FA_276 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_275 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_275;

architecture SYN_BEHAVIORAL of FA_275 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_274 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_274;

architecture SYN_BEHAVIORAL of FA_274 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_273 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_273;

architecture SYN_BEHAVIORAL of FA_273 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_272 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_272;

architecture SYN_BEHAVIORAL of FA_272 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_271 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_271;

architecture SYN_BEHAVIORAL of FA_271 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_270 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_270;

architecture SYN_BEHAVIORAL of FA_270 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_269 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_269;

architecture SYN_BEHAVIORAL of FA_269 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_268 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_268;

architecture SYN_BEHAVIORAL of FA_268 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_267 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_267;

architecture SYN_BEHAVIORAL of FA_267 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_266 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_266;

architecture SYN_BEHAVIORAL of FA_266 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_265 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_265;

architecture SYN_BEHAVIORAL of FA_265 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_264 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_264;

architecture SYN_BEHAVIORAL of FA_264 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_263 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_263;

architecture SYN_BEHAVIORAL of FA_263 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_262 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_262;

architecture SYN_BEHAVIORAL of FA_262 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_261 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_261;

architecture SYN_BEHAVIORAL of FA_261 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_260 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_260;

architecture SYN_BEHAVIORAL of FA_260 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_259 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_259;

architecture SYN_BEHAVIORAL of FA_259 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_258 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_258;

architecture SYN_BEHAVIORAL of FA_258 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_257 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_257;

architecture SYN_BEHAVIORAL of FA_257 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_256 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_256;

architecture SYN_BEHAVIORAL of FA_256 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_255 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_255;

architecture SYN_BEHAVIORAL of FA_255 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_254 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_254;

architecture SYN_BEHAVIORAL of FA_254 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_253 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_253;

architecture SYN_BEHAVIORAL of FA_253 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_252 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_252;

architecture SYN_BEHAVIORAL of FA_252 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_251 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_251;

architecture SYN_BEHAVIORAL of FA_251 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_250 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_250;

architecture SYN_BEHAVIORAL of FA_250 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_249 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_249;

architecture SYN_BEHAVIORAL of FA_249 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_248 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_248;

architecture SYN_BEHAVIORAL of FA_248 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_247 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_247;

architecture SYN_BEHAVIORAL of FA_247 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_246 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_246;

architecture SYN_BEHAVIORAL of FA_246 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_245 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_245;

architecture SYN_BEHAVIORAL of FA_245 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_244 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_244;

architecture SYN_BEHAVIORAL of FA_244 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_243 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_243;

architecture SYN_BEHAVIORAL of FA_243 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_242 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_242;

architecture SYN_BEHAVIORAL of FA_242 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_241 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_241;

architecture SYN_BEHAVIORAL of FA_241 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_240 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_240;

architecture SYN_BEHAVIORAL of FA_240 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_239 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_239;

architecture SYN_BEHAVIORAL of FA_239 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_238 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_238;

architecture SYN_BEHAVIORAL of FA_238 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_237 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_237;

architecture SYN_BEHAVIORAL of FA_237 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_236 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_236;

architecture SYN_BEHAVIORAL of FA_236 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_235 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_235;

architecture SYN_BEHAVIORAL of FA_235 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_234 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_234;

architecture SYN_BEHAVIORAL of FA_234 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_233 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_233;

architecture SYN_BEHAVIORAL of FA_233 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_232 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_232;

architecture SYN_BEHAVIORAL of FA_232 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_231 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_231;

architecture SYN_BEHAVIORAL of FA_231 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_230 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_230;

architecture SYN_BEHAVIORAL of FA_230 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_229 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_229;

architecture SYN_BEHAVIORAL of FA_229 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_228 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_228;

architecture SYN_BEHAVIORAL of FA_228 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_227 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_227;

architecture SYN_BEHAVIORAL of FA_227 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_226 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_226;

architecture SYN_BEHAVIORAL of FA_226 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_225 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_225;

architecture SYN_BEHAVIORAL of FA_225 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_224 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_224;

architecture SYN_BEHAVIORAL of FA_224 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_223 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_223;

architecture SYN_BEHAVIORAL of FA_223 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_222 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_222;

architecture SYN_BEHAVIORAL of FA_222 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_221 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_221;

architecture SYN_BEHAVIORAL of FA_221 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_220 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_220;

architecture SYN_BEHAVIORAL of FA_220 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_219 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_219;

architecture SYN_BEHAVIORAL of FA_219 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_218 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_218;

architecture SYN_BEHAVIORAL of FA_218 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_217 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_217;

architecture SYN_BEHAVIORAL of FA_217 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_216 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_216;

architecture SYN_BEHAVIORAL of FA_216 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_215 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_215;

architecture SYN_BEHAVIORAL of FA_215 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_214 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_214;

architecture SYN_BEHAVIORAL of FA_214 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_213 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_213;

architecture SYN_BEHAVIORAL of FA_213 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_212 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_212;

architecture SYN_BEHAVIORAL of FA_212 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_211 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_211;

architecture SYN_BEHAVIORAL of FA_211 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_210 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_210;

architecture SYN_BEHAVIORAL of FA_210 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_209 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_209;

architecture SYN_BEHAVIORAL of FA_209 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_208 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_208;

architecture SYN_BEHAVIORAL of FA_208 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_207 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_207;

architecture SYN_BEHAVIORAL of FA_207 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_206 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_206;

architecture SYN_BEHAVIORAL of FA_206 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_205 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_205;

architecture SYN_BEHAVIORAL of FA_205 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_204 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_204;

architecture SYN_BEHAVIORAL of FA_204 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_203 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_203;

architecture SYN_BEHAVIORAL of FA_203 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_202 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_202;

architecture SYN_BEHAVIORAL of FA_202 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_201 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_201;

architecture SYN_BEHAVIORAL of FA_201 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_200 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_200;

architecture SYN_BEHAVIORAL of FA_200 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_199 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_199;

architecture SYN_BEHAVIORAL of FA_199 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_198 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_198;

architecture SYN_BEHAVIORAL of FA_198 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_197 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_197;

architecture SYN_BEHAVIORAL of FA_197 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_196 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_196;

architecture SYN_BEHAVIORAL of FA_196 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_195 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_195;

architecture SYN_BEHAVIORAL of FA_195 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_194 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_194;

architecture SYN_BEHAVIORAL of FA_194 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_193 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_193;

architecture SYN_BEHAVIORAL of FA_193 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_192 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_192;

architecture SYN_BEHAVIORAL of FA_192 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_191 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_191;

architecture SYN_BEHAVIORAL of FA_191 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_190 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_190;

architecture SYN_BEHAVIORAL of FA_190 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_189 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_189;

architecture SYN_BEHAVIORAL of FA_189 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_188 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_188;

architecture SYN_BEHAVIORAL of FA_188 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_187 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_187;

architecture SYN_BEHAVIORAL of FA_187 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_186 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_186;

architecture SYN_BEHAVIORAL of FA_186 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_185 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_185;

architecture SYN_BEHAVIORAL of FA_185 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_184 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_184;

architecture SYN_BEHAVIORAL of FA_184 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_183 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_183;

architecture SYN_BEHAVIORAL of FA_183 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_182 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_182;

architecture SYN_BEHAVIORAL of FA_182 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_181 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_181;

architecture SYN_BEHAVIORAL of FA_181 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_180 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_180;

architecture SYN_BEHAVIORAL of FA_180 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_179 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_179;

architecture SYN_BEHAVIORAL of FA_179 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_178 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_178;

architecture SYN_BEHAVIORAL of FA_178 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_177 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_177;

architecture SYN_BEHAVIORAL of FA_177 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_176 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_176;

architecture SYN_BEHAVIORAL of FA_176 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_175 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_175;

architecture SYN_BEHAVIORAL of FA_175 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_174 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_174;

architecture SYN_BEHAVIORAL of FA_174 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_173 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_173;

architecture SYN_BEHAVIORAL of FA_173 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_172 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_172;

architecture SYN_BEHAVIORAL of FA_172 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_171 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_171;

architecture SYN_BEHAVIORAL of FA_171 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_170 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_170;

architecture SYN_BEHAVIORAL of FA_170 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_169 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_169;

architecture SYN_BEHAVIORAL of FA_169 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_168 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_168;

architecture SYN_BEHAVIORAL of FA_168 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_167 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_167;

architecture SYN_BEHAVIORAL of FA_167 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_166 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_166;

architecture SYN_BEHAVIORAL of FA_166 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_165 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_165;

architecture SYN_BEHAVIORAL of FA_165 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_164 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_164;

architecture SYN_BEHAVIORAL of FA_164 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_163 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_163;

architecture SYN_BEHAVIORAL of FA_163 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_162 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_162;

architecture SYN_BEHAVIORAL of FA_162 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_161 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_161;

architecture SYN_BEHAVIORAL of FA_161 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_160 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_160;

architecture SYN_BEHAVIORAL of FA_160 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_159 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_159;

architecture SYN_BEHAVIORAL of FA_159 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_158 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_158;

architecture SYN_BEHAVIORAL of FA_158 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_157 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_157;

architecture SYN_BEHAVIORAL of FA_157 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_156 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_156;

architecture SYN_BEHAVIORAL of FA_156 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_155 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_155;

architecture SYN_BEHAVIORAL of FA_155 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_154 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_154;

architecture SYN_BEHAVIORAL of FA_154 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_153 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_153;

architecture SYN_BEHAVIORAL of FA_153 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_152 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_152;

architecture SYN_BEHAVIORAL of FA_152 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_151 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_151;

architecture SYN_BEHAVIORAL of FA_151 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_150 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_150;

architecture SYN_BEHAVIORAL of FA_150 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_149 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_149;

architecture SYN_BEHAVIORAL of FA_149 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_148 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_148;

architecture SYN_BEHAVIORAL of FA_148 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_147 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_147;

architecture SYN_BEHAVIORAL of FA_147 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_146 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_146;

architecture SYN_BEHAVIORAL of FA_146 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_145 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_145;

architecture SYN_BEHAVIORAL of FA_145 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_144 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_144;

architecture SYN_BEHAVIORAL of FA_144 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_143 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_143;

architecture SYN_BEHAVIORAL of FA_143 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_142 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_142;

architecture SYN_BEHAVIORAL of FA_142 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_141 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_141;

architecture SYN_BEHAVIORAL of FA_141 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_140 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_140;

architecture SYN_BEHAVIORAL of FA_140 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_139 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_139;

architecture SYN_BEHAVIORAL of FA_139 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_138 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_138;

architecture SYN_BEHAVIORAL of FA_138 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_137 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_137;

architecture SYN_BEHAVIORAL of FA_137 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_136 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_136;

architecture SYN_BEHAVIORAL of FA_136 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_135 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_135;

architecture SYN_BEHAVIORAL of FA_135 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_134 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_134;

architecture SYN_BEHAVIORAL of FA_134 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_133 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_133;

architecture SYN_BEHAVIORAL of FA_133 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_132 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_132;

architecture SYN_BEHAVIORAL of FA_132 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_131 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_131;

architecture SYN_BEHAVIORAL of FA_131 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_130 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_130;

architecture SYN_BEHAVIORAL of FA_130 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_129 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_129;

architecture SYN_BEHAVIORAL of FA_129 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_128 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_128;

architecture SYN_BEHAVIORAL of FA_128 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_127 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_127;

architecture SYN_BEHAVIORAL of FA_127 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_126 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_126;

architecture SYN_BEHAVIORAL of FA_126 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_125 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_125;

architecture SYN_BEHAVIORAL of FA_125 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_124 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_124;

architecture SYN_BEHAVIORAL of FA_124 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_123 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_123;

architecture SYN_BEHAVIORAL of FA_123 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_122 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_122;

architecture SYN_BEHAVIORAL of FA_122 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_121 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_121;

architecture SYN_BEHAVIORAL of FA_121 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_120 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_120;

architecture SYN_BEHAVIORAL of FA_120 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_119 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_119;

architecture SYN_BEHAVIORAL of FA_119 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_118 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_118;

architecture SYN_BEHAVIORAL of FA_118 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_117 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_117;

architecture SYN_BEHAVIORAL of FA_117 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_116 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_116;

architecture SYN_BEHAVIORAL of FA_116 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_115 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_115;

architecture SYN_BEHAVIORAL of FA_115 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_114 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_114;

architecture SYN_BEHAVIORAL of FA_114 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_113 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_113;

architecture SYN_BEHAVIORAL of FA_113 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_112 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_112;

architecture SYN_BEHAVIORAL of FA_112 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_111 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_111;

architecture SYN_BEHAVIORAL of FA_111 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_110 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_110;

architecture SYN_BEHAVIORAL of FA_110 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_109 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_109;

architecture SYN_BEHAVIORAL of FA_109 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_108 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_108;

architecture SYN_BEHAVIORAL of FA_108 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_107 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_107;

architecture SYN_BEHAVIORAL of FA_107 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_106 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_106;

architecture SYN_BEHAVIORAL of FA_106 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_105 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_105;

architecture SYN_BEHAVIORAL of FA_105 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_104 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_104;

architecture SYN_BEHAVIORAL of FA_104 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_103 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_103;

architecture SYN_BEHAVIORAL of FA_103 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_102 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_102;

architecture SYN_BEHAVIORAL of FA_102 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_101 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_101;

architecture SYN_BEHAVIORAL of FA_101 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_100 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_100;

architecture SYN_BEHAVIORAL of FA_100 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_99 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_99;

architecture SYN_BEHAVIORAL of FA_99 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_98 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_98;

architecture SYN_BEHAVIORAL of FA_98 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_97 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_97;

architecture SYN_BEHAVIORAL of FA_97 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_96 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_96;

architecture SYN_BEHAVIORAL of FA_96 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_95 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_95;

architecture SYN_BEHAVIORAL of FA_95 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_94 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_94;

architecture SYN_BEHAVIORAL of FA_94 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_93 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_93;

architecture SYN_BEHAVIORAL of FA_93 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_92 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_92;

architecture SYN_BEHAVIORAL of FA_92 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_91 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_91;

architecture SYN_BEHAVIORAL of FA_91 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_90 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_90;

architecture SYN_BEHAVIORAL of FA_90 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_89 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_89;

architecture SYN_BEHAVIORAL of FA_89 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_88 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_88;

architecture SYN_BEHAVIORAL of FA_88 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_87 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_87;

architecture SYN_BEHAVIORAL of FA_87 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_86 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_86;

architecture SYN_BEHAVIORAL of FA_86 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_85 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_85;

architecture SYN_BEHAVIORAL of FA_85 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_84 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_84;

architecture SYN_BEHAVIORAL of FA_84 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_83 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_83;

architecture SYN_BEHAVIORAL of FA_83 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_82 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_82;

architecture SYN_BEHAVIORAL of FA_82 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_81 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_81;

architecture SYN_BEHAVIORAL of FA_81 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_80 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_80;

architecture SYN_BEHAVIORAL of FA_80 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_79 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_79;

architecture SYN_BEHAVIORAL of FA_79 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_78 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_78;

architecture SYN_BEHAVIORAL of FA_78 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_77 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_77;

architecture SYN_BEHAVIORAL of FA_77 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_76 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_76;

architecture SYN_BEHAVIORAL of FA_76 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_75 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_75;

architecture SYN_BEHAVIORAL of FA_75 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_74 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_74;

architecture SYN_BEHAVIORAL of FA_74 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_73 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_73;

architecture SYN_BEHAVIORAL of FA_73 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_72 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_72;

architecture SYN_BEHAVIORAL of FA_72 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_71 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_71;

architecture SYN_BEHAVIORAL of FA_71 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_70 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_70;

architecture SYN_BEHAVIORAL of FA_70 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_69 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_69;

architecture SYN_BEHAVIORAL of FA_69 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_68 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_68;

architecture SYN_BEHAVIORAL of FA_68 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_67 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_67;

architecture SYN_BEHAVIORAL of FA_67 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_66 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_66;

architecture SYN_BEHAVIORAL of FA_66 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_65 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_65;

architecture SYN_BEHAVIORAL of FA_65 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_64 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_64;

architecture SYN_BEHAVIORAL of FA_64 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_63 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_63;

architecture SYN_BEHAVIORAL of FA_63 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_62 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_62;

architecture SYN_BEHAVIORAL of FA_62 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_61 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_61;

architecture SYN_BEHAVIORAL of FA_61 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_60 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_60;

architecture SYN_BEHAVIORAL of FA_60 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_59 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_59;

architecture SYN_BEHAVIORAL of FA_59 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_58 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_58;

architecture SYN_BEHAVIORAL of FA_58 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_57 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_57;

architecture SYN_BEHAVIORAL of FA_57 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_56 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_56;

architecture SYN_BEHAVIORAL of FA_56 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_55 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_55;

architecture SYN_BEHAVIORAL of FA_55 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_54 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_54;

architecture SYN_BEHAVIORAL of FA_54 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_53 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_53;

architecture SYN_BEHAVIORAL of FA_53 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_52 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_52;

architecture SYN_BEHAVIORAL of FA_52 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_51 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_51;

architecture SYN_BEHAVIORAL of FA_51 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_50 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_50;

architecture SYN_BEHAVIORAL of FA_50 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_49 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_49;

architecture SYN_BEHAVIORAL of FA_49 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_48 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_48;

architecture SYN_BEHAVIORAL of FA_48 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_47 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_47;

architecture SYN_BEHAVIORAL of FA_47 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_46 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_46;

architecture SYN_BEHAVIORAL of FA_46 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_45 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_45;

architecture SYN_BEHAVIORAL of FA_45 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_44 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_44;

architecture SYN_BEHAVIORAL of FA_44 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_43 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_43;

architecture SYN_BEHAVIORAL of FA_43 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_42 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_42;

architecture SYN_BEHAVIORAL of FA_42 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_41 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_41;

architecture SYN_BEHAVIORAL of FA_41 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_40 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_40;

architecture SYN_BEHAVIORAL of FA_40 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_39 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_39;

architecture SYN_BEHAVIORAL of FA_39 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_38 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_38;

architecture SYN_BEHAVIORAL of FA_38 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_37 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_37;

architecture SYN_BEHAVIORAL of FA_37 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_36 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_36;

architecture SYN_BEHAVIORAL of FA_36 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_35 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_35;

architecture SYN_BEHAVIORAL of FA_35 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_34 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_34;

architecture SYN_BEHAVIORAL of FA_34 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_33 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_33;

architecture SYN_BEHAVIORAL of FA_33 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_32 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_32;

architecture SYN_BEHAVIORAL of FA_32 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_31 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_31;

architecture SYN_BEHAVIORAL of FA_31 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_30 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_30;

architecture SYN_BEHAVIORAL of FA_30 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_29 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_29;

architecture SYN_BEHAVIORAL of FA_29 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_28 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_28;

architecture SYN_BEHAVIORAL of FA_28 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_27 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_27;

architecture SYN_BEHAVIORAL of FA_27 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_26 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_26;

architecture SYN_BEHAVIORAL of FA_26 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_25 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_25;

architecture SYN_BEHAVIORAL of FA_25 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_24 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_24;

architecture SYN_BEHAVIORAL of FA_24 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_23 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_23;

architecture SYN_BEHAVIORAL of FA_23 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_22 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_22;

architecture SYN_BEHAVIORAL of FA_22 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_21 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_21;

architecture SYN_BEHAVIORAL of FA_21 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_20 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_20;

architecture SYN_BEHAVIORAL of FA_20 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_19 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_19;

architecture SYN_BEHAVIORAL of FA_19 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_18 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_18;

architecture SYN_BEHAVIORAL of FA_18 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_17 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_17;

architecture SYN_BEHAVIORAL of FA_17 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_16 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_16;

architecture SYN_BEHAVIORAL of FA_16 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_15 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_15;

architecture SYN_BEHAVIORAL of FA_15 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_14 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_14;

architecture SYN_BEHAVIORAL of FA_14 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_13 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_13;

architecture SYN_BEHAVIORAL of FA_13 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_12 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_12;

architecture SYN_BEHAVIORAL of FA_12 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_11 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_11;

architecture SYN_BEHAVIORAL of FA_11 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_10 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_10;

architecture SYN_BEHAVIORAL of FA_10 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_9 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_9;

architecture SYN_BEHAVIORAL of FA_9 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_8 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_8;

architecture SYN_BEHAVIORAL of FA_8 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_7 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_7;

architecture SYN_BEHAVIORAL of FA_7 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_6 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_6;

architecture SYN_BEHAVIORAL of FA_6 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_5 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_5;

architecture SYN_BEHAVIORAL of FA_5 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_4 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_4;

architecture SYN_BEHAVIORAL of FA_4 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_3 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_3;

architecture SYN_BEHAVIORAL of FA_3 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_2 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2;

architecture SYN_BEHAVIORAL of FA_2 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_1 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1;

architecture SYN_BEHAVIORAL of FA_1 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n5, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n5, B2 => Ci, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity sum_generator_n_bit64_n_CSB16_2 is

   port( A, B : in std_logic_vector (63 downto 0);  C_in : in std_logic_vector 
         (15 downto 0);  S : out std_logic_vector (63 downto 0));

end sum_generator_n_bit64_n_CSB16_2;

architecture SYN_STRUCTURAL of sum_generator_n_bit64_n_CSB16_2 is

   component carry_select_block_n4_17
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_n4_18
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_n4_19
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_n4_20
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_n4_21
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_n4_22
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_n4_23
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_n4_24
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_n4_25
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_n4_26
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_n4_27
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_n4_28
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_n4_29
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_n4_30
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_n4_31
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_n4_32
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;

begin
   
   csb_0 : carry_select_block_n4_32 port map( A(3) => A(3), A(2) => A(2), A(1) 
                           => A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), 
                           B(1) => B(1), B(0) => B(0), C_sel => C_in(0), S(3) 
                           => S(3), S(2) => S(2), S(1) => S(1), S(0) => S(0));
   csb_1 : carry_select_block_n4_31 port map( A(3) => A(7), A(2) => A(6), A(1) 
                           => A(5), A(0) => A(4), B(3) => B(7), B(2) => B(6), 
                           B(1) => B(5), B(0) => B(4), C_sel => C_in(1), S(3) 
                           => S(7), S(2) => S(6), S(1) => S(5), S(0) => S(4));
   csb_2 : carry_select_block_n4_30 port map( A(3) => A(11), A(2) => A(10), 
                           A(1) => A(9), A(0) => A(8), B(3) => B(11), B(2) => 
                           B(10), B(1) => B(9), B(0) => B(8), C_sel => C_in(2),
                           S(3) => S(11), S(2) => S(10), S(1) => S(9), S(0) => 
                           S(8));
   csb_3 : carry_select_block_n4_29 port map( A(3) => A(15), A(2) => A(14), 
                           A(1) => A(13), A(0) => A(12), B(3) => B(15), B(2) =>
                           B(14), B(1) => B(13), B(0) => B(12), C_sel => 
                           C_in(3), S(3) => S(15), S(2) => S(14), S(1) => S(13)
                           , S(0) => S(12));
   csb_4 : carry_select_block_n4_28 port map( A(3) => A(19), A(2) => A(18), 
                           A(1) => A(17), A(0) => A(16), B(3) => B(19), B(2) =>
                           B(18), B(1) => B(17), B(0) => B(16), C_sel => 
                           C_in(4), S(3) => S(19), S(2) => S(18), S(1) => S(17)
                           , S(0) => S(16));
   csb_5 : carry_select_block_n4_27 port map( A(3) => A(23), A(2) => A(22), 
                           A(1) => A(21), A(0) => A(20), B(3) => B(23), B(2) =>
                           B(22), B(1) => B(21), B(0) => B(20), C_sel => 
                           C_in(5), S(3) => S(23), S(2) => S(22), S(1) => S(21)
                           , S(0) => S(20));
   csb_6 : carry_select_block_n4_26 port map( A(3) => A(27), A(2) => A(26), 
                           A(1) => A(25), A(0) => A(24), B(3) => B(27), B(2) =>
                           B(26), B(1) => B(25), B(0) => B(24), C_sel => 
                           C_in(6), S(3) => S(27), S(2) => S(26), S(1) => S(25)
                           , S(0) => S(24));
   csb_7 : carry_select_block_n4_25 port map( A(3) => A(31), A(2) => A(30), 
                           A(1) => A(29), A(0) => A(28), B(3) => B(31), B(2) =>
                           B(30), B(1) => B(29), B(0) => B(28), C_sel => 
                           C_in(7), S(3) => S(31), S(2) => S(30), S(1) => S(29)
                           , S(0) => S(28));
   csb_8 : carry_select_block_n4_24 port map( A(3) => A(35), A(2) => A(34), 
                           A(1) => A(33), A(0) => A(32), B(3) => B(35), B(2) =>
                           B(34), B(1) => B(33), B(0) => B(32), C_sel => 
                           C_in(8), S(3) => S(35), S(2) => S(34), S(1) => S(33)
                           , S(0) => S(32));
   csb_9 : carry_select_block_n4_23 port map( A(3) => A(39), A(2) => A(38), 
                           A(1) => A(37), A(0) => A(36), B(3) => B(39), B(2) =>
                           B(38), B(1) => B(37), B(0) => B(36), C_sel => 
                           C_in(9), S(3) => S(39), S(2) => S(38), S(1) => S(37)
                           , S(0) => S(36));
   csb_10 : carry_select_block_n4_22 port map( A(3) => A(43), A(2) => A(42), 
                           A(1) => A(41), A(0) => A(40), B(3) => B(43), B(2) =>
                           B(42), B(1) => B(41), B(0) => B(40), C_sel => 
                           C_in(10), S(3) => S(43), S(2) => S(42), S(1) => 
                           S(41), S(0) => S(40));
   csb_11 : carry_select_block_n4_21 port map( A(3) => A(47), A(2) => A(46), 
                           A(1) => A(45), A(0) => A(44), B(3) => B(47), B(2) =>
                           B(46), B(1) => B(45), B(0) => B(44), C_sel => 
                           C_in(11), S(3) => S(47), S(2) => S(46), S(1) => 
                           S(45), S(0) => S(44));
   csb_12 : carry_select_block_n4_20 port map( A(3) => A(51), A(2) => A(50), 
                           A(1) => A(49), A(0) => A(48), B(3) => B(51), B(2) =>
                           B(50), B(1) => B(49), B(0) => B(48), C_sel => 
                           C_in(12), S(3) => S(51), S(2) => S(50), S(1) => 
                           S(49), S(0) => S(48));
   csb_13 : carry_select_block_n4_19 port map( A(3) => A(55), A(2) => A(54), 
                           A(1) => A(53), A(0) => A(52), B(3) => B(55), B(2) =>
                           B(54), B(1) => B(53), B(0) => B(52), C_sel => 
                           C_in(13), S(3) => S(55), S(2) => S(54), S(1) => 
                           S(53), S(0) => S(52));
   csb_14 : carry_select_block_n4_18 port map( A(3) => A(59), A(2) => A(58), 
                           A(1) => A(57), A(0) => A(56), B(3) => B(59), B(2) =>
                           B(58), B(1) => B(57), B(0) => B(56), C_sel => 
                           C_in(14), S(3) => S(59), S(2) => S(58), S(1) => 
                           S(57), S(0) => S(56));
   csb_15 : carry_select_block_n4_17 port map( A(3) => A(63), A(2) => A(62), 
                           A(1) => A(61), A(0) => A(60), B(3) => B(63), B(2) =>
                           B(62), B(1) => B(61), B(0) => B(60), C_sel => 
                           C_in(15), S(3) => S(63), S(2) => S(62), S(1) => 
                           S(61), S(0) => S(60));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity sum_generator_n_bit64_n_CSB16_1 is

   port( A, B : in std_logic_vector (63 downto 0);  C_in : in std_logic_vector 
         (15 downto 0);  S : out std_logic_vector (63 downto 0));

end sum_generator_n_bit64_n_CSB16_1;

architecture SYN_STRUCTURAL of sum_generator_n_bit64_n_CSB16_1 is

   component carry_select_block_n4_1
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_n4_2
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_n4_3
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_n4_4
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_n4_5
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_n4_6
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_n4_7
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_n4_8
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_n4_9
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_n4_10
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_n4_11
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_n4_12
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_n4_13
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_n4_14
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_n4_15
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_n4_16
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;

begin
   
   csb_0 : carry_select_block_n4_16 port map( A(3) => A(3), A(2) => A(2), A(1) 
                           => A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), 
                           B(1) => B(1), B(0) => B(0), C_sel => C_in(0), S(3) 
                           => S(3), S(2) => S(2), S(1) => S(1), S(0) => S(0));
   csb_1 : carry_select_block_n4_15 port map( A(3) => A(7), A(2) => A(6), A(1) 
                           => A(5), A(0) => A(4), B(3) => B(7), B(2) => B(6), 
                           B(1) => B(5), B(0) => B(4), C_sel => C_in(1), S(3) 
                           => S(7), S(2) => S(6), S(1) => S(5), S(0) => S(4));
   csb_2 : carry_select_block_n4_14 port map( A(3) => A(11), A(2) => A(10), 
                           A(1) => A(9), A(0) => A(8), B(3) => B(11), B(2) => 
                           B(10), B(1) => B(9), B(0) => B(8), C_sel => C_in(2),
                           S(3) => S(11), S(2) => S(10), S(1) => S(9), S(0) => 
                           S(8));
   csb_3 : carry_select_block_n4_13 port map( A(3) => A(15), A(2) => A(14), 
                           A(1) => A(13), A(0) => A(12), B(3) => B(15), B(2) =>
                           B(14), B(1) => B(13), B(0) => B(12), C_sel => 
                           C_in(3), S(3) => S(15), S(2) => S(14), S(1) => S(13)
                           , S(0) => S(12));
   csb_4 : carry_select_block_n4_12 port map( A(3) => A(19), A(2) => A(18), 
                           A(1) => A(17), A(0) => A(16), B(3) => B(19), B(2) =>
                           B(18), B(1) => B(17), B(0) => B(16), C_sel => 
                           C_in(4), S(3) => S(19), S(2) => S(18), S(1) => S(17)
                           , S(0) => S(16));
   csb_5 : carry_select_block_n4_11 port map( A(3) => A(23), A(2) => A(22), 
                           A(1) => A(21), A(0) => A(20), B(3) => B(23), B(2) =>
                           B(22), B(1) => B(21), B(0) => B(20), C_sel => 
                           C_in(5), S(3) => S(23), S(2) => S(22), S(1) => S(21)
                           , S(0) => S(20));
   csb_6 : carry_select_block_n4_10 port map( A(3) => A(27), A(2) => A(26), 
                           A(1) => A(25), A(0) => A(24), B(3) => B(27), B(2) =>
                           B(26), B(1) => B(25), B(0) => B(24), C_sel => 
                           C_in(6), S(3) => S(27), S(2) => S(26), S(1) => S(25)
                           , S(0) => S(24));
   csb_7 : carry_select_block_n4_9 port map( A(3) => A(31), A(2) => A(30), A(1)
                           => A(29), A(0) => A(28), B(3) => B(31), B(2) => 
                           B(30), B(1) => B(29), B(0) => B(28), C_sel => 
                           C_in(7), S(3) => S(31), S(2) => S(30), S(1) => S(29)
                           , S(0) => S(28));
   csb_8 : carry_select_block_n4_8 port map( A(3) => A(35), A(2) => A(34), A(1)
                           => A(33), A(0) => A(32), B(3) => B(35), B(2) => 
                           B(34), B(1) => B(33), B(0) => B(32), C_sel => 
                           C_in(8), S(3) => S(35), S(2) => S(34), S(1) => S(33)
                           , S(0) => S(32));
   csb_9 : carry_select_block_n4_7 port map( A(3) => A(39), A(2) => A(38), A(1)
                           => A(37), A(0) => A(36), B(3) => B(39), B(2) => 
                           B(38), B(1) => B(37), B(0) => B(36), C_sel => 
                           C_in(9), S(3) => S(39), S(2) => S(38), S(1) => S(37)
                           , S(0) => S(36));
   csb_10 : carry_select_block_n4_6 port map( A(3) => A(43), A(2) => A(42), 
                           A(1) => A(41), A(0) => A(40), B(3) => B(43), B(2) =>
                           B(42), B(1) => B(41), B(0) => B(40), C_sel => 
                           C_in(10), S(3) => S(43), S(2) => S(42), S(1) => 
                           S(41), S(0) => S(40));
   csb_11 : carry_select_block_n4_5 port map( A(3) => A(47), A(2) => A(46), 
                           A(1) => A(45), A(0) => A(44), B(3) => B(47), B(2) =>
                           B(46), B(1) => B(45), B(0) => B(44), C_sel => 
                           C_in(11), S(3) => S(47), S(2) => S(46), S(1) => 
                           S(45), S(0) => S(44));
   csb_12 : carry_select_block_n4_4 port map( A(3) => A(51), A(2) => A(50), 
                           A(1) => A(49), A(0) => A(48), B(3) => B(51), B(2) =>
                           B(50), B(1) => B(49), B(0) => B(48), C_sel => 
                           C_in(12), S(3) => S(51), S(2) => S(50), S(1) => 
                           S(49), S(0) => S(48));
   csb_13 : carry_select_block_n4_3 port map( A(3) => A(55), A(2) => A(54), 
                           A(1) => A(53), A(0) => A(52), B(3) => B(55), B(2) =>
                           B(54), B(1) => B(53), B(0) => B(52), C_sel => 
                           C_in(13), S(3) => S(55), S(2) => S(54), S(1) => 
                           S(53), S(0) => S(52));
   csb_14 : carry_select_block_n4_2 port map( A(3) => A(59), A(2) => A(58), 
                           A(1) => A(57), A(0) => A(56), B(3) => B(59), B(2) =>
                           B(58), B(1) => B(57), B(0) => B(56), C_sel => 
                           C_in(14), S(3) => S(59), S(2) => S(58), S(1) => 
                           S(57), S(0) => S(56));
   csb_15 : carry_select_block_n4_1 port map( A(3) => A(63), A(2) => A(62), 
                           A(1) => A(61), A(0) => A(60), B(3) => B(63), B(2) =>
                           B(62), B(1) => B(61), B(0) => B(60), C_sel => 
                           C_in(15), S(3) => S(63), S(2) => S(62), S(1) => 
                           S(61), S(0) => S(60));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity CARRY_GENERATOR_NBIT64_NBIT_PER_BLOCK4_2 is

   port( A, B : in std_logic_vector (63 downto 0);  Cin : in std_logic;  Co : 
         out std_logic_vector (15 downto 0));

end CARRY_GENERATOR_NBIT64_NBIT_PER_BLOCK4_2;

architecture SYN_structural of CARRY_GENERATOR_NBIT64_NBIT_PER_BLOCK4_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component G_BLOCK_18
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component G_BLOCK_19
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component G_BLOCK_20
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component G_BLOCK_21
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component G_BLOCK_22
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component G_BLOCK_23
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component G_BLOCK_24
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component G_BLOCK_25
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component G_BLOCK_26
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component G_BLOCK_27
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component G_BLOCK_28
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component G_BLOCK_29
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component PG_BLOCK_64
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_65
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_66
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_67
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component G_BLOCK_30
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component G_BLOCK_31
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component PG_BLOCK_68
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_69
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_70
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_71
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_72
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_73
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component G_BLOCK_32
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component PG_BLOCK_74
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_75
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_76
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_77
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_78
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_79
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_80
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component G_BLOCK_33
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component PG_BLOCK_81
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_82
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_83
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_84
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_85
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_86
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_87
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_88
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_89
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_90
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_91
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_92
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_93
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_94
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_95
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component G_BLOCK_34
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component PG_BLOCK_96
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_97
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_98
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_99
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_100
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_101
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_102
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_103
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_104
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_105
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_106
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_107
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_108
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_109
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_110
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_111
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_112
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_113
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_114
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_115
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_116
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_117
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_118
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_119
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_120
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_121
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_122
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_123
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_124
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_125
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_126
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component pg_net_64
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_65
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_66
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_67
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_68
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_69
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_70
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_71
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_72
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_73
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_74
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_75
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_76
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_77
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_78
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_79
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_80
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_81
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_82
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_83
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_84
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_85
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_86
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_87
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_88
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_89
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_90
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_91
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_92
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_93
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_94
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_95
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_96
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_97
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_98
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_99
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_100
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_101
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_102
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_103
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_104
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_105
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_106
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_107
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_108
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_109
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_110
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_111
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_112
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_113
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_114
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_115
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_116
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_117
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_118
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_119
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_120
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_121
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_122
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_123
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_124
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_125
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_126
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   signal Co_15_port, Co_14_port, Co_13_port, Co_12_port, Co_11_port, 
      Co_10_port, Co_9_port, Co_8_port, Co_7_port, Co_6_port, Co_5_port, 
      Co_4_port, Co_3_port, Co_2_port, Co_1_port, Co_0_port, g_vector_5_63_port
      , g_vector_5_59_port, g_vector_5_55_port, g_vector_5_51_port, 
      g_vector_4_63_port, g_vector_4_59_port, g_vector_4_47_port, 
      g_vector_4_43_port, g_vector_4_31_port, g_vector_4_27_port, 
      g_vector_3_63_port, g_vector_3_55_port, g_vector_3_47_port, 
      g_vector_3_39_port, g_vector_3_31_port, g_vector_3_23_port, 
      g_vector_3_15_port, g_vector_2_63_port, g_vector_2_59_port, 
      g_vector_2_55_port, g_vector_2_51_port, g_vector_2_47_port, 
      g_vector_2_43_port, g_vector_2_39_port, g_vector_2_35_port, 
      g_vector_2_31_port, g_vector_2_27_port, g_vector_2_23_port, 
      g_vector_2_19_port, g_vector_2_15_port, g_vector_2_11_port, 
      g_vector_2_7_port, g_vector_1_63_port, g_vector_1_61_port, 
      g_vector_1_59_port, g_vector_1_57_port, g_vector_1_55_port, 
      g_vector_1_53_port, g_vector_1_51_port, g_vector_1_49_port, 
      g_vector_1_47_port, g_vector_1_45_port, g_vector_1_43_port, 
      g_vector_1_41_port, g_vector_1_39_port, g_vector_1_37_port, 
      g_vector_1_35_port, g_vector_1_33_port, g_vector_1_31_port, 
      g_vector_1_29_port, g_vector_1_27_port, g_vector_1_25_port, 
      g_vector_1_23_port, g_vector_1_21_port, g_vector_1_19_port, 
      g_vector_1_17_port, g_vector_1_15_port, g_vector_1_13_port, 
      g_vector_1_11_port, g_vector_1_9_port, g_vector_1_7_port, 
      g_vector_1_5_port, g_vector_1_3_port, g_vector_1_1_port, 
      g_vector_0_63_port, g_vector_0_62_port, g_vector_0_61_port, 
      g_vector_0_60_port, g_vector_0_59_port, g_vector_0_58_port, 
      g_vector_0_57_port, g_vector_0_56_port, g_vector_0_55_port, 
      g_vector_0_54_port, g_vector_0_53_port, g_vector_0_52_port, 
      g_vector_0_51_port, g_vector_0_50_port, g_vector_0_49_port, 
      g_vector_0_48_port, g_vector_0_47_port, g_vector_0_46_port, 
      g_vector_0_45_port, g_vector_0_44_port, g_vector_0_43_port, 
      g_vector_0_42_port, g_vector_0_41_port, g_vector_0_40_port, 
      g_vector_0_39_port, g_vector_0_38_port, g_vector_0_37_port, 
      g_vector_0_36_port, g_vector_0_35_port, g_vector_0_34_port, 
      g_vector_0_33_port, g_vector_0_32_port, g_vector_0_31_port, 
      g_vector_0_30_port, g_vector_0_29_port, g_vector_0_28_port, 
      g_vector_0_27_port, g_vector_0_26_port, g_vector_0_25_port, 
      g_vector_0_24_port, g_vector_0_23_port, g_vector_0_22_port, 
      g_vector_0_21_port, g_vector_0_20_port, g_vector_0_19_port, 
      g_vector_0_18_port, g_vector_0_17_port, g_vector_0_16_port, 
      g_vector_0_15_port, g_vector_0_14_port, g_vector_0_13_port, 
      g_vector_0_12_port, g_vector_0_11_port, g_vector_0_10_port, 
      g_vector_0_9_port, g_vector_0_8_port, g_vector_0_7_port, 
      g_vector_0_6_port, g_vector_0_5_port, g_vector_0_4_port, 
      g_vector_0_3_port, g_vector_0_2_port, g_vector_0_1_port, 
      g_vector_0_0_port, p_vector_5_63_port, p_vector_5_59_port, 
      p_vector_5_55_port, p_vector_5_51_port, p_vector_4_63_port, 
      p_vector_4_59_port, p_vector_4_47_port, p_vector_4_43_port, 
      p_vector_4_31_port, p_vector_4_27_port, p_vector_3_63_port, 
      p_vector_3_55_port, p_vector_3_47_port, p_vector_3_39_port, 
      p_vector_3_31_port, p_vector_3_23_port, p_vector_3_15_port, 
      p_vector_2_63_port, p_vector_2_59_port, p_vector_2_55_port, 
      p_vector_2_51_port, p_vector_2_47_port, p_vector_2_43_port, 
      p_vector_2_39_port, p_vector_2_35_port, p_vector_2_31_port, 
      p_vector_2_27_port, p_vector_2_23_port, p_vector_2_19_port, 
      p_vector_2_15_port, p_vector_2_11_port, p_vector_2_7_port, 
      p_vector_1_63_port, p_vector_1_61_port, p_vector_1_59_port, 
      p_vector_1_57_port, p_vector_1_55_port, p_vector_1_53_port, 
      p_vector_1_51_port, p_vector_1_49_port, p_vector_1_47_port, 
      p_vector_1_45_port, p_vector_1_43_port, p_vector_1_41_port, 
      p_vector_1_39_port, p_vector_1_37_port, p_vector_1_35_port, 
      p_vector_1_33_port, p_vector_1_31_port, p_vector_1_29_port, 
      p_vector_1_27_port, p_vector_1_25_port, p_vector_1_23_port, 
      p_vector_1_21_port, p_vector_1_19_port, p_vector_1_17_port, 
      p_vector_1_15_port, p_vector_1_13_port, p_vector_1_11_port, 
      p_vector_1_9_port, p_vector_1_7_port, p_vector_1_5_port, 
      p_vector_1_3_port, p_vector_0_63_port, p_vector_0_62_port, 
      p_vector_0_61_port, p_vector_0_60_port, p_vector_0_59_port, 
      p_vector_0_58_port, p_vector_0_57_port, p_vector_0_56_port, 
      p_vector_0_55_port, p_vector_0_54_port, p_vector_0_53_port, 
      p_vector_0_52_port, p_vector_0_51_port, p_vector_0_50_port, 
      p_vector_0_49_port, p_vector_0_48_port, p_vector_0_47_port, 
      p_vector_0_46_port, p_vector_0_45_port, p_vector_0_44_port, 
      p_vector_0_43_port, p_vector_0_42_port, p_vector_0_41_port, 
      p_vector_0_40_port, p_vector_0_39_port, p_vector_0_38_port, 
      p_vector_0_37_port, p_vector_0_36_port, p_vector_0_35_port, 
      p_vector_0_34_port, p_vector_0_33_port, p_vector_0_32_port, 
      p_vector_0_31_port, p_vector_0_30_port, p_vector_0_29_port, 
      p_vector_0_28_port, p_vector_0_27_port, p_vector_0_26_port, 
      p_vector_0_25_port, p_vector_0_24_port, p_vector_0_23_port, 
      p_vector_0_22_port, p_vector_0_21_port, p_vector_0_20_port, 
      p_vector_0_19_port, p_vector_0_18_port, p_vector_0_17_port, 
      p_vector_0_16_port, p_vector_0_15_port, p_vector_0_14_port, 
      p_vector_0_13_port, p_vector_0_12_port, p_vector_0_11_port, 
      p_vector_0_10_port, p_vector_0_9_port, p_vector_0_8_port, 
      p_vector_0_7_port, p_vector_0_6_port, p_vector_0_5_port, 
      p_vector_0_4_port, p_vector_0_3_port, p_vector_0_2_port, 
      p_vector_0_1_port, n1, n2, n4 : std_logic;

begin
   Co <= ( Co_15_port, Co_14_port, Co_13_port, Co_12_port, Co_11_port, 
      Co_10_port, Co_9_port, Co_8_port, Co_7_port, Co_6_port, Co_5_port, 
      Co_4_port, Co_3_port, Co_2_port, Co_1_port, Co_0_port );
   
   pg_network_63 : pg_net_126 port map( a => A(63), b => B(63), p => 
                           p_vector_0_63_port, g => g_vector_0_63_port);
   pg_network_62 : pg_net_125 port map( a => A(62), b => B(62), p => 
                           p_vector_0_62_port, g => g_vector_0_62_port);
   pg_network_61 : pg_net_124 port map( a => A(61), b => B(61), p => 
                           p_vector_0_61_port, g => g_vector_0_61_port);
   pg_network_60 : pg_net_123 port map( a => A(60), b => B(60), p => 
                           p_vector_0_60_port, g => g_vector_0_60_port);
   pg_network_59 : pg_net_122 port map( a => A(59), b => B(59), p => 
                           p_vector_0_59_port, g => g_vector_0_59_port);
   pg_network_58 : pg_net_121 port map( a => A(58), b => B(58), p => 
                           p_vector_0_58_port, g => g_vector_0_58_port);
   pg_network_57 : pg_net_120 port map( a => A(57), b => B(57), p => 
                           p_vector_0_57_port, g => g_vector_0_57_port);
   pg_network_56 : pg_net_119 port map( a => A(56), b => B(56), p => 
                           p_vector_0_56_port, g => g_vector_0_56_port);
   pg_network_55 : pg_net_118 port map( a => A(55), b => B(55), p => 
                           p_vector_0_55_port, g => g_vector_0_55_port);
   pg_network_54 : pg_net_117 port map( a => A(54), b => B(54), p => 
                           p_vector_0_54_port, g => g_vector_0_54_port);
   pg_network_53 : pg_net_116 port map( a => A(53), b => B(53), p => 
                           p_vector_0_53_port, g => g_vector_0_53_port);
   pg_network_52 : pg_net_115 port map( a => A(52), b => B(52), p => 
                           p_vector_0_52_port, g => g_vector_0_52_port);
   pg_network_51 : pg_net_114 port map( a => A(51), b => B(51), p => 
                           p_vector_0_51_port, g => g_vector_0_51_port);
   pg_network_50 : pg_net_113 port map( a => A(50), b => B(50), p => 
                           p_vector_0_50_port, g => g_vector_0_50_port);
   pg_network_49 : pg_net_112 port map( a => A(49), b => B(49), p => 
                           p_vector_0_49_port, g => g_vector_0_49_port);
   pg_network_48 : pg_net_111 port map( a => A(48), b => B(48), p => 
                           p_vector_0_48_port, g => g_vector_0_48_port);
   pg_network_47 : pg_net_110 port map( a => A(47), b => B(47), p => 
                           p_vector_0_47_port, g => g_vector_0_47_port);
   pg_network_46 : pg_net_109 port map( a => A(46), b => B(46), p => 
                           p_vector_0_46_port, g => g_vector_0_46_port);
   pg_network_45 : pg_net_108 port map( a => A(45), b => B(45), p => 
                           p_vector_0_45_port, g => g_vector_0_45_port);
   pg_network_44 : pg_net_107 port map( a => A(44), b => B(44), p => 
                           p_vector_0_44_port, g => g_vector_0_44_port);
   pg_network_43 : pg_net_106 port map( a => A(43), b => B(43), p => 
                           p_vector_0_43_port, g => g_vector_0_43_port);
   pg_network_42 : pg_net_105 port map( a => A(42), b => B(42), p => 
                           p_vector_0_42_port, g => g_vector_0_42_port);
   pg_network_41 : pg_net_104 port map( a => A(41), b => B(41), p => 
                           p_vector_0_41_port, g => g_vector_0_41_port);
   pg_network_40 : pg_net_103 port map( a => A(40), b => B(40), p => 
                           p_vector_0_40_port, g => g_vector_0_40_port);
   pg_network_39 : pg_net_102 port map( a => A(39), b => B(39), p => 
                           p_vector_0_39_port, g => g_vector_0_39_port);
   pg_network_38 : pg_net_101 port map( a => A(38), b => B(38), p => 
                           p_vector_0_38_port, g => g_vector_0_38_port);
   pg_network_37 : pg_net_100 port map( a => A(37), b => B(37), p => 
                           p_vector_0_37_port, g => g_vector_0_37_port);
   pg_network_36 : pg_net_99 port map( a => A(36), b => B(36), p => 
                           p_vector_0_36_port, g => g_vector_0_36_port);
   pg_network_35 : pg_net_98 port map( a => A(35), b => B(35), p => 
                           p_vector_0_35_port, g => g_vector_0_35_port);
   pg_network_34 : pg_net_97 port map( a => A(34), b => B(34), p => 
                           p_vector_0_34_port, g => g_vector_0_34_port);
   pg_network_33 : pg_net_96 port map( a => A(33), b => B(33), p => 
                           p_vector_0_33_port, g => g_vector_0_33_port);
   pg_network_32 : pg_net_95 port map( a => A(32), b => B(32), p => 
                           p_vector_0_32_port, g => g_vector_0_32_port);
   pg_network_31 : pg_net_94 port map( a => A(31), b => B(31), p => 
                           p_vector_0_31_port, g => g_vector_0_31_port);
   pg_network_30 : pg_net_93 port map( a => A(30), b => B(30), p => 
                           p_vector_0_30_port, g => g_vector_0_30_port);
   pg_network_29 : pg_net_92 port map( a => A(29), b => B(29), p => 
                           p_vector_0_29_port, g => g_vector_0_29_port);
   pg_network_28 : pg_net_91 port map( a => A(28), b => B(28), p => 
                           p_vector_0_28_port, g => g_vector_0_28_port);
   pg_network_27 : pg_net_90 port map( a => A(27), b => B(27), p => 
                           p_vector_0_27_port, g => g_vector_0_27_port);
   pg_network_26 : pg_net_89 port map( a => A(26), b => B(26), p => 
                           p_vector_0_26_port, g => g_vector_0_26_port);
   pg_network_25 : pg_net_88 port map( a => A(25), b => B(25), p => 
                           p_vector_0_25_port, g => g_vector_0_25_port);
   pg_network_24 : pg_net_87 port map( a => A(24), b => B(24), p => 
                           p_vector_0_24_port, g => g_vector_0_24_port);
   pg_network_23 : pg_net_86 port map( a => A(23), b => B(23), p => 
                           p_vector_0_23_port, g => g_vector_0_23_port);
   pg_network_22 : pg_net_85 port map( a => A(22), b => B(22), p => 
                           p_vector_0_22_port, g => g_vector_0_22_port);
   pg_network_21 : pg_net_84 port map( a => A(21), b => B(21), p => 
                           p_vector_0_21_port, g => g_vector_0_21_port);
   pg_network_20 : pg_net_83 port map( a => A(20), b => B(20), p => 
                           p_vector_0_20_port, g => g_vector_0_20_port);
   pg_network_19 : pg_net_82 port map( a => A(19), b => B(19), p => 
                           p_vector_0_19_port, g => g_vector_0_19_port);
   pg_network_18 : pg_net_81 port map( a => A(18), b => B(18), p => 
                           p_vector_0_18_port, g => g_vector_0_18_port);
   pg_network_17 : pg_net_80 port map( a => A(17), b => B(17), p => 
                           p_vector_0_17_port, g => g_vector_0_17_port);
   pg_network_16 : pg_net_79 port map( a => A(16), b => B(16), p => 
                           p_vector_0_16_port, g => g_vector_0_16_port);
   pg_network_15 : pg_net_78 port map( a => A(15), b => B(15), p => 
                           p_vector_0_15_port, g => g_vector_0_15_port);
   pg_network_14 : pg_net_77 port map( a => A(14), b => B(14), p => 
                           p_vector_0_14_port, g => g_vector_0_14_port);
   pg_network_13 : pg_net_76 port map( a => A(13), b => B(13), p => 
                           p_vector_0_13_port, g => g_vector_0_13_port);
   pg_network_12 : pg_net_75 port map( a => A(12), b => B(12), p => 
                           p_vector_0_12_port, g => g_vector_0_12_port);
   pg_network_11 : pg_net_74 port map( a => A(11), b => B(11), p => 
                           p_vector_0_11_port, g => g_vector_0_11_port);
   pg_network_10 : pg_net_73 port map( a => A(10), b => B(10), p => 
                           p_vector_0_10_port, g => g_vector_0_10_port);
   pg_network_9 : pg_net_72 port map( a => A(9), b => B(9), p => 
                           p_vector_0_9_port, g => g_vector_0_9_port);
   pg_network_8 : pg_net_71 port map( a => A(8), b => B(8), p => 
                           p_vector_0_8_port, g => g_vector_0_8_port);
   pg_network_7 : pg_net_70 port map( a => A(7), b => B(7), p => 
                           p_vector_0_7_port, g => g_vector_0_7_port);
   pg_network_6 : pg_net_69 port map( a => A(6), b => B(6), p => 
                           p_vector_0_6_port, g => g_vector_0_6_port);
   pg_network_5 : pg_net_68 port map( a => A(5), b => B(5), p => 
                           p_vector_0_5_port, g => g_vector_0_5_port);
   pg_network_4 : pg_net_67 port map( a => A(4), b => B(4), p => 
                           p_vector_0_4_port, g => g_vector_0_4_port);
   pg_network_3 : pg_net_66 port map( a => A(3), b => B(3), p => 
                           p_vector_0_3_port, g => g_vector_0_3_port);
   pg_network_2 : pg_net_65 port map( a => A(2), b => B(2), p => 
                           p_vector_0_2_port, g => g_vector_0_2_port);
   pg_network_1 : pg_net_64 port map( a => A(1), b => B(1), p => 
                           p_vector_0_1_port, g => g_vector_0_1_port);
   std_PG_1_63 : PG_BLOCK_126 port map( p2 => p_vector_0_63_port, g2 => 
                           g_vector_0_63_port, p1 => p_vector_0_62_port, g1 => 
                           g_vector_0_62_port, PG_P => p_vector_1_63_port, PG_G
                           => g_vector_1_63_port);
   std_PG_1_61 : PG_BLOCK_125 port map( p2 => p_vector_0_61_port, g2 => 
                           g_vector_0_61_port, p1 => p_vector_0_60_port, g1 => 
                           g_vector_0_60_port, PG_P => p_vector_1_61_port, PG_G
                           => g_vector_1_61_port);
   std_PG_1_59 : PG_BLOCK_124 port map( p2 => p_vector_0_59_port, g2 => 
                           g_vector_0_59_port, p1 => p_vector_0_58_port, g1 => 
                           g_vector_0_58_port, PG_P => p_vector_1_59_port, PG_G
                           => g_vector_1_59_port);
   std_PG_1_57 : PG_BLOCK_123 port map( p2 => p_vector_0_57_port, g2 => 
                           g_vector_0_57_port, p1 => p_vector_0_56_port, g1 => 
                           g_vector_0_56_port, PG_P => p_vector_1_57_port, PG_G
                           => g_vector_1_57_port);
   std_PG_1_55 : PG_BLOCK_122 port map( p2 => p_vector_0_55_port, g2 => 
                           g_vector_0_55_port, p1 => p_vector_0_54_port, g1 => 
                           g_vector_0_54_port, PG_P => p_vector_1_55_port, PG_G
                           => g_vector_1_55_port);
   std_PG_1_53 : PG_BLOCK_121 port map( p2 => p_vector_0_53_port, g2 => 
                           g_vector_0_53_port, p1 => p_vector_0_52_port, g1 => 
                           g_vector_0_52_port, PG_P => p_vector_1_53_port, PG_G
                           => g_vector_1_53_port);
   std_PG_1_51 : PG_BLOCK_120 port map( p2 => p_vector_0_51_port, g2 => 
                           g_vector_0_51_port, p1 => p_vector_0_50_port, g1 => 
                           g_vector_0_50_port, PG_P => p_vector_1_51_port, PG_G
                           => g_vector_1_51_port);
   std_PG_1_49 : PG_BLOCK_119 port map( p2 => p_vector_0_49_port, g2 => 
                           g_vector_0_49_port, p1 => p_vector_0_48_port, g1 => 
                           g_vector_0_48_port, PG_P => p_vector_1_49_port, PG_G
                           => g_vector_1_49_port);
   std_PG_1_47 : PG_BLOCK_118 port map( p2 => p_vector_0_47_port, g2 => 
                           g_vector_0_47_port, p1 => p_vector_0_46_port, g1 => 
                           g_vector_0_46_port, PG_P => p_vector_1_47_port, PG_G
                           => g_vector_1_47_port);
   std_PG_1_45 : PG_BLOCK_117 port map( p2 => p_vector_0_45_port, g2 => 
                           g_vector_0_45_port, p1 => p_vector_0_44_port, g1 => 
                           g_vector_0_44_port, PG_P => p_vector_1_45_port, PG_G
                           => g_vector_1_45_port);
   std_PG_1_43 : PG_BLOCK_116 port map( p2 => p_vector_0_43_port, g2 => 
                           g_vector_0_43_port, p1 => p_vector_0_42_port, g1 => 
                           g_vector_0_42_port, PG_P => p_vector_1_43_port, PG_G
                           => g_vector_1_43_port);
   std_PG_1_41 : PG_BLOCK_115 port map( p2 => p_vector_0_41_port, g2 => 
                           g_vector_0_41_port, p1 => p_vector_0_40_port, g1 => 
                           g_vector_0_40_port, PG_P => p_vector_1_41_port, PG_G
                           => g_vector_1_41_port);
   std_PG_1_39 : PG_BLOCK_114 port map( p2 => p_vector_0_39_port, g2 => 
                           g_vector_0_39_port, p1 => p_vector_0_38_port, g1 => 
                           g_vector_0_38_port, PG_P => p_vector_1_39_port, PG_G
                           => g_vector_1_39_port);
   std_PG_1_37 : PG_BLOCK_113 port map( p2 => p_vector_0_37_port, g2 => 
                           g_vector_0_37_port, p1 => p_vector_0_36_port, g1 => 
                           g_vector_0_36_port, PG_P => p_vector_1_37_port, PG_G
                           => g_vector_1_37_port);
   std_PG_1_35 : PG_BLOCK_112 port map( p2 => p_vector_0_35_port, g2 => 
                           g_vector_0_35_port, p1 => p_vector_0_34_port, g1 => 
                           g_vector_0_34_port, PG_P => p_vector_1_35_port, PG_G
                           => g_vector_1_35_port);
   std_PG_1_33 : PG_BLOCK_111 port map( p2 => p_vector_0_33_port, g2 => 
                           g_vector_0_33_port, p1 => p_vector_0_32_port, g1 => 
                           g_vector_0_32_port, PG_P => p_vector_1_33_port, PG_G
                           => g_vector_1_33_port);
   std_PG_1_31 : PG_BLOCK_110 port map( p2 => p_vector_0_31_port, g2 => 
                           g_vector_0_31_port, p1 => p_vector_0_30_port, g1 => 
                           g_vector_0_30_port, PG_P => p_vector_1_31_port, PG_G
                           => g_vector_1_31_port);
   std_PG_1_29 : PG_BLOCK_109 port map( p2 => p_vector_0_29_port, g2 => 
                           g_vector_0_29_port, p1 => p_vector_0_28_port, g1 => 
                           g_vector_0_28_port, PG_P => p_vector_1_29_port, PG_G
                           => g_vector_1_29_port);
   std_PG_1_27 : PG_BLOCK_108 port map( p2 => p_vector_0_27_port, g2 => 
                           g_vector_0_27_port, p1 => p_vector_0_26_port, g1 => 
                           g_vector_0_26_port, PG_P => p_vector_1_27_port, PG_G
                           => g_vector_1_27_port);
   std_PG_1_25 : PG_BLOCK_107 port map( p2 => p_vector_0_25_port, g2 => 
                           g_vector_0_25_port, p1 => p_vector_0_24_port, g1 => 
                           g_vector_0_24_port, PG_P => p_vector_1_25_port, PG_G
                           => g_vector_1_25_port);
   std_PG_1_23 : PG_BLOCK_106 port map( p2 => p_vector_0_23_port, g2 => 
                           g_vector_0_23_port, p1 => p_vector_0_22_port, g1 => 
                           g_vector_0_22_port, PG_P => p_vector_1_23_port, PG_G
                           => g_vector_1_23_port);
   std_PG_1_21 : PG_BLOCK_105 port map( p2 => p_vector_0_21_port, g2 => 
                           g_vector_0_21_port, p1 => p_vector_0_20_port, g1 => 
                           g_vector_0_20_port, PG_P => p_vector_1_21_port, PG_G
                           => g_vector_1_21_port);
   std_PG_1_19 : PG_BLOCK_104 port map( p2 => p_vector_0_19_port, g2 => 
                           g_vector_0_19_port, p1 => p_vector_0_18_port, g1 => 
                           g_vector_0_18_port, PG_P => p_vector_1_19_port, PG_G
                           => g_vector_1_19_port);
   std_PG_1_17 : PG_BLOCK_103 port map( p2 => p_vector_0_17_port, g2 => 
                           g_vector_0_17_port, p1 => p_vector_0_16_port, g1 => 
                           g_vector_0_16_port, PG_P => p_vector_1_17_port, PG_G
                           => g_vector_1_17_port);
   std_PG_1_15 : PG_BLOCK_102 port map( p2 => p_vector_0_15_port, g2 => 
                           g_vector_0_15_port, p1 => p_vector_0_14_port, g1 => 
                           g_vector_0_14_port, PG_P => p_vector_1_15_port, PG_G
                           => g_vector_1_15_port);
   std_PG_1_13 : PG_BLOCK_101 port map( p2 => p_vector_0_13_port, g2 => 
                           g_vector_0_13_port, p1 => p_vector_0_12_port, g1 => 
                           g_vector_0_12_port, PG_P => p_vector_1_13_port, PG_G
                           => g_vector_1_13_port);
   std_PG_1_11 : PG_BLOCK_100 port map( p2 => p_vector_0_11_port, g2 => 
                           g_vector_0_11_port, p1 => p_vector_0_10_port, g1 => 
                           g_vector_0_10_port, PG_P => p_vector_1_11_port, PG_G
                           => g_vector_1_11_port);
   std_PG_1_9 : PG_BLOCK_99 port map( p2 => p_vector_0_9_port, g2 => 
                           g_vector_0_9_port, p1 => p_vector_0_8_port, g1 => 
                           g_vector_0_8_port, PG_P => p_vector_1_9_port, PG_G 
                           => g_vector_1_9_port);
   std_PG_1_7 : PG_BLOCK_98 port map( p2 => p_vector_0_7_port, g2 => 
                           g_vector_0_7_port, p1 => p_vector_0_6_port, g1 => 
                           g_vector_0_6_port, PG_P => p_vector_1_7_port, PG_G 
                           => g_vector_1_7_port);
   std_PG_1_5 : PG_BLOCK_97 port map( p2 => p_vector_0_5_port, g2 => 
                           g_vector_0_5_port, p1 => p_vector_0_4_port, g1 => 
                           g_vector_0_4_port, PG_P => p_vector_1_5_port, PG_G 
                           => g_vector_1_5_port);
   std_PG_1_3 : PG_BLOCK_96 port map( p2 => p_vector_0_3_port, g2 => 
                           g_vector_0_3_port, p1 => p_vector_0_2_port, g1 => 
                           g_vector_0_2_port, PG_P => p_vector_1_3_port, PG_G 
                           => g_vector_1_3_port);
   std_G_1_1 : G_BLOCK_34 port map( p2 => p_vector_0_1_port, g2 => 
                           g_vector_0_1_port, g1 => g_vector_0_0_port, G => 
                           g_vector_1_1_port);
   std_PG_2_63 : PG_BLOCK_95 port map( p2 => p_vector_1_63_port, g2 => 
                           g_vector_1_63_port, p1 => p_vector_1_61_port, g1 => 
                           g_vector_1_61_port, PG_P => p_vector_2_63_port, PG_G
                           => g_vector_2_63_port);
   std_PG_2_59 : PG_BLOCK_94 port map( p2 => p_vector_1_59_port, g2 => 
                           g_vector_1_59_port, p1 => p_vector_1_57_port, g1 => 
                           g_vector_1_57_port, PG_P => p_vector_2_59_port, PG_G
                           => g_vector_2_59_port);
   std_PG_2_55 : PG_BLOCK_93 port map( p2 => p_vector_1_55_port, g2 => 
                           g_vector_1_55_port, p1 => p_vector_1_53_port, g1 => 
                           g_vector_1_53_port, PG_P => p_vector_2_55_port, PG_G
                           => g_vector_2_55_port);
   std_PG_2_51 : PG_BLOCK_92 port map( p2 => p_vector_1_51_port, g2 => 
                           g_vector_1_51_port, p1 => p_vector_1_49_port, g1 => 
                           g_vector_1_49_port, PG_P => p_vector_2_51_port, PG_G
                           => g_vector_2_51_port);
   std_PG_2_47 : PG_BLOCK_91 port map( p2 => p_vector_1_47_port, g2 => 
                           g_vector_1_47_port, p1 => p_vector_1_45_port, g1 => 
                           g_vector_1_45_port, PG_P => p_vector_2_47_port, PG_G
                           => g_vector_2_47_port);
   std_PG_2_43 : PG_BLOCK_90 port map( p2 => p_vector_1_43_port, g2 => 
                           g_vector_1_43_port, p1 => p_vector_1_41_port, g1 => 
                           g_vector_1_41_port, PG_P => p_vector_2_43_port, PG_G
                           => g_vector_2_43_port);
   std_PG_2_39 : PG_BLOCK_89 port map( p2 => p_vector_1_39_port, g2 => 
                           g_vector_1_39_port, p1 => p_vector_1_37_port, g1 => 
                           g_vector_1_37_port, PG_P => p_vector_2_39_port, PG_G
                           => g_vector_2_39_port);
   std_PG_2_35 : PG_BLOCK_88 port map( p2 => p_vector_1_35_port, g2 => 
                           g_vector_1_35_port, p1 => p_vector_1_33_port, g1 => 
                           g_vector_1_33_port, PG_P => p_vector_2_35_port, PG_G
                           => g_vector_2_35_port);
   std_PG_2_31 : PG_BLOCK_87 port map( p2 => p_vector_1_31_port, g2 => 
                           g_vector_1_31_port, p1 => p_vector_1_29_port, g1 => 
                           g_vector_1_29_port, PG_P => p_vector_2_31_port, PG_G
                           => g_vector_2_31_port);
   std_PG_2_27 : PG_BLOCK_86 port map( p2 => p_vector_1_27_port, g2 => 
                           g_vector_1_27_port, p1 => p_vector_1_25_port, g1 => 
                           g_vector_1_25_port, PG_P => p_vector_2_27_port, PG_G
                           => g_vector_2_27_port);
   std_PG_2_23 : PG_BLOCK_85 port map( p2 => p_vector_1_23_port, g2 => 
                           g_vector_1_23_port, p1 => p_vector_1_21_port, g1 => 
                           g_vector_1_21_port, PG_P => p_vector_2_23_port, PG_G
                           => g_vector_2_23_port);
   std_PG_2_19 : PG_BLOCK_84 port map( p2 => p_vector_1_19_port, g2 => 
                           g_vector_1_19_port, p1 => p_vector_1_17_port, g1 => 
                           g_vector_1_17_port, PG_P => p_vector_2_19_port, PG_G
                           => g_vector_2_19_port);
   std_PG_2_15 : PG_BLOCK_83 port map( p2 => p_vector_1_15_port, g2 => 
                           g_vector_1_15_port, p1 => p_vector_1_13_port, g1 => 
                           g_vector_1_13_port, PG_P => p_vector_2_15_port, PG_G
                           => g_vector_2_15_port);
   std_PG_2_11 : PG_BLOCK_82 port map( p2 => p_vector_1_11_port, g2 => 
                           g_vector_1_11_port, p1 => p_vector_1_9_port, g1 => 
                           g_vector_1_9_port, PG_P => p_vector_2_11_port, PG_G 
                           => g_vector_2_11_port);
   std_PG_2_7 : PG_BLOCK_81 port map( p2 => p_vector_1_7_port, g2 => 
                           g_vector_1_7_port, p1 => p_vector_1_5_port, g1 => 
                           g_vector_1_5_port, PG_P => p_vector_2_7_port, PG_G 
                           => g_vector_2_7_port);
   std_G_2_3 : G_BLOCK_33 port map( p2 => p_vector_1_3_port, g2 => 
                           g_vector_1_3_port, g1 => g_vector_1_1_port, G => 
                           Co_0_port);
   std_PG_3_63 : PG_BLOCK_80 port map( p2 => p_vector_2_63_port, g2 => 
                           g_vector_2_63_port, p1 => p_vector_2_59_port, g1 => 
                           g_vector_2_59_port, PG_P => p_vector_3_63_port, PG_G
                           => g_vector_3_63_port);
   std_PG_3_55 : PG_BLOCK_79 port map( p2 => p_vector_2_55_port, g2 => 
                           g_vector_2_55_port, p1 => p_vector_2_51_port, g1 => 
                           g_vector_2_51_port, PG_P => p_vector_3_55_port, PG_G
                           => g_vector_3_55_port);
   std_PG_3_47 : PG_BLOCK_78 port map( p2 => p_vector_2_47_port, g2 => 
                           g_vector_2_47_port, p1 => p_vector_2_43_port, g1 => 
                           g_vector_2_43_port, PG_P => p_vector_3_47_port, PG_G
                           => g_vector_3_47_port);
   std_PG_3_39 : PG_BLOCK_77 port map( p2 => p_vector_2_39_port, g2 => 
                           g_vector_2_39_port, p1 => p_vector_2_35_port, g1 => 
                           g_vector_2_35_port, PG_P => p_vector_3_39_port, PG_G
                           => g_vector_3_39_port);
   std_PG_3_31 : PG_BLOCK_76 port map( p2 => p_vector_2_31_port, g2 => 
                           g_vector_2_31_port, p1 => p_vector_2_27_port, g1 => 
                           g_vector_2_27_port, PG_P => p_vector_3_31_port, PG_G
                           => g_vector_3_31_port);
   std_PG_3_23 : PG_BLOCK_75 port map( p2 => p_vector_2_23_port, g2 => 
                           g_vector_2_23_port, p1 => p_vector_2_19_port, g1 => 
                           g_vector_2_19_port, PG_P => p_vector_3_23_port, PG_G
                           => g_vector_3_23_port);
   std_PG_3_15 : PG_BLOCK_74 port map( p2 => p_vector_2_15_port, g2 => 
                           g_vector_2_15_port, p1 => p_vector_2_11_port, g1 => 
                           g_vector_2_11_port, PG_P => p_vector_3_15_port, PG_G
                           => g_vector_3_15_port);
   std_G_3_7 : G_BLOCK_32 port map( p2 => p_vector_2_7_port, g2 => 
                           g_vector_2_7_port, g1 => Co_0_port, G => Co_1_port);
   std_PG_4_63 : PG_BLOCK_73 port map( p2 => p_vector_3_63_port, g2 => 
                           g_vector_3_63_port, p1 => p_vector_3_55_port, g1 => 
                           g_vector_3_55_port, PG_P => p_vector_4_63_port, PG_G
                           => g_vector_4_63_port);
   add_PG_4_63_1 : PG_BLOCK_72 port map( p2 => p_vector_2_59_port, g2 => 
                           g_vector_2_59_port, p1 => p_vector_3_55_port, g1 => 
                           g_vector_3_55_port, PG_P => p_vector_4_59_port, PG_G
                           => g_vector_4_59_port);
   std_PG_4_47 : PG_BLOCK_71 port map( p2 => p_vector_3_47_port, g2 => 
                           g_vector_3_47_port, p1 => p_vector_3_39_port, g1 => 
                           g_vector_3_39_port, PG_P => p_vector_4_47_port, PG_G
                           => g_vector_4_47_port);
   add_PG_4_47_1 : PG_BLOCK_70 port map( p2 => p_vector_2_43_port, g2 => 
                           g_vector_2_43_port, p1 => p_vector_3_39_port, g1 => 
                           g_vector_3_39_port, PG_P => p_vector_4_43_port, PG_G
                           => g_vector_4_43_port);
   std_PG_4_31 : PG_BLOCK_69 port map( p2 => p_vector_3_31_port, g2 => 
                           g_vector_3_31_port, p1 => p_vector_3_23_port, g1 => 
                           g_vector_3_23_port, PG_P => p_vector_4_31_port, PG_G
                           => g_vector_4_31_port);
   add_PG_4_31_1 : PG_BLOCK_68 port map( p2 => p_vector_2_27_port, g2 => 
                           g_vector_2_27_port, p1 => p_vector_3_23_port, g1 => 
                           g_vector_3_23_port, PG_P => p_vector_4_27_port, PG_G
                           => g_vector_4_27_port);
   std_G_4_15 : G_BLOCK_31 port map( p2 => p_vector_3_15_port, g2 => 
                           g_vector_3_15_port, g1 => Co_1_port, G => Co_3_port)
                           ;
   add_G_4_15_1 : G_BLOCK_30 port map( p2 => p_vector_2_11_port, g2 => 
                           g_vector_2_11_port, g1 => Co_1_port, G => Co_2_port)
                           ;
   std_PG_5_63 : PG_BLOCK_67 port map( p2 => p_vector_4_63_port, g2 => 
                           g_vector_4_63_port, p1 => p_vector_4_47_port, g1 => 
                           g_vector_4_47_port, PG_P => p_vector_5_63_port, PG_G
                           => g_vector_5_63_port);
   add_PG_5_63_1 : PG_BLOCK_66 port map( p2 => p_vector_4_59_port, g2 => 
                           g_vector_4_59_port, p1 => p_vector_4_47_port, g1 => 
                           g_vector_4_47_port, PG_P => p_vector_5_59_port, PG_G
                           => g_vector_5_59_port);
   add_PG_5_63_2 : PG_BLOCK_65 port map( p2 => p_vector_3_55_port, g2 => 
                           g_vector_3_55_port, p1 => p_vector_4_47_port, g1 => 
                           g_vector_4_47_port, PG_P => p_vector_5_55_port, PG_G
                           => g_vector_5_55_port);
   add_PG_5_63_3 : PG_BLOCK_64 port map( p2 => p_vector_2_51_port, g2 => 
                           g_vector_2_51_port, p1 => p_vector_4_47_port, g1 => 
                           g_vector_4_47_port, PG_P => p_vector_5_51_port, PG_G
                           => g_vector_5_51_port);
   std_G_5_31 : G_BLOCK_29 port map( p2 => p_vector_4_31_port, g2 => 
                           g_vector_4_31_port, g1 => Co_3_port, G => Co_7_port)
                           ;
   add_G_5_31_1 : G_BLOCK_28 port map( p2 => p_vector_4_27_port, g2 => 
                           g_vector_4_27_port, g1 => Co_3_port, G => Co_6_port)
                           ;
   add_G_5_31_2 : G_BLOCK_27 port map( p2 => p_vector_3_23_port, g2 => 
                           g_vector_3_23_port, g1 => Co_3_port, G => Co_5_port)
                           ;
   add_G_5_31_3 : G_BLOCK_26 port map( p2 => p_vector_2_19_port, g2 => 
                           g_vector_2_19_port, g1 => Co_3_port, G => Co_4_port)
                           ;
   std_G_6_63 : G_BLOCK_25 port map( p2 => p_vector_5_63_port, g2 => 
                           g_vector_5_63_port, g1 => Co_7_port, G => Co_15_port
                           );
   add_G_6_63_1 : G_BLOCK_24 port map( p2 => p_vector_5_59_port, g2 => 
                           g_vector_5_59_port, g1 => Co_7_port, G => Co_14_port
                           );
   add_G_6_63_2 : G_BLOCK_23 port map( p2 => p_vector_5_55_port, g2 => 
                           g_vector_5_55_port, g1 => Co_7_port, G => Co_13_port
                           );
   add_G_6_63_3 : G_BLOCK_22 port map( p2 => p_vector_5_51_port, g2 => 
                           g_vector_5_51_port, g1 => Co_7_port, G => Co_12_port
                           );
   add_G_6_63_4 : G_BLOCK_21 port map( p2 => p_vector_4_47_port, g2 => 
                           g_vector_4_47_port, g1 => Co_7_port, G => Co_11_port
                           );
   add_G_6_63_5 : G_BLOCK_20 port map( p2 => p_vector_4_43_port, g2 => 
                           g_vector_4_43_port, g1 => Co_7_port, G => Co_10_port
                           );
   add_G_6_63_6 : G_BLOCK_19 port map( p2 => p_vector_3_39_port, g2 => 
                           g_vector_3_39_port, g1 => Co_7_port, G => Co_9_port)
                           ;
   add_G_6_63_7 : G_BLOCK_18 port map( p2 => p_vector_2_35_port, g2 => 
                           g_vector_2_35_port, g1 => Co_7_port, G => Co_8_port)
                           ;
   U1 : OAI21_X1 port map( B1 => n2, B2 => n1, A => n4, ZN => g_vector_0_0_port
                           );
   U2 : OAI21_X1 port map( B1 => A(0), B2 => B(0), A => Cin, ZN => n4);
   U3 : INV_X1 port map( A => A(0), ZN => n2);
   U4 : INV_X1 port map( A => B(0), ZN => n1);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity CARRY_GENERATOR_NBIT64_NBIT_PER_BLOCK4_1 is

   port( A, B : in std_logic_vector (63 downto 0);  Cin : in std_logic;  Co : 
         out std_logic_vector (15 downto 0));

end CARRY_GENERATOR_NBIT64_NBIT_PER_BLOCK4_1;

architecture SYN_structural of CARRY_GENERATOR_NBIT64_NBIT_PER_BLOCK4_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component G_BLOCK_1
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component G_BLOCK_2
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component G_BLOCK_3
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component G_BLOCK_4
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component G_BLOCK_5
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component G_BLOCK_6
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component G_BLOCK_7
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component G_BLOCK_8
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component G_BLOCK_9
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component G_BLOCK_10
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component G_BLOCK_11
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component G_BLOCK_12
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component PG_BLOCK_1
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_2
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_3
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_4
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component G_BLOCK_13
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component G_BLOCK_14
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component PG_BLOCK_5
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_6
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_7
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_8
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_9
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_10
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component G_BLOCK_15
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component PG_BLOCK_11
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_12
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_13
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_14
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_15
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_16
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_17
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component G_BLOCK_16
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component PG_BLOCK_18
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_19
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_20
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_21
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_22
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_23
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_24
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_25
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_26
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_27
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_28
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_29
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_30
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_31
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_32
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component G_BLOCK_17
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component PG_BLOCK_33
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_34
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_35
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_36
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_37
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_38
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_39
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_40
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_41
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_42
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_43
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_44
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_45
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_46
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_47
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_48
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_49
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_50
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_51
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_52
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_53
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_54
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_55
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_56
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_57
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_58
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_59
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_60
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_61
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_62
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_63
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component pg_net_1
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_2
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_3
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_4
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_5
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_6
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_7
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_8
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_9
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_10
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_11
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_12
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_13
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_14
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_15
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_16
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_17
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_18
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_19
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_20
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_21
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_22
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_23
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_24
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_25
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_26
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_27
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_28
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_29
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_30
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_31
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_32
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_33
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_34
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_35
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_36
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_37
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_38
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_39
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_40
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_41
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_42
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_43
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_44
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_45
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_46
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_47
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_48
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_49
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_50
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_51
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_52
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_53
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_54
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_55
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_56
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_57
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_58
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_59
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_60
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_61
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_62
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_63
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   signal Co_15_port, Co_14_port, Co_13_port, Co_12_port, Co_11_port, 
      Co_10_port, Co_9_port, Co_8_port, Co_7_port, Co_6_port, Co_5_port, 
      Co_4_port, Co_3_port, Co_2_port, Co_1_port, Co_0_port, g_vector_5_63_port
      , g_vector_5_59_port, g_vector_5_55_port, g_vector_5_51_port, 
      g_vector_4_63_port, g_vector_4_59_port, g_vector_4_47_port, 
      g_vector_4_43_port, g_vector_4_31_port, g_vector_4_27_port, 
      g_vector_3_63_port, g_vector_3_55_port, g_vector_3_47_port, 
      g_vector_3_39_port, g_vector_3_31_port, g_vector_3_23_port, 
      g_vector_3_15_port, g_vector_2_63_port, g_vector_2_59_port, 
      g_vector_2_55_port, g_vector_2_51_port, g_vector_2_47_port, 
      g_vector_2_43_port, g_vector_2_39_port, g_vector_2_35_port, 
      g_vector_2_31_port, g_vector_2_27_port, g_vector_2_23_port, 
      g_vector_2_19_port, g_vector_2_15_port, g_vector_2_11_port, 
      g_vector_2_7_port, g_vector_1_63_port, g_vector_1_61_port, 
      g_vector_1_59_port, g_vector_1_57_port, g_vector_1_55_port, 
      g_vector_1_53_port, g_vector_1_51_port, g_vector_1_49_port, 
      g_vector_1_47_port, g_vector_1_45_port, g_vector_1_43_port, 
      g_vector_1_41_port, g_vector_1_39_port, g_vector_1_37_port, 
      g_vector_1_35_port, g_vector_1_33_port, g_vector_1_31_port, 
      g_vector_1_29_port, g_vector_1_27_port, g_vector_1_25_port, 
      g_vector_1_23_port, g_vector_1_21_port, g_vector_1_19_port, 
      g_vector_1_17_port, g_vector_1_15_port, g_vector_1_13_port, 
      g_vector_1_11_port, g_vector_1_9_port, g_vector_1_7_port, 
      g_vector_1_5_port, g_vector_1_3_port, g_vector_1_1_port, 
      g_vector_0_63_port, g_vector_0_62_port, g_vector_0_61_port, 
      g_vector_0_60_port, g_vector_0_59_port, g_vector_0_58_port, 
      g_vector_0_57_port, g_vector_0_56_port, g_vector_0_55_port, 
      g_vector_0_54_port, g_vector_0_53_port, g_vector_0_52_port, 
      g_vector_0_51_port, g_vector_0_50_port, g_vector_0_49_port, 
      g_vector_0_48_port, g_vector_0_47_port, g_vector_0_46_port, 
      g_vector_0_45_port, g_vector_0_44_port, g_vector_0_43_port, 
      g_vector_0_42_port, g_vector_0_41_port, g_vector_0_40_port, 
      g_vector_0_39_port, g_vector_0_38_port, g_vector_0_37_port, 
      g_vector_0_36_port, g_vector_0_35_port, g_vector_0_34_port, 
      g_vector_0_33_port, g_vector_0_32_port, g_vector_0_31_port, 
      g_vector_0_30_port, g_vector_0_29_port, g_vector_0_28_port, 
      g_vector_0_27_port, g_vector_0_26_port, g_vector_0_25_port, 
      g_vector_0_24_port, g_vector_0_23_port, g_vector_0_22_port, 
      g_vector_0_21_port, g_vector_0_20_port, g_vector_0_19_port, 
      g_vector_0_18_port, g_vector_0_17_port, g_vector_0_16_port, 
      g_vector_0_15_port, g_vector_0_14_port, g_vector_0_13_port, 
      g_vector_0_12_port, g_vector_0_11_port, g_vector_0_10_port, 
      g_vector_0_9_port, g_vector_0_8_port, g_vector_0_7_port, 
      g_vector_0_6_port, g_vector_0_5_port, g_vector_0_4_port, 
      g_vector_0_3_port, g_vector_0_2_port, g_vector_0_1_port, 
      g_vector_0_0_port, p_vector_5_63_port, p_vector_5_59_port, 
      p_vector_5_55_port, p_vector_5_51_port, p_vector_4_63_port, 
      p_vector_4_59_port, p_vector_4_47_port, p_vector_4_43_port, 
      p_vector_4_31_port, p_vector_4_27_port, p_vector_3_63_port, 
      p_vector_3_55_port, p_vector_3_47_port, p_vector_3_39_port, 
      p_vector_3_31_port, p_vector_3_23_port, p_vector_3_15_port, 
      p_vector_2_63_port, p_vector_2_59_port, p_vector_2_55_port, 
      p_vector_2_51_port, p_vector_2_47_port, p_vector_2_43_port, 
      p_vector_2_39_port, p_vector_2_35_port, p_vector_2_31_port, 
      p_vector_2_27_port, p_vector_2_23_port, p_vector_2_19_port, 
      p_vector_2_15_port, p_vector_2_11_port, p_vector_2_7_port, 
      p_vector_1_63_port, p_vector_1_61_port, p_vector_1_59_port, 
      p_vector_1_57_port, p_vector_1_55_port, p_vector_1_53_port, 
      p_vector_1_51_port, p_vector_1_49_port, p_vector_1_47_port, 
      p_vector_1_45_port, p_vector_1_43_port, p_vector_1_41_port, 
      p_vector_1_39_port, p_vector_1_37_port, p_vector_1_35_port, 
      p_vector_1_33_port, p_vector_1_31_port, p_vector_1_29_port, 
      p_vector_1_27_port, p_vector_1_25_port, p_vector_1_23_port, 
      p_vector_1_21_port, p_vector_1_19_port, p_vector_1_17_port, 
      p_vector_1_15_port, p_vector_1_13_port, p_vector_1_11_port, 
      p_vector_1_9_port, p_vector_1_7_port, p_vector_1_5_port, 
      p_vector_1_3_port, p_vector_0_63_port, p_vector_0_62_port, 
      p_vector_0_61_port, p_vector_0_60_port, p_vector_0_59_port, 
      p_vector_0_58_port, p_vector_0_57_port, p_vector_0_56_port, 
      p_vector_0_55_port, p_vector_0_54_port, p_vector_0_53_port, 
      p_vector_0_52_port, p_vector_0_51_port, p_vector_0_50_port, 
      p_vector_0_49_port, p_vector_0_48_port, p_vector_0_47_port, 
      p_vector_0_46_port, p_vector_0_45_port, p_vector_0_44_port, 
      p_vector_0_43_port, p_vector_0_42_port, p_vector_0_41_port, 
      p_vector_0_40_port, p_vector_0_39_port, p_vector_0_38_port, 
      p_vector_0_37_port, p_vector_0_36_port, p_vector_0_35_port, 
      p_vector_0_34_port, p_vector_0_33_port, p_vector_0_32_port, 
      p_vector_0_31_port, p_vector_0_30_port, p_vector_0_29_port, 
      p_vector_0_28_port, p_vector_0_27_port, p_vector_0_26_port, 
      p_vector_0_25_port, p_vector_0_24_port, p_vector_0_23_port, 
      p_vector_0_22_port, p_vector_0_21_port, p_vector_0_20_port, 
      p_vector_0_19_port, p_vector_0_18_port, p_vector_0_17_port, 
      p_vector_0_16_port, p_vector_0_15_port, p_vector_0_14_port, 
      p_vector_0_13_port, p_vector_0_12_port, p_vector_0_11_port, 
      p_vector_0_10_port, p_vector_0_9_port, p_vector_0_8_port, 
      p_vector_0_7_port, p_vector_0_6_port, p_vector_0_5_port, 
      p_vector_0_4_port, p_vector_0_3_port, p_vector_0_2_port, 
      p_vector_0_1_port, n1, n2, n4 : std_logic;

begin
   Co <= ( Co_15_port, Co_14_port, Co_13_port, Co_12_port, Co_11_port, 
      Co_10_port, Co_9_port, Co_8_port, Co_7_port, Co_6_port, Co_5_port, 
      Co_4_port, Co_3_port, Co_2_port, Co_1_port, Co_0_port );
   
   pg_network_63 : pg_net_63 port map( a => A(63), b => B(63), p => 
                           p_vector_0_63_port, g => g_vector_0_63_port);
   pg_network_62 : pg_net_62 port map( a => A(62), b => B(62), p => 
                           p_vector_0_62_port, g => g_vector_0_62_port);
   pg_network_61 : pg_net_61 port map( a => A(61), b => B(61), p => 
                           p_vector_0_61_port, g => g_vector_0_61_port);
   pg_network_60 : pg_net_60 port map( a => A(60), b => B(60), p => 
                           p_vector_0_60_port, g => g_vector_0_60_port);
   pg_network_59 : pg_net_59 port map( a => A(59), b => B(59), p => 
                           p_vector_0_59_port, g => g_vector_0_59_port);
   pg_network_58 : pg_net_58 port map( a => A(58), b => B(58), p => 
                           p_vector_0_58_port, g => g_vector_0_58_port);
   pg_network_57 : pg_net_57 port map( a => A(57), b => B(57), p => 
                           p_vector_0_57_port, g => g_vector_0_57_port);
   pg_network_56 : pg_net_56 port map( a => A(56), b => B(56), p => 
                           p_vector_0_56_port, g => g_vector_0_56_port);
   pg_network_55 : pg_net_55 port map( a => A(55), b => B(55), p => 
                           p_vector_0_55_port, g => g_vector_0_55_port);
   pg_network_54 : pg_net_54 port map( a => A(54), b => B(54), p => 
                           p_vector_0_54_port, g => g_vector_0_54_port);
   pg_network_53 : pg_net_53 port map( a => A(53), b => B(53), p => 
                           p_vector_0_53_port, g => g_vector_0_53_port);
   pg_network_52 : pg_net_52 port map( a => A(52), b => B(52), p => 
                           p_vector_0_52_port, g => g_vector_0_52_port);
   pg_network_51 : pg_net_51 port map( a => A(51), b => B(51), p => 
                           p_vector_0_51_port, g => g_vector_0_51_port);
   pg_network_50 : pg_net_50 port map( a => A(50), b => B(50), p => 
                           p_vector_0_50_port, g => g_vector_0_50_port);
   pg_network_49 : pg_net_49 port map( a => A(49), b => B(49), p => 
                           p_vector_0_49_port, g => g_vector_0_49_port);
   pg_network_48 : pg_net_48 port map( a => A(48), b => B(48), p => 
                           p_vector_0_48_port, g => g_vector_0_48_port);
   pg_network_47 : pg_net_47 port map( a => A(47), b => B(47), p => 
                           p_vector_0_47_port, g => g_vector_0_47_port);
   pg_network_46 : pg_net_46 port map( a => A(46), b => B(46), p => 
                           p_vector_0_46_port, g => g_vector_0_46_port);
   pg_network_45 : pg_net_45 port map( a => A(45), b => B(45), p => 
                           p_vector_0_45_port, g => g_vector_0_45_port);
   pg_network_44 : pg_net_44 port map( a => A(44), b => B(44), p => 
                           p_vector_0_44_port, g => g_vector_0_44_port);
   pg_network_43 : pg_net_43 port map( a => A(43), b => B(43), p => 
                           p_vector_0_43_port, g => g_vector_0_43_port);
   pg_network_42 : pg_net_42 port map( a => A(42), b => B(42), p => 
                           p_vector_0_42_port, g => g_vector_0_42_port);
   pg_network_41 : pg_net_41 port map( a => A(41), b => B(41), p => 
                           p_vector_0_41_port, g => g_vector_0_41_port);
   pg_network_40 : pg_net_40 port map( a => A(40), b => B(40), p => 
                           p_vector_0_40_port, g => g_vector_0_40_port);
   pg_network_39 : pg_net_39 port map( a => A(39), b => B(39), p => 
                           p_vector_0_39_port, g => g_vector_0_39_port);
   pg_network_38 : pg_net_38 port map( a => A(38), b => B(38), p => 
                           p_vector_0_38_port, g => g_vector_0_38_port);
   pg_network_37 : pg_net_37 port map( a => A(37), b => B(37), p => 
                           p_vector_0_37_port, g => g_vector_0_37_port);
   pg_network_36 : pg_net_36 port map( a => A(36), b => B(36), p => 
                           p_vector_0_36_port, g => g_vector_0_36_port);
   pg_network_35 : pg_net_35 port map( a => A(35), b => B(35), p => 
                           p_vector_0_35_port, g => g_vector_0_35_port);
   pg_network_34 : pg_net_34 port map( a => A(34), b => B(34), p => 
                           p_vector_0_34_port, g => g_vector_0_34_port);
   pg_network_33 : pg_net_33 port map( a => A(33), b => B(33), p => 
                           p_vector_0_33_port, g => g_vector_0_33_port);
   pg_network_32 : pg_net_32 port map( a => A(32), b => B(32), p => 
                           p_vector_0_32_port, g => g_vector_0_32_port);
   pg_network_31 : pg_net_31 port map( a => A(31), b => B(31), p => 
                           p_vector_0_31_port, g => g_vector_0_31_port);
   pg_network_30 : pg_net_30 port map( a => A(30), b => B(30), p => 
                           p_vector_0_30_port, g => g_vector_0_30_port);
   pg_network_29 : pg_net_29 port map( a => A(29), b => B(29), p => 
                           p_vector_0_29_port, g => g_vector_0_29_port);
   pg_network_28 : pg_net_28 port map( a => A(28), b => B(28), p => 
                           p_vector_0_28_port, g => g_vector_0_28_port);
   pg_network_27 : pg_net_27 port map( a => A(27), b => B(27), p => 
                           p_vector_0_27_port, g => g_vector_0_27_port);
   pg_network_26 : pg_net_26 port map( a => A(26), b => B(26), p => 
                           p_vector_0_26_port, g => g_vector_0_26_port);
   pg_network_25 : pg_net_25 port map( a => A(25), b => B(25), p => 
                           p_vector_0_25_port, g => g_vector_0_25_port);
   pg_network_24 : pg_net_24 port map( a => A(24), b => B(24), p => 
                           p_vector_0_24_port, g => g_vector_0_24_port);
   pg_network_23 : pg_net_23 port map( a => A(23), b => B(23), p => 
                           p_vector_0_23_port, g => g_vector_0_23_port);
   pg_network_22 : pg_net_22 port map( a => A(22), b => B(22), p => 
                           p_vector_0_22_port, g => g_vector_0_22_port);
   pg_network_21 : pg_net_21 port map( a => A(21), b => B(21), p => 
                           p_vector_0_21_port, g => g_vector_0_21_port);
   pg_network_20 : pg_net_20 port map( a => A(20), b => B(20), p => 
                           p_vector_0_20_port, g => g_vector_0_20_port);
   pg_network_19 : pg_net_19 port map( a => A(19), b => B(19), p => 
                           p_vector_0_19_port, g => g_vector_0_19_port);
   pg_network_18 : pg_net_18 port map( a => A(18), b => B(18), p => 
                           p_vector_0_18_port, g => g_vector_0_18_port);
   pg_network_17 : pg_net_17 port map( a => A(17), b => B(17), p => 
                           p_vector_0_17_port, g => g_vector_0_17_port);
   pg_network_16 : pg_net_16 port map( a => A(16), b => B(16), p => 
                           p_vector_0_16_port, g => g_vector_0_16_port);
   pg_network_15 : pg_net_15 port map( a => A(15), b => B(15), p => 
                           p_vector_0_15_port, g => g_vector_0_15_port);
   pg_network_14 : pg_net_14 port map( a => A(14), b => B(14), p => 
                           p_vector_0_14_port, g => g_vector_0_14_port);
   pg_network_13 : pg_net_13 port map( a => A(13), b => B(13), p => 
                           p_vector_0_13_port, g => g_vector_0_13_port);
   pg_network_12 : pg_net_12 port map( a => A(12), b => B(12), p => 
                           p_vector_0_12_port, g => g_vector_0_12_port);
   pg_network_11 : pg_net_11 port map( a => A(11), b => B(11), p => 
                           p_vector_0_11_port, g => g_vector_0_11_port);
   pg_network_10 : pg_net_10 port map( a => A(10), b => B(10), p => 
                           p_vector_0_10_port, g => g_vector_0_10_port);
   pg_network_9 : pg_net_9 port map( a => A(9), b => B(9), p => 
                           p_vector_0_9_port, g => g_vector_0_9_port);
   pg_network_8 : pg_net_8 port map( a => A(8), b => B(8), p => 
                           p_vector_0_8_port, g => g_vector_0_8_port);
   pg_network_7 : pg_net_7 port map( a => A(7), b => B(7), p => 
                           p_vector_0_7_port, g => g_vector_0_7_port);
   pg_network_6 : pg_net_6 port map( a => A(6), b => B(6), p => 
                           p_vector_0_6_port, g => g_vector_0_6_port);
   pg_network_5 : pg_net_5 port map( a => A(5), b => B(5), p => 
                           p_vector_0_5_port, g => g_vector_0_5_port);
   pg_network_4 : pg_net_4 port map( a => A(4), b => B(4), p => 
                           p_vector_0_4_port, g => g_vector_0_4_port);
   pg_network_3 : pg_net_3 port map( a => A(3), b => B(3), p => 
                           p_vector_0_3_port, g => g_vector_0_3_port);
   pg_network_2 : pg_net_2 port map( a => A(2), b => B(2), p => 
                           p_vector_0_2_port, g => g_vector_0_2_port);
   pg_network_1 : pg_net_1 port map( a => A(1), b => B(1), p => 
                           p_vector_0_1_port, g => g_vector_0_1_port);
   std_PG_1_63 : PG_BLOCK_63 port map( p2 => p_vector_0_63_port, g2 => 
                           g_vector_0_63_port, p1 => p_vector_0_62_port, g1 => 
                           g_vector_0_62_port, PG_P => p_vector_1_63_port, PG_G
                           => g_vector_1_63_port);
   std_PG_1_61 : PG_BLOCK_62 port map( p2 => p_vector_0_61_port, g2 => 
                           g_vector_0_61_port, p1 => p_vector_0_60_port, g1 => 
                           g_vector_0_60_port, PG_P => p_vector_1_61_port, PG_G
                           => g_vector_1_61_port);
   std_PG_1_59 : PG_BLOCK_61 port map( p2 => p_vector_0_59_port, g2 => 
                           g_vector_0_59_port, p1 => p_vector_0_58_port, g1 => 
                           g_vector_0_58_port, PG_P => p_vector_1_59_port, PG_G
                           => g_vector_1_59_port);
   std_PG_1_57 : PG_BLOCK_60 port map( p2 => p_vector_0_57_port, g2 => 
                           g_vector_0_57_port, p1 => p_vector_0_56_port, g1 => 
                           g_vector_0_56_port, PG_P => p_vector_1_57_port, PG_G
                           => g_vector_1_57_port);
   std_PG_1_55 : PG_BLOCK_59 port map( p2 => p_vector_0_55_port, g2 => 
                           g_vector_0_55_port, p1 => p_vector_0_54_port, g1 => 
                           g_vector_0_54_port, PG_P => p_vector_1_55_port, PG_G
                           => g_vector_1_55_port);
   std_PG_1_53 : PG_BLOCK_58 port map( p2 => p_vector_0_53_port, g2 => 
                           g_vector_0_53_port, p1 => p_vector_0_52_port, g1 => 
                           g_vector_0_52_port, PG_P => p_vector_1_53_port, PG_G
                           => g_vector_1_53_port);
   std_PG_1_51 : PG_BLOCK_57 port map( p2 => p_vector_0_51_port, g2 => 
                           g_vector_0_51_port, p1 => p_vector_0_50_port, g1 => 
                           g_vector_0_50_port, PG_P => p_vector_1_51_port, PG_G
                           => g_vector_1_51_port);
   std_PG_1_49 : PG_BLOCK_56 port map( p2 => p_vector_0_49_port, g2 => 
                           g_vector_0_49_port, p1 => p_vector_0_48_port, g1 => 
                           g_vector_0_48_port, PG_P => p_vector_1_49_port, PG_G
                           => g_vector_1_49_port);
   std_PG_1_47 : PG_BLOCK_55 port map( p2 => p_vector_0_47_port, g2 => 
                           g_vector_0_47_port, p1 => p_vector_0_46_port, g1 => 
                           g_vector_0_46_port, PG_P => p_vector_1_47_port, PG_G
                           => g_vector_1_47_port);
   std_PG_1_45 : PG_BLOCK_54 port map( p2 => p_vector_0_45_port, g2 => 
                           g_vector_0_45_port, p1 => p_vector_0_44_port, g1 => 
                           g_vector_0_44_port, PG_P => p_vector_1_45_port, PG_G
                           => g_vector_1_45_port);
   std_PG_1_43 : PG_BLOCK_53 port map( p2 => p_vector_0_43_port, g2 => 
                           g_vector_0_43_port, p1 => p_vector_0_42_port, g1 => 
                           g_vector_0_42_port, PG_P => p_vector_1_43_port, PG_G
                           => g_vector_1_43_port);
   std_PG_1_41 : PG_BLOCK_52 port map( p2 => p_vector_0_41_port, g2 => 
                           g_vector_0_41_port, p1 => p_vector_0_40_port, g1 => 
                           g_vector_0_40_port, PG_P => p_vector_1_41_port, PG_G
                           => g_vector_1_41_port);
   std_PG_1_39 : PG_BLOCK_51 port map( p2 => p_vector_0_39_port, g2 => 
                           g_vector_0_39_port, p1 => p_vector_0_38_port, g1 => 
                           g_vector_0_38_port, PG_P => p_vector_1_39_port, PG_G
                           => g_vector_1_39_port);
   std_PG_1_37 : PG_BLOCK_50 port map( p2 => p_vector_0_37_port, g2 => 
                           g_vector_0_37_port, p1 => p_vector_0_36_port, g1 => 
                           g_vector_0_36_port, PG_P => p_vector_1_37_port, PG_G
                           => g_vector_1_37_port);
   std_PG_1_35 : PG_BLOCK_49 port map( p2 => p_vector_0_35_port, g2 => 
                           g_vector_0_35_port, p1 => p_vector_0_34_port, g1 => 
                           g_vector_0_34_port, PG_P => p_vector_1_35_port, PG_G
                           => g_vector_1_35_port);
   std_PG_1_33 : PG_BLOCK_48 port map( p2 => p_vector_0_33_port, g2 => 
                           g_vector_0_33_port, p1 => p_vector_0_32_port, g1 => 
                           g_vector_0_32_port, PG_P => p_vector_1_33_port, PG_G
                           => g_vector_1_33_port);
   std_PG_1_31 : PG_BLOCK_47 port map( p2 => p_vector_0_31_port, g2 => 
                           g_vector_0_31_port, p1 => p_vector_0_30_port, g1 => 
                           g_vector_0_30_port, PG_P => p_vector_1_31_port, PG_G
                           => g_vector_1_31_port);
   std_PG_1_29 : PG_BLOCK_46 port map( p2 => p_vector_0_29_port, g2 => 
                           g_vector_0_29_port, p1 => p_vector_0_28_port, g1 => 
                           g_vector_0_28_port, PG_P => p_vector_1_29_port, PG_G
                           => g_vector_1_29_port);
   std_PG_1_27 : PG_BLOCK_45 port map( p2 => p_vector_0_27_port, g2 => 
                           g_vector_0_27_port, p1 => p_vector_0_26_port, g1 => 
                           g_vector_0_26_port, PG_P => p_vector_1_27_port, PG_G
                           => g_vector_1_27_port);
   std_PG_1_25 : PG_BLOCK_44 port map( p2 => p_vector_0_25_port, g2 => 
                           g_vector_0_25_port, p1 => p_vector_0_24_port, g1 => 
                           g_vector_0_24_port, PG_P => p_vector_1_25_port, PG_G
                           => g_vector_1_25_port);
   std_PG_1_23 : PG_BLOCK_43 port map( p2 => p_vector_0_23_port, g2 => 
                           g_vector_0_23_port, p1 => p_vector_0_22_port, g1 => 
                           g_vector_0_22_port, PG_P => p_vector_1_23_port, PG_G
                           => g_vector_1_23_port);
   std_PG_1_21 : PG_BLOCK_42 port map( p2 => p_vector_0_21_port, g2 => 
                           g_vector_0_21_port, p1 => p_vector_0_20_port, g1 => 
                           g_vector_0_20_port, PG_P => p_vector_1_21_port, PG_G
                           => g_vector_1_21_port);
   std_PG_1_19 : PG_BLOCK_41 port map( p2 => p_vector_0_19_port, g2 => 
                           g_vector_0_19_port, p1 => p_vector_0_18_port, g1 => 
                           g_vector_0_18_port, PG_P => p_vector_1_19_port, PG_G
                           => g_vector_1_19_port);
   std_PG_1_17 : PG_BLOCK_40 port map( p2 => p_vector_0_17_port, g2 => 
                           g_vector_0_17_port, p1 => p_vector_0_16_port, g1 => 
                           g_vector_0_16_port, PG_P => p_vector_1_17_port, PG_G
                           => g_vector_1_17_port);
   std_PG_1_15 : PG_BLOCK_39 port map( p2 => p_vector_0_15_port, g2 => 
                           g_vector_0_15_port, p1 => p_vector_0_14_port, g1 => 
                           g_vector_0_14_port, PG_P => p_vector_1_15_port, PG_G
                           => g_vector_1_15_port);
   std_PG_1_13 : PG_BLOCK_38 port map( p2 => p_vector_0_13_port, g2 => 
                           g_vector_0_13_port, p1 => p_vector_0_12_port, g1 => 
                           g_vector_0_12_port, PG_P => p_vector_1_13_port, PG_G
                           => g_vector_1_13_port);
   std_PG_1_11 : PG_BLOCK_37 port map( p2 => p_vector_0_11_port, g2 => 
                           g_vector_0_11_port, p1 => p_vector_0_10_port, g1 => 
                           g_vector_0_10_port, PG_P => p_vector_1_11_port, PG_G
                           => g_vector_1_11_port);
   std_PG_1_9 : PG_BLOCK_36 port map( p2 => p_vector_0_9_port, g2 => 
                           g_vector_0_9_port, p1 => p_vector_0_8_port, g1 => 
                           g_vector_0_8_port, PG_P => p_vector_1_9_port, PG_G 
                           => g_vector_1_9_port);
   std_PG_1_7 : PG_BLOCK_35 port map( p2 => p_vector_0_7_port, g2 => 
                           g_vector_0_7_port, p1 => p_vector_0_6_port, g1 => 
                           g_vector_0_6_port, PG_P => p_vector_1_7_port, PG_G 
                           => g_vector_1_7_port);
   std_PG_1_5 : PG_BLOCK_34 port map( p2 => p_vector_0_5_port, g2 => 
                           g_vector_0_5_port, p1 => p_vector_0_4_port, g1 => 
                           g_vector_0_4_port, PG_P => p_vector_1_5_port, PG_G 
                           => g_vector_1_5_port);
   std_PG_1_3 : PG_BLOCK_33 port map( p2 => p_vector_0_3_port, g2 => 
                           g_vector_0_3_port, p1 => p_vector_0_2_port, g1 => 
                           g_vector_0_2_port, PG_P => p_vector_1_3_port, PG_G 
                           => g_vector_1_3_port);
   std_G_1_1 : G_BLOCK_17 port map( p2 => p_vector_0_1_port, g2 => 
                           g_vector_0_1_port, g1 => g_vector_0_0_port, G => 
                           g_vector_1_1_port);
   std_PG_2_63 : PG_BLOCK_32 port map( p2 => p_vector_1_63_port, g2 => 
                           g_vector_1_63_port, p1 => p_vector_1_61_port, g1 => 
                           g_vector_1_61_port, PG_P => p_vector_2_63_port, PG_G
                           => g_vector_2_63_port);
   std_PG_2_59 : PG_BLOCK_31 port map( p2 => p_vector_1_59_port, g2 => 
                           g_vector_1_59_port, p1 => p_vector_1_57_port, g1 => 
                           g_vector_1_57_port, PG_P => p_vector_2_59_port, PG_G
                           => g_vector_2_59_port);
   std_PG_2_55 : PG_BLOCK_30 port map( p2 => p_vector_1_55_port, g2 => 
                           g_vector_1_55_port, p1 => p_vector_1_53_port, g1 => 
                           g_vector_1_53_port, PG_P => p_vector_2_55_port, PG_G
                           => g_vector_2_55_port);
   std_PG_2_51 : PG_BLOCK_29 port map( p2 => p_vector_1_51_port, g2 => 
                           g_vector_1_51_port, p1 => p_vector_1_49_port, g1 => 
                           g_vector_1_49_port, PG_P => p_vector_2_51_port, PG_G
                           => g_vector_2_51_port);
   std_PG_2_47 : PG_BLOCK_28 port map( p2 => p_vector_1_47_port, g2 => 
                           g_vector_1_47_port, p1 => p_vector_1_45_port, g1 => 
                           g_vector_1_45_port, PG_P => p_vector_2_47_port, PG_G
                           => g_vector_2_47_port);
   std_PG_2_43 : PG_BLOCK_27 port map( p2 => p_vector_1_43_port, g2 => 
                           g_vector_1_43_port, p1 => p_vector_1_41_port, g1 => 
                           g_vector_1_41_port, PG_P => p_vector_2_43_port, PG_G
                           => g_vector_2_43_port);
   std_PG_2_39 : PG_BLOCK_26 port map( p2 => p_vector_1_39_port, g2 => 
                           g_vector_1_39_port, p1 => p_vector_1_37_port, g1 => 
                           g_vector_1_37_port, PG_P => p_vector_2_39_port, PG_G
                           => g_vector_2_39_port);
   std_PG_2_35 : PG_BLOCK_25 port map( p2 => p_vector_1_35_port, g2 => 
                           g_vector_1_35_port, p1 => p_vector_1_33_port, g1 => 
                           g_vector_1_33_port, PG_P => p_vector_2_35_port, PG_G
                           => g_vector_2_35_port);
   std_PG_2_31 : PG_BLOCK_24 port map( p2 => p_vector_1_31_port, g2 => 
                           g_vector_1_31_port, p1 => p_vector_1_29_port, g1 => 
                           g_vector_1_29_port, PG_P => p_vector_2_31_port, PG_G
                           => g_vector_2_31_port);
   std_PG_2_27 : PG_BLOCK_23 port map( p2 => p_vector_1_27_port, g2 => 
                           g_vector_1_27_port, p1 => p_vector_1_25_port, g1 => 
                           g_vector_1_25_port, PG_P => p_vector_2_27_port, PG_G
                           => g_vector_2_27_port);
   std_PG_2_23 : PG_BLOCK_22 port map( p2 => p_vector_1_23_port, g2 => 
                           g_vector_1_23_port, p1 => p_vector_1_21_port, g1 => 
                           g_vector_1_21_port, PG_P => p_vector_2_23_port, PG_G
                           => g_vector_2_23_port);
   std_PG_2_19 : PG_BLOCK_21 port map( p2 => p_vector_1_19_port, g2 => 
                           g_vector_1_19_port, p1 => p_vector_1_17_port, g1 => 
                           g_vector_1_17_port, PG_P => p_vector_2_19_port, PG_G
                           => g_vector_2_19_port);
   std_PG_2_15 : PG_BLOCK_20 port map( p2 => p_vector_1_15_port, g2 => 
                           g_vector_1_15_port, p1 => p_vector_1_13_port, g1 => 
                           g_vector_1_13_port, PG_P => p_vector_2_15_port, PG_G
                           => g_vector_2_15_port);
   std_PG_2_11 : PG_BLOCK_19 port map( p2 => p_vector_1_11_port, g2 => 
                           g_vector_1_11_port, p1 => p_vector_1_9_port, g1 => 
                           g_vector_1_9_port, PG_P => p_vector_2_11_port, PG_G 
                           => g_vector_2_11_port);
   std_PG_2_7 : PG_BLOCK_18 port map( p2 => p_vector_1_7_port, g2 => 
                           g_vector_1_7_port, p1 => p_vector_1_5_port, g1 => 
                           g_vector_1_5_port, PG_P => p_vector_2_7_port, PG_G 
                           => g_vector_2_7_port);
   std_G_2_3 : G_BLOCK_16 port map( p2 => p_vector_1_3_port, g2 => 
                           g_vector_1_3_port, g1 => g_vector_1_1_port, G => 
                           Co_0_port);
   std_PG_3_63 : PG_BLOCK_17 port map( p2 => p_vector_2_63_port, g2 => 
                           g_vector_2_63_port, p1 => p_vector_2_59_port, g1 => 
                           g_vector_2_59_port, PG_P => p_vector_3_63_port, PG_G
                           => g_vector_3_63_port);
   std_PG_3_55 : PG_BLOCK_16 port map( p2 => p_vector_2_55_port, g2 => 
                           g_vector_2_55_port, p1 => p_vector_2_51_port, g1 => 
                           g_vector_2_51_port, PG_P => p_vector_3_55_port, PG_G
                           => g_vector_3_55_port);
   std_PG_3_47 : PG_BLOCK_15 port map( p2 => p_vector_2_47_port, g2 => 
                           g_vector_2_47_port, p1 => p_vector_2_43_port, g1 => 
                           g_vector_2_43_port, PG_P => p_vector_3_47_port, PG_G
                           => g_vector_3_47_port);
   std_PG_3_39 : PG_BLOCK_14 port map( p2 => p_vector_2_39_port, g2 => 
                           g_vector_2_39_port, p1 => p_vector_2_35_port, g1 => 
                           g_vector_2_35_port, PG_P => p_vector_3_39_port, PG_G
                           => g_vector_3_39_port);
   std_PG_3_31 : PG_BLOCK_13 port map( p2 => p_vector_2_31_port, g2 => 
                           g_vector_2_31_port, p1 => p_vector_2_27_port, g1 => 
                           g_vector_2_27_port, PG_P => p_vector_3_31_port, PG_G
                           => g_vector_3_31_port);
   std_PG_3_23 : PG_BLOCK_12 port map( p2 => p_vector_2_23_port, g2 => 
                           g_vector_2_23_port, p1 => p_vector_2_19_port, g1 => 
                           g_vector_2_19_port, PG_P => p_vector_3_23_port, PG_G
                           => g_vector_3_23_port);
   std_PG_3_15 : PG_BLOCK_11 port map( p2 => p_vector_2_15_port, g2 => 
                           g_vector_2_15_port, p1 => p_vector_2_11_port, g1 => 
                           g_vector_2_11_port, PG_P => p_vector_3_15_port, PG_G
                           => g_vector_3_15_port);
   std_G_3_7 : G_BLOCK_15 port map( p2 => p_vector_2_7_port, g2 => 
                           g_vector_2_7_port, g1 => Co_0_port, G => Co_1_port);
   std_PG_4_63 : PG_BLOCK_10 port map( p2 => p_vector_3_63_port, g2 => 
                           g_vector_3_63_port, p1 => p_vector_3_55_port, g1 => 
                           g_vector_3_55_port, PG_P => p_vector_4_63_port, PG_G
                           => g_vector_4_63_port);
   add_PG_4_63_1 : PG_BLOCK_9 port map( p2 => p_vector_2_59_port, g2 => 
                           g_vector_2_59_port, p1 => p_vector_3_55_port, g1 => 
                           g_vector_3_55_port, PG_P => p_vector_4_59_port, PG_G
                           => g_vector_4_59_port);
   std_PG_4_47 : PG_BLOCK_8 port map( p2 => p_vector_3_47_port, g2 => 
                           g_vector_3_47_port, p1 => p_vector_3_39_port, g1 => 
                           g_vector_3_39_port, PG_P => p_vector_4_47_port, PG_G
                           => g_vector_4_47_port);
   add_PG_4_47_1 : PG_BLOCK_7 port map( p2 => p_vector_2_43_port, g2 => 
                           g_vector_2_43_port, p1 => p_vector_3_39_port, g1 => 
                           g_vector_3_39_port, PG_P => p_vector_4_43_port, PG_G
                           => g_vector_4_43_port);
   std_PG_4_31 : PG_BLOCK_6 port map( p2 => p_vector_3_31_port, g2 => 
                           g_vector_3_31_port, p1 => p_vector_3_23_port, g1 => 
                           g_vector_3_23_port, PG_P => p_vector_4_31_port, PG_G
                           => g_vector_4_31_port);
   add_PG_4_31_1 : PG_BLOCK_5 port map( p2 => p_vector_2_27_port, g2 => 
                           g_vector_2_27_port, p1 => p_vector_3_23_port, g1 => 
                           g_vector_3_23_port, PG_P => p_vector_4_27_port, PG_G
                           => g_vector_4_27_port);
   std_G_4_15 : G_BLOCK_14 port map( p2 => p_vector_3_15_port, g2 => 
                           g_vector_3_15_port, g1 => Co_1_port, G => Co_3_port)
                           ;
   add_G_4_15_1 : G_BLOCK_13 port map( p2 => p_vector_2_11_port, g2 => 
                           g_vector_2_11_port, g1 => Co_1_port, G => Co_2_port)
                           ;
   std_PG_5_63 : PG_BLOCK_4 port map( p2 => p_vector_4_63_port, g2 => 
                           g_vector_4_63_port, p1 => p_vector_4_47_port, g1 => 
                           g_vector_4_47_port, PG_P => p_vector_5_63_port, PG_G
                           => g_vector_5_63_port);
   add_PG_5_63_1 : PG_BLOCK_3 port map( p2 => p_vector_4_59_port, g2 => 
                           g_vector_4_59_port, p1 => p_vector_4_47_port, g1 => 
                           g_vector_4_47_port, PG_P => p_vector_5_59_port, PG_G
                           => g_vector_5_59_port);
   add_PG_5_63_2 : PG_BLOCK_2 port map( p2 => p_vector_3_55_port, g2 => 
                           g_vector_3_55_port, p1 => p_vector_4_47_port, g1 => 
                           g_vector_4_47_port, PG_P => p_vector_5_55_port, PG_G
                           => g_vector_5_55_port);
   add_PG_5_63_3 : PG_BLOCK_1 port map( p2 => p_vector_2_51_port, g2 => 
                           g_vector_2_51_port, p1 => p_vector_4_47_port, g1 => 
                           g_vector_4_47_port, PG_P => p_vector_5_51_port, PG_G
                           => g_vector_5_51_port);
   std_G_5_31 : G_BLOCK_12 port map( p2 => p_vector_4_31_port, g2 => 
                           g_vector_4_31_port, g1 => Co_3_port, G => Co_7_port)
                           ;
   add_G_5_31_1 : G_BLOCK_11 port map( p2 => p_vector_4_27_port, g2 => 
                           g_vector_4_27_port, g1 => Co_3_port, G => Co_6_port)
                           ;
   add_G_5_31_2 : G_BLOCK_10 port map( p2 => p_vector_3_23_port, g2 => 
                           g_vector_3_23_port, g1 => Co_3_port, G => Co_5_port)
                           ;
   add_G_5_31_3 : G_BLOCK_9 port map( p2 => p_vector_2_19_port, g2 => 
                           g_vector_2_19_port, g1 => Co_3_port, G => Co_4_port)
                           ;
   std_G_6_63 : G_BLOCK_8 port map( p2 => p_vector_5_63_port, g2 => 
                           g_vector_5_63_port, g1 => Co_7_port, G => Co_15_port
                           );
   add_G_6_63_1 : G_BLOCK_7 port map( p2 => p_vector_5_59_port, g2 => 
                           g_vector_5_59_port, g1 => Co_7_port, G => Co_14_port
                           );
   add_G_6_63_2 : G_BLOCK_6 port map( p2 => p_vector_5_55_port, g2 => 
                           g_vector_5_55_port, g1 => Co_7_port, G => Co_13_port
                           );
   add_G_6_63_3 : G_BLOCK_5 port map( p2 => p_vector_5_51_port, g2 => 
                           g_vector_5_51_port, g1 => Co_7_port, G => Co_12_port
                           );
   add_G_6_63_4 : G_BLOCK_4 port map( p2 => p_vector_4_47_port, g2 => 
                           g_vector_4_47_port, g1 => Co_7_port, G => Co_11_port
                           );
   add_G_6_63_5 : G_BLOCK_3 port map( p2 => p_vector_4_43_port, g2 => 
                           g_vector_4_43_port, g1 => Co_7_port, G => Co_10_port
                           );
   add_G_6_63_6 : G_BLOCK_2 port map( p2 => p_vector_3_39_port, g2 => 
                           g_vector_3_39_port, g1 => Co_7_port, G => Co_9_port)
                           ;
   add_G_6_63_7 : G_BLOCK_1 port map( p2 => p_vector_2_35_port, g2 => 
                           g_vector_2_35_port, g1 => Co_7_port, G => Co_8_port)
                           ;
   U1 : OAI21_X1 port map( B1 => n2, B2 => n1, A => n4, ZN => g_vector_0_0_port
                           );
   U2 : OAI21_X1 port map( B1 => A(0), B2 => B(0), A => Cin, ZN => n4);
   U3 : INV_X1 port map( A => A(0), ZN => n2);
   U4 : INV_X1 port map( A => B(0), ZN => n1);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand41_31 is

   port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);

end nand41_31;

architecture SYN_behavioral of nand41_31 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => in4, A2 => in3, A3 => in2, A4 => in1, ZN => o)
                           ;

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand41_30 is

   port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);

end nand41_30;

architecture SYN_behavioral of nand41_30 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => in4, A2 => in3, A3 => in2, A4 => in1, ZN => o)
                           ;

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand41_29 is

   port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);

end nand41_29;

architecture SYN_behavioral of nand41_29 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => in4, A2 => in3, A3 => in2, A4 => in1, ZN => o)
                           ;

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand41_28 is

   port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);

end nand41_28;

architecture SYN_behavioral of nand41_28 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => in4, A2 => in3, A3 => in2, A4 => in1, ZN => o)
                           ;

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand41_27 is

   port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);

end nand41_27;

architecture SYN_behavioral of nand41_27 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => in4, A2 => in3, A3 => in2, A4 => in1, ZN => o)
                           ;

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand41_26 is

   port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);

end nand41_26;

architecture SYN_behavioral of nand41_26 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => in4, A2 => in3, A3 => in2, A4 => in1, ZN => o)
                           ;

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand41_25 is

   port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);

end nand41_25;

architecture SYN_behavioral of nand41_25 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => in4, A2 => in3, A3 => in2, A4 => in1, ZN => o)
                           ;

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand41_24 is

   port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);

end nand41_24;

architecture SYN_behavioral of nand41_24 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => in4, A2 => in3, A3 => in2, A4 => in1, ZN => o)
                           ;

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand41_23 is

   port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);

end nand41_23;

architecture SYN_behavioral of nand41_23 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => in4, A2 => in3, A3 => in2, A4 => in1, ZN => o)
                           ;

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand41_22 is

   port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);

end nand41_22;

architecture SYN_behavioral of nand41_22 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => in4, A2 => in3, A3 => in2, A4 => in1, ZN => o)
                           ;

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand41_21 is

   port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);

end nand41_21;

architecture SYN_behavioral of nand41_21 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => in4, A2 => in3, A3 => in2, A4 => in1, ZN => o)
                           ;

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand41_20 is

   port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);

end nand41_20;

architecture SYN_behavioral of nand41_20 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => in4, A2 => in3, A3 => in2, A4 => in1, ZN => o)
                           ;

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand41_19 is

   port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);

end nand41_19;

architecture SYN_behavioral of nand41_19 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => in4, A2 => in3, A3 => in2, A4 => in1, ZN => o)
                           ;

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand41_18 is

   port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);

end nand41_18;

architecture SYN_behavioral of nand41_18 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => in4, A2 => in3, A3 => in2, A4 => in1, ZN => o)
                           ;

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand41_17 is

   port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);

end nand41_17;

architecture SYN_behavioral of nand41_17 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => in4, A2 => in3, A3 => in2, A4 => in1, ZN => o)
                           ;

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand41_16 is

   port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);

end nand41_16;

architecture SYN_behavioral of nand41_16 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => in4, A2 => in3, A3 => in2, A4 => in1, ZN => o)
                           ;

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand41_15 is

   port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);

end nand41_15;

architecture SYN_behavioral of nand41_15 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => in4, A2 => in3, A3 => in2, A4 => in1, ZN => o)
                           ;

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand41_14 is

   port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);

end nand41_14;

architecture SYN_behavioral of nand41_14 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => in4, A2 => in3, A3 => in2, A4 => in1, ZN => o)
                           ;

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand41_13 is

   port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);

end nand41_13;

architecture SYN_behavioral of nand41_13 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => in4, A2 => in3, A3 => in2, A4 => in1, ZN => o)
                           ;

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand41_12 is

   port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);

end nand41_12;

architecture SYN_behavioral of nand41_12 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => in4, A2 => in3, A3 => in2, A4 => in1, ZN => o)
                           ;

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand41_11 is

   port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);

end nand41_11;

architecture SYN_behavioral of nand41_11 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => in4, A2 => in3, A3 => in2, A4 => in1, ZN => o)
                           ;

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand41_10 is

   port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);

end nand41_10;

architecture SYN_behavioral of nand41_10 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => in4, A2 => in3, A3 => in2, A4 => in1, ZN => o)
                           ;

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand41_9 is

   port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);

end nand41_9;

architecture SYN_behavioral of nand41_9 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => in4, A2 => in3, A3 => in2, A4 => in1, ZN => o)
                           ;

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand41_8 is

   port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);

end nand41_8;

architecture SYN_behavioral of nand41_8 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => in4, A2 => in3, A3 => in2, A4 => in1, ZN => o)
                           ;

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand41_7 is

   port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);

end nand41_7;

architecture SYN_behavioral of nand41_7 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => in4, A2 => in3, A3 => in2, A4 => in1, ZN => o)
                           ;

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand41_6 is

   port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);

end nand41_6;

architecture SYN_behavioral of nand41_6 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => in4, A2 => in3, A3 => in2, A4 => in1, ZN => o)
                           ;

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand41_5 is

   port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);

end nand41_5;

architecture SYN_behavioral of nand41_5 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => in4, A2 => in3, A3 => in2, A4 => in1, ZN => o)
                           ;

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand41_4 is

   port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);

end nand41_4;

architecture SYN_behavioral of nand41_4 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => in4, A2 => in3, A3 => in2, A4 => in1, ZN => o)
                           ;

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand41_3 is

   port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);

end nand41_3;

architecture SYN_behavioral of nand41_3 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => in4, A2 => in3, A3 => in2, A4 => in1, ZN => o)
                           ;

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand41_2 is

   port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);

end nand41_2;

architecture SYN_behavioral of nand41_2 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => in4, A2 => in3, A3 => in2, A4 => in1, ZN => o)
                           ;

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand41_1 is

   port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);

end nand41_1;

architecture SYN_behavioral of nand41_1 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => in4, A2 => in3, A3 => in2, A4 => in1, ZN => o)
                           ;

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_127 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_127;

architecture SYN_behavioral of nand31_127 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_126 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_126;

architecture SYN_behavioral of nand31_126 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_125 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_125;

architecture SYN_behavioral of nand31_125 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_124 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_124;

architecture SYN_behavioral of nand31_124 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_123 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_123;

architecture SYN_behavioral of nand31_123 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_122 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_122;

architecture SYN_behavioral of nand31_122 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_121 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_121;

architecture SYN_behavioral of nand31_121 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_120 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_120;

architecture SYN_behavioral of nand31_120 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_119 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_119;

architecture SYN_behavioral of nand31_119 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_118 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_118;

architecture SYN_behavioral of nand31_118 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_117 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_117;

architecture SYN_behavioral of nand31_117 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_116 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_116;

architecture SYN_behavioral of nand31_116 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_115 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_115;

architecture SYN_behavioral of nand31_115 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_114 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_114;

architecture SYN_behavioral of nand31_114 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_113 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_113;

architecture SYN_behavioral of nand31_113 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_112 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_112;

architecture SYN_behavioral of nand31_112 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_111 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_111;

architecture SYN_behavioral of nand31_111 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_110 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_110;

architecture SYN_behavioral of nand31_110 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_109 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_109;

architecture SYN_behavioral of nand31_109 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_108 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_108;

architecture SYN_behavioral of nand31_108 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_107 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_107;

architecture SYN_behavioral of nand31_107 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_106 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_106;

architecture SYN_behavioral of nand31_106 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_105 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_105;

architecture SYN_behavioral of nand31_105 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_104 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_104;

architecture SYN_behavioral of nand31_104 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_103 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_103;

architecture SYN_behavioral of nand31_103 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_102 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_102;

architecture SYN_behavioral of nand31_102 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_101 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_101;

architecture SYN_behavioral of nand31_101 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_100 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_100;

architecture SYN_behavioral of nand31_100 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_99 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_99;

architecture SYN_behavioral of nand31_99 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_98 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_98;

architecture SYN_behavioral of nand31_98 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_97 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_97;

architecture SYN_behavioral of nand31_97 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_96 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_96;

architecture SYN_behavioral of nand31_96 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_95 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_95;

architecture SYN_behavioral of nand31_95 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_94 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_94;

architecture SYN_behavioral of nand31_94 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_93 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_93;

architecture SYN_behavioral of nand31_93 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_92 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_92;

architecture SYN_behavioral of nand31_92 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_91 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_91;

architecture SYN_behavioral of nand31_91 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_90 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_90;

architecture SYN_behavioral of nand31_90 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_89 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_89;

architecture SYN_behavioral of nand31_89 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_88 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_88;

architecture SYN_behavioral of nand31_88 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_87 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_87;

architecture SYN_behavioral of nand31_87 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_86 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_86;

architecture SYN_behavioral of nand31_86 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_85 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_85;

architecture SYN_behavioral of nand31_85 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_84 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_84;

architecture SYN_behavioral of nand31_84 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_83 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_83;

architecture SYN_behavioral of nand31_83 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_82 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_82;

architecture SYN_behavioral of nand31_82 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_81 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_81;

architecture SYN_behavioral of nand31_81 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_80 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_80;

architecture SYN_behavioral of nand31_80 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_79 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_79;

architecture SYN_behavioral of nand31_79 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_78 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_78;

architecture SYN_behavioral of nand31_78 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_77 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_77;

architecture SYN_behavioral of nand31_77 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_76 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_76;

architecture SYN_behavioral of nand31_76 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_75 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_75;

architecture SYN_behavioral of nand31_75 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_74 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_74;

architecture SYN_behavioral of nand31_74 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_73 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_73;

architecture SYN_behavioral of nand31_73 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_72 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_72;

architecture SYN_behavioral of nand31_72 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_71 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_71;

architecture SYN_behavioral of nand31_71 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_70 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_70;

architecture SYN_behavioral of nand31_70 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_69 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_69;

architecture SYN_behavioral of nand31_69 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_68 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_68;

architecture SYN_behavioral of nand31_68 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_67 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_67;

architecture SYN_behavioral of nand31_67 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_66 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_66;

architecture SYN_behavioral of nand31_66 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_65 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_65;

architecture SYN_behavioral of nand31_65 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_64 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_64;

architecture SYN_behavioral of nand31_64 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_63 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_63;

architecture SYN_behavioral of nand31_63 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_62 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_62;

architecture SYN_behavioral of nand31_62 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_61 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_61;

architecture SYN_behavioral of nand31_61 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_60 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_60;

architecture SYN_behavioral of nand31_60 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_59 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_59;

architecture SYN_behavioral of nand31_59 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_58 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_58;

architecture SYN_behavioral of nand31_58 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_57 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_57;

architecture SYN_behavioral of nand31_57 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_56 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_56;

architecture SYN_behavioral of nand31_56 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_55 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_55;

architecture SYN_behavioral of nand31_55 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_54 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_54;

architecture SYN_behavioral of nand31_54 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_53 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_53;

architecture SYN_behavioral of nand31_53 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_52 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_52;

architecture SYN_behavioral of nand31_52 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_51 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_51;

architecture SYN_behavioral of nand31_51 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_50 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_50;

architecture SYN_behavioral of nand31_50 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_49 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_49;

architecture SYN_behavioral of nand31_49 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_48 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_48;

architecture SYN_behavioral of nand31_48 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_47 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_47;

architecture SYN_behavioral of nand31_47 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_46 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_46;

architecture SYN_behavioral of nand31_46 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_45 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_45;

architecture SYN_behavioral of nand31_45 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_44 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_44;

architecture SYN_behavioral of nand31_44 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_43 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_43;

architecture SYN_behavioral of nand31_43 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_42 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_42;

architecture SYN_behavioral of nand31_42 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_41 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_41;

architecture SYN_behavioral of nand31_41 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_40 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_40;

architecture SYN_behavioral of nand31_40 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_39 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_39;

architecture SYN_behavioral of nand31_39 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_38 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_38;

architecture SYN_behavioral of nand31_38 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_37 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_37;

architecture SYN_behavioral of nand31_37 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_36 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_36;

architecture SYN_behavioral of nand31_36 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_35 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_35;

architecture SYN_behavioral of nand31_35 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_34 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_34;

architecture SYN_behavioral of nand31_34 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_33 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_33;

architecture SYN_behavioral of nand31_33 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_32 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_32;

architecture SYN_behavioral of nand31_32 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_31 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_31;

architecture SYN_behavioral of nand31_31 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_30 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_30;

architecture SYN_behavioral of nand31_30 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_29 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_29;

architecture SYN_behavioral of nand31_29 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_28 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_28;

architecture SYN_behavioral of nand31_28 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_27 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_27;

architecture SYN_behavioral of nand31_27 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_26 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_26;

architecture SYN_behavioral of nand31_26 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_25 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_25;

architecture SYN_behavioral of nand31_25 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_24 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_24;

architecture SYN_behavioral of nand31_24 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_23 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_23;

architecture SYN_behavioral of nand31_23 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_22 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_22;

architecture SYN_behavioral of nand31_22 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_21 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_21;

architecture SYN_behavioral of nand31_21 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_20 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_20;

architecture SYN_behavioral of nand31_20 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_19 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_19;

architecture SYN_behavioral of nand31_19 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_18 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_18;

architecture SYN_behavioral of nand31_18 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_17 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_17;

architecture SYN_behavioral of nand31_17 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_16 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_16;

architecture SYN_behavioral of nand31_16 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_15 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_15;

architecture SYN_behavioral of nand31_15 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_14 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_14;

architecture SYN_behavioral of nand31_14 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_13 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_13;

architecture SYN_behavioral of nand31_13 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_12 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_12;

architecture SYN_behavioral of nand31_12 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_11 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_11;

architecture SYN_behavioral of nand31_11 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_10 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_10;

architecture SYN_behavioral of nand31_10 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_9 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_9;

architecture SYN_behavioral of nand31_9 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_8 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_8;

architecture SYN_behavioral of nand31_8 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_7 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_7;

architecture SYN_behavioral of nand31_7 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_6 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_6;

architecture SYN_behavioral of nand31_6 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_5 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_5;

architecture SYN_behavioral of nand31_5 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_4 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_4;

architecture SYN_behavioral of nand31_4 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_3 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_3;

architecture SYN_behavioral of nand31_3 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_2 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_2;

architecture SYN_behavioral of nand31_2 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_1 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_1;

architecture SYN_behavioral of nand31_1 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_63 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_63;

architecture SYN_structural of MUX21_GENERIC_NBIT4_63 is

   component MUX21_385
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_386
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_387
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_388
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_388 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_387 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_386 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_385 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_62 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_62;

architecture SYN_structural of MUX21_GENERIC_NBIT4_62 is

   component MUX21_381
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_382
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_383
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_384
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_384 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_383 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_382 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_381 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_61 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_61;

architecture SYN_structural of MUX21_GENERIC_NBIT4_61 is

   component MUX21_377
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_378
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_379
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_380
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_380 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_379 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_378 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_377 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_60 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_60;

architecture SYN_structural of MUX21_GENERIC_NBIT4_60 is

   component MUX21_373
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_374
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_375
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_376
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_376 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_375 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_374 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_373 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_59 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_59;

architecture SYN_structural of MUX21_GENERIC_NBIT4_59 is

   component MUX21_369
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_370
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_371
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_372
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_372 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_371 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_370 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_369 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_58 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_58;

architecture SYN_structural of MUX21_GENERIC_NBIT4_58 is

   component MUX21_365
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_366
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_367
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_368
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_368 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_367 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_366 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_365 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_57 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_57;

architecture SYN_structural of MUX21_GENERIC_NBIT4_57 is

   component MUX21_361
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_362
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_363
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_364
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_364 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_363 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_362 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_361 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_56 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_56;

architecture SYN_structural of MUX21_GENERIC_NBIT4_56 is

   component MUX21_221
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_222
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_223
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_224
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_224 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_223 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_222 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_221 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_55 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_55;

architecture SYN_structural of MUX21_GENERIC_NBIT4_55 is

   component MUX21_217
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_218
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_219
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_220
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_220 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_219 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_218 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_217 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_54 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_54;

architecture SYN_structural of MUX21_GENERIC_NBIT4_54 is

   component MUX21_213
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_214
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_215
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_216
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_216 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_215 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_214 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_213 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_53 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_53;

architecture SYN_structural of MUX21_GENERIC_NBIT4_53 is

   component MUX21_209
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_210
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_211
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_212
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_212 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_211 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_210 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_209 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_52 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_52;

architecture SYN_structural of MUX21_GENERIC_NBIT4_52 is

   component MUX21_205
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_206
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_207
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_208
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_208 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_207 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_206 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_205 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_51 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_51;

architecture SYN_structural of MUX21_GENERIC_NBIT4_51 is

   component MUX21_201
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_202
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_203
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_204
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_204 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_203 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_202 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_201 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_50 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_50;

architecture SYN_structural of MUX21_GENERIC_NBIT4_50 is

   component MUX21_197
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_198
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_199
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_200
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_200 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_199 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_198 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_197 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_49 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_49;

architecture SYN_structural of MUX21_GENERIC_NBIT4_49 is

   component MUX21_193
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_194
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_195
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_196
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_196 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_195 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_194 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_193 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_48 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_48;

architecture SYN_structural of MUX21_GENERIC_NBIT4_48 is

   component MUX21_189
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_190
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_191
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_192
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_192 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_191 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_190 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_189 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_47 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_47;

architecture SYN_structural of MUX21_GENERIC_NBIT4_47 is

   component MUX21_185
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_186
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_187
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_188
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_188 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_187 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_186 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_185 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_46 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_46;

architecture SYN_structural of MUX21_GENERIC_NBIT4_46 is

   component MUX21_181
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_182
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_183
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_184
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_184 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_183 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_182 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_181 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_45 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_45;

architecture SYN_structural of MUX21_GENERIC_NBIT4_45 is

   component MUX21_177
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_178
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_179
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_180
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_180 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_179 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_178 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_177 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_44 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_44;

architecture SYN_structural of MUX21_GENERIC_NBIT4_44 is

   component MUX21_173
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_174
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_175
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_176
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_176 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_175 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_174 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_173 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_43 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_43;

architecture SYN_structural of MUX21_GENERIC_NBIT4_43 is

   component MUX21_169
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_170
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_171
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_172
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_172 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_171 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_170 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_169 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_42 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_42;

architecture SYN_structural of MUX21_GENERIC_NBIT4_42 is

   component MUX21_165
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_166
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_167
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_168
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_168 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_167 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_166 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_165 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_41 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_41;

architecture SYN_structural of MUX21_GENERIC_NBIT4_41 is

   component MUX21_161
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_162
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_163
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_164
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_164 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_163 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_162 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_161 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_40 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_40;

architecture SYN_structural of MUX21_GENERIC_NBIT4_40 is

   component MUX21_157
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_158
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_159
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_160
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_160 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_159 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_158 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_157 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_39 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_39;

architecture SYN_structural of MUX21_GENERIC_NBIT4_39 is

   component MUX21_153
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_154
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_155
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_156
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_156 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_155 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_154 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_153 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_38 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_38;

architecture SYN_structural of MUX21_GENERIC_NBIT4_38 is

   component MUX21_149
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_150
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_151
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_152
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_152 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_151 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_150 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_149 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_37 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_37;

architecture SYN_structural of MUX21_GENERIC_NBIT4_37 is

   component MUX21_145
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_146
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_147
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_148
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_148 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_147 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_146 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_145 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_36 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_36;

architecture SYN_structural of MUX21_GENERIC_NBIT4_36 is

   component MUX21_141
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_142
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_143
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_144
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_144 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_143 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_142 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_141 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_35 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_35;

architecture SYN_structural of MUX21_GENERIC_NBIT4_35 is

   component MUX21_137
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_138
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_139
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_140
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_140 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_139 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_138 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_137 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_34 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_34;

architecture SYN_structural of MUX21_GENERIC_NBIT4_34 is

   component MUX21_133
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_134
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_135
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_136
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_136 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_135 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_134 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_133 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_33 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_33;

architecture SYN_structural of MUX21_GENERIC_NBIT4_33 is

   component MUX21_129
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_130
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_131
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_132
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_132 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_131 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_130 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_129 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_32 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_32;

architecture SYN_structural of MUX21_GENERIC_NBIT4_32 is

   component MUX21_125
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_126
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_127
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_128
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_128 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_127 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_126 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_125 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_31 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_31;

architecture SYN_structural of MUX21_GENERIC_NBIT4_31 is

   component MUX21_121
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_122
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_123
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_124
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_124 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_123 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_122 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_121 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_30 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_30;

architecture SYN_structural of MUX21_GENERIC_NBIT4_30 is

   component MUX21_117
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_118
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_119
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_120
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_120 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_119 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_118 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_117 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_29 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_29;

architecture SYN_structural of MUX21_GENERIC_NBIT4_29 is

   component MUX21_113
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_114
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_115
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_116
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_116 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_115 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_114 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_113 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_28 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_28;

architecture SYN_structural of MUX21_GENERIC_NBIT4_28 is

   component MUX21_109
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_110
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_111
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_112
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_112 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_111 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_110 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_109 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_27 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_27;

architecture SYN_structural of MUX21_GENERIC_NBIT4_27 is

   component MUX21_105
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_106
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_107
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_108
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_108 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_107 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_106 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_105 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_26 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_26;

architecture SYN_structural of MUX21_GENERIC_NBIT4_26 is

   component MUX21_101
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_102
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_103
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_104
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_104 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_103 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_102 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_101 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_25 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_25;

architecture SYN_structural of MUX21_GENERIC_NBIT4_25 is

   component MUX21_97
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_98
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_99
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_100
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_100 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_99 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_98 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_97 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_24 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_24;

architecture SYN_structural of MUX21_GENERIC_NBIT4_24 is

   component MUX21_93
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_94
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_95
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_96
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_96 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_95 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_94 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_93 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_23 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_23;

architecture SYN_structural of MUX21_GENERIC_NBIT4_23 is

   component MUX21_89
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_90
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_91
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_92
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_92 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_91 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_90 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_89 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_22 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_22;

architecture SYN_structural of MUX21_GENERIC_NBIT4_22 is

   component MUX21_85
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_86
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_87
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_88
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_88 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_87 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_86 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_85 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_21 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_21;

architecture SYN_structural of MUX21_GENERIC_NBIT4_21 is

   component MUX21_81
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_82
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_83
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_84
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_84 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_83 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_82 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_81 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_20 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_20;

architecture SYN_structural of MUX21_GENERIC_NBIT4_20 is

   component MUX21_77
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_78
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_79
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_80
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_80 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_79 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_78 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_77 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_19 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_19;

architecture SYN_structural of MUX21_GENERIC_NBIT4_19 is

   component MUX21_73
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_74
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_75
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_76
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_76 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_75 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_74 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_73 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_18 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_18;

architecture SYN_structural of MUX21_GENERIC_NBIT4_18 is

   component MUX21_69
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_70
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_71
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_72
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_72 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_71 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_70 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_69 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_17 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_17;

architecture SYN_structural of MUX21_GENERIC_NBIT4_17 is

   component MUX21_65
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_66
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_67
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_68
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_68 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_67 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_66 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_65 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_16 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_16;

architecture SYN_structural of MUX21_GENERIC_NBIT4_16 is

   component MUX21_61
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_62
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_63
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_64
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_64 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_63 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_62 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_61 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_15 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_15;

architecture SYN_structural of MUX21_GENERIC_NBIT4_15 is

   component MUX21_57
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_58
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_59
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_60
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_60 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_59 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_58 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_57 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_14 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_14;

architecture SYN_structural of MUX21_GENERIC_NBIT4_14 is

   component MUX21_53
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_54
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_55
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_56
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_56 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_55 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_54 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_53 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_13 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_13;

architecture SYN_structural of MUX21_GENERIC_NBIT4_13 is

   component MUX21_49
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_50
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_51
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_52
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_52 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_51 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_50 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_49 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_12 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_12;

architecture SYN_structural of MUX21_GENERIC_NBIT4_12 is

   component MUX21_45
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_46
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_47
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_48
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_48 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_47 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_46 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_45 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_11 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_11;

architecture SYN_structural of MUX21_GENERIC_NBIT4_11 is

   component MUX21_41
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_42
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_43
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_44
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_44 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_43 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_42 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_41 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_10 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_10;

architecture SYN_structural of MUX21_GENERIC_NBIT4_10 is

   component MUX21_37
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_38
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_39
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_40
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_40 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_39 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_38 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_37 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_9 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_9;

architecture SYN_structural of MUX21_GENERIC_NBIT4_9 is

   component MUX21_33
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_34
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_35
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_36
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_36 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_35 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_34 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_33 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_8 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_8;

architecture SYN_structural of MUX21_GENERIC_NBIT4_8 is

   component MUX21_29
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_30
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_31
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_32
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_32 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_31 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_30 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_29 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_7;

architecture SYN_structural of MUX21_GENERIC_NBIT4_7 is

   component MUX21_25
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_26
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_27
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_28
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_28 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_27 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_26 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_25 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_6;

architecture SYN_structural of MUX21_GENERIC_NBIT4_6 is

   component MUX21_21
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_22
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_23
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_24
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_24 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_23 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_22 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_21 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_5;

architecture SYN_structural of MUX21_GENERIC_NBIT4_5 is

   component MUX21_17
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_18
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_19
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_20
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_20 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_19 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_18 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_17 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_4;

architecture SYN_structural of MUX21_GENERIC_NBIT4_4 is

   component MUX21_13
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_14
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_15
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_16
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_16 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_15 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_14 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_13 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_3;

architecture SYN_structural of MUX21_GENERIC_NBIT4_3 is

   component MUX21_9
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_10
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_11
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_12
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_12 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_11 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_10 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_9 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_2;

architecture SYN_structural of MUX21_GENERIC_NBIT4_2 is

   component MUX21_5
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_6
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_7
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_8
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_8 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_7 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_6 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_5 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_1;

architecture SYN_structural of MUX21_GENERIC_NBIT4_1 is

   component MUX21_1
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_2
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_3
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_4
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_4 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_3 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_2 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_1 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_127 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_127;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_127 is

   component FA_505
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_506
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_507
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_508
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_508 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_507 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_506 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_505 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_126 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_126;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_126 is

   component FA_501
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_502
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_503
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_504
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_504 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_503 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_502 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_501 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_125 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_125;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_125 is

   component FA_497
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_498
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_499
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_500
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_500 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_499 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_498 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_497 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_124 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_124;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_124 is

   component FA_493
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_494
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_495
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_496
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_496 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_495 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_494 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_493 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_123 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_123;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_123 is

   component FA_489
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_490
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_491
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_492
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_492 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_491 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_490 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_489 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_122 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_122;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_122 is

   component FA_485
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_486
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_487
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_488
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_488 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_487 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_486 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_485 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_121 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_121;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_121 is

   component FA_481
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_482
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_483
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_484
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_484 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_483 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_482 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_481 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_120 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_120;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_120 is

   component FA_477
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_478
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_479
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_480
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_480 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_479 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_478 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_477 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_119 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_119;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_119 is

   component FA_473
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_474
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_475
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_476
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_476 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_475 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_474 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_473 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_118 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_118;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_118 is

   component FA_469
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_470
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_471
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_472
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_472 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_471 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_470 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_469 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_117 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_117;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_117 is

   component FA_465
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_466
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_467
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_468
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_468 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_467 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_466 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_465 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_116 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_116;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_116 is

   component FA_461
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_462
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_463
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_464
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_464 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_463 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_462 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_461 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_115 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_115;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_115 is

   component FA_457
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_458
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_459
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_460
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_460 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_459 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_458 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_457 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_114 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_114;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_114 is

   component FA_453
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_454
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_455
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_456
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_456 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_455 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_454 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_453 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_113 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_113;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_113 is

   component FA_449
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_450
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_451
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_452
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_452 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_451 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_450 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_449 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_112 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_112;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_112 is

   component FA_445
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_446
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_447
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_448
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_448 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_447 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_446 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_445 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_111 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_111;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_111 is

   component FA_441
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_442
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_443
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_444
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_444 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_443 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_442 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_441 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_110 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_110;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_110 is

   component FA_437
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_438
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_439
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_440
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_440 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_439 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_438 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_437 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_109 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_109;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_109 is

   component FA_433
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_434
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_435
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_436
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_436 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_435 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_434 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_433 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_108 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_108;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_108 is

   component FA_429
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_430
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_431
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_432
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_432 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_431 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_430 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_429 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_107 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_107;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_107 is

   component FA_425
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_426
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_427
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_428
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_428 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_427 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_426 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_425 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_106 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_106;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_106 is

   component FA_421
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_422
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_423
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_424
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_424 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_423 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_422 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_421 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_105 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_105;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_105 is

   component FA_417
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_418
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_419
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_420
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_420 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_419 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_418 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_417 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_104 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_104;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_104 is

   component FA_413
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_414
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_415
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_416
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_416 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_415 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_414 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_413 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_103 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_103;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_103 is

   component FA_409
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_410
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_411
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_412
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_412 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_411 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_410 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_409 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_102 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_102;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_102 is

   component FA_405
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_406
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_407
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_408
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_408 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_407 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_406 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_405 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_101 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_101;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_101 is

   component FA_401
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_402
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_403
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_404
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_404 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_403 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_402 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_401 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_100 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_100;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_100 is

   component FA_397
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_398
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_399
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_400
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_400 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_399 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_398 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_397 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_99 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_99;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_99 is

   component FA_393
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_394
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_395
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_396
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_396 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_395 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_394 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_393 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_98 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_98;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_98 is

   component FA_389
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_390
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_391
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_392
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_392 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_391 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_390 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_389 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_97 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_97;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_97 is

   component FA_385
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_386
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_387
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_388
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_388 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_387 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_386 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_385 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_96 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_96;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_96 is

   component FA_381
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_382
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_383
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_384
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_384 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_383 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_382 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_381 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_95 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_95;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_95 is

   component FA_377
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_378
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_379
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_380
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_380 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_379 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_378 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_377 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_94 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_94;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_94 is

   component FA_373
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_374
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_375
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_376
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_376 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_375 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_374 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_373 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_93 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_93;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_93 is

   component FA_369
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_370
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_371
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_372
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_372 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_371 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_370 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_369 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_92 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_92;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_92 is

   component FA_365
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_366
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_367
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_368
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_368 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_367 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_366 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_365 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_91 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_91;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_91 is

   component FA_361
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_362
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_363
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_364
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_364 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_363 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_362 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_361 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_90 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_90;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_90 is

   component FA_357
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_358
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_359
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_360
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_360 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_359 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_358 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_357 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_89 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_89;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_89 is

   component FA_353
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_354
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_355
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_356
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_356 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_355 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_354 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_353 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_88 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_88;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_88 is

   component FA_349
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_350
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_351
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_352
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_352 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_351 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_350 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_349 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_87 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_87;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_87 is

   component FA_345
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_346
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_347
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_348
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_348 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_347 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_346 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_345 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_86 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_86;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_86 is

   component FA_341
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_342
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_343
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_344
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_344 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_343 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_342 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_341 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_85 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_85;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_85 is

   component FA_337
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_338
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_339
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_340
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_340 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_339 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_338 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_337 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_84 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_84;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_84 is

   component FA_333
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_334
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_335
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_336
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_336 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_335 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_334 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_333 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_83 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_83;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_83 is

   component FA_329
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_330
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_331
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_332
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_332 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_331 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_330 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_329 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_82 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_82;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_82 is

   component FA_325
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_326
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_327
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_328
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_328 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_327 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_326 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_325 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_81 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_81;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_81 is

   component FA_321
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_322
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_323
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_324
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_324 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_323 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_322 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_321 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_80 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_80;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_80 is

   component FA_317
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_318
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_319
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_320
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_320 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_319 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_318 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_317 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_79 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_79;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_79 is

   component FA_313
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_314
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_315
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_316
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_316 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_315 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_314 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_313 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_78 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_78;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_78 is

   component FA_309
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_310
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_311
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_312
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_312 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_311 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_310 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_309 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_77 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_77;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_77 is

   component FA_305
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_306
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_307
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_308
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_308 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_307 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_306 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_305 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_76 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_76;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_76 is

   component FA_301
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_302
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_303
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_304
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_304 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_303 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_302 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_301 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_75 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_75;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_75 is

   component FA_297
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_298
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_299
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_300
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_300 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_299 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_298 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_297 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_74 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_74;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_74 is

   component FA_293
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_294
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_295
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_296
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_296 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_295 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_294 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_293 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_73 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_73;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_73 is

   component FA_289
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_290
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_291
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_292
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_292 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_291 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_290 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_289 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_72 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_72;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_72 is

   component FA_285
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_286
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_287
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_288
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_288 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_287 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_286 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_285 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_71 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_71;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_71 is

   component FA_281
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_282
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_283
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_284
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_284 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_283 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_282 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_281 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_70 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_70;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_70 is

   component FA_277
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_278
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_279
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_280
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_280 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_279 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_278 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_277 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_69 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_69;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_69 is

   component FA_273
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_274
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_275
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_276
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_276 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_275 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_274 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_273 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_68 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_68;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_68 is

   component FA_269
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_270
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_271
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_272
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_272 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_271 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_270 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_269 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_67 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_67;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_67 is

   component FA_265
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_266
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_267
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_268
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_268 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_267 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_266 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_265 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_66 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_66;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_66 is

   component FA_261
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_262
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_263
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_264
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_264 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_263 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_262 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_261 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_65 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_65;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_65 is

   component FA_257
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_258
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_259
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_260
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_260 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_259 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_258 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_257 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_64 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_64;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_64 is

   component FA_253
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_254
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_255
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_256
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_256 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_255 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_254 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_253 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_63 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_63;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_63 is

   component FA_249
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_250
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_251
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_252
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_252 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_251 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_250 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_249 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_62 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_62;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_62 is

   component FA_245
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_246
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_247
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_248
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_248 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_247 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_246 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_245 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_61 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_61;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_61 is

   component FA_241
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_242
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_243
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_244
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_244 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_243 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_242 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_241 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_60 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_60;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_60 is

   component FA_237
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_238
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_239
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_240
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_240 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_239 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_238 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_237 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_59 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_59;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_59 is

   component FA_233
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_234
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_235
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_236
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_236 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_235 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_234 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_233 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_58 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_58;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_58 is

   component FA_229
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_230
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_231
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_232
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_232 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_231 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_230 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_229 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_57 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_57;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_57 is

   component FA_225
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_226
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_227
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_228
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_228 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_227 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_226 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_225 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_56 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_56;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_56 is

   component FA_221
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_222
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_223
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_224
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_224 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_223 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_222 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_221 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_55 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_55;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_55 is

   component FA_217
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_218
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_219
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_220
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_220 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_219 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_218 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_217 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_54 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_54;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_54 is

   component FA_213
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_214
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_215
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_216
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_216 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_215 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_214 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_213 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_53 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_53;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_53 is

   component FA_209
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_210
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_211
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_212
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_212 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_211 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_210 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_209 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_52 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_52;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_52 is

   component FA_205
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_206
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_207
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_208
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_208 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_207 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_206 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_205 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_51 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_51;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_51 is

   component FA_201
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_202
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_203
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_204
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_204 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_203 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_202 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_201 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_50 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_50;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_50 is

   component FA_197
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_198
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_199
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_200
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_200 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_199 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_198 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_197 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_49 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_49;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_49 is

   component FA_193
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_194
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_195
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_196
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_196 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_195 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_194 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_193 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_48 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_48;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_48 is

   component FA_189
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_190
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_191
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_192
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_192 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_191 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_190 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_189 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_47 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_47;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_47 is

   component FA_185
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_186
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_187
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_188
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_188 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_187 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_186 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_185 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_46 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_46;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_46 is

   component FA_181
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_182
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_183
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_184
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_184 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_183 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_182 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_181 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_45 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_45;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_45 is

   component FA_177
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_178
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_179
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_180
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_180 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_179 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_178 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_177 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_44 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_44;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_44 is

   component FA_173
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_174
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_175
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_176
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_176 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_175 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_174 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_173 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_43 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_43;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_43 is

   component FA_169
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_170
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_171
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_172
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_172 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_171 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_170 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_169 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_42 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_42;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_42 is

   component FA_165
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_166
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_167
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_168
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_168 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_167 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_166 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_165 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_41 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_41;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_41 is

   component FA_161
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_162
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_163
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_164
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_164 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_163 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_162 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_161 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_40 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_40;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_40 is

   component FA_157
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_158
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_159
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_160
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_160 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_159 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_158 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_157 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_39 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_39;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_39 is

   component FA_153
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_154
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_155
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_156
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_156 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_155 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_154 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_153 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_38 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_38;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_38 is

   component FA_149
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_150
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_151
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_152
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_152 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_151 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_150 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_149 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_37 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_37;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_37 is

   component FA_145
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_146
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_147
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_148
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_148 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_147 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_146 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_145 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_36 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_36;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_36 is

   component FA_141
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_142
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_143
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_144
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_144 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_143 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_142 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_141 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_35 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_35;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_35 is

   component FA_137
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_138
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_139
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_140
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_140 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_139 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_138 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_137 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_34 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_34;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_34 is

   component FA_133
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_134
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_135
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_136
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_136 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_135 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_134 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_133 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_33 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_33;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_33 is

   component FA_129
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_130
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_131
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_132
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_132 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_131 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_130 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_129 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_32 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_32;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_32 is

   component FA_125
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_126
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_127
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_128
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_128 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_127 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_126 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_125 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_31 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_31;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_31 is

   component FA_121
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_122
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_123
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_124
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_124 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_123 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_122 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_121 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_30 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_30;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_30 is

   component FA_117
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_118
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_119
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_120
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_120 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_119 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_118 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_117 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_29 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_29;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_29 is

   component FA_113
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_114
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_115
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_116
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_116 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_115 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_114 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_113 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_28 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_28;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_28 is

   component FA_109
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_110
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_111
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_112
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_112 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_111 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_110 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_109 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_27 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_27;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_27 is

   component FA_105
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_106
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_107
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_108
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_108 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_107 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_106 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_105 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_26 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_26;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_26 is

   component FA_101
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_102
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_103
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_104
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_104 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_103 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_102 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_101 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_25 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_25;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_25 is

   component FA_97
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_98
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_99
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_100
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_100 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_99 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_98 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_97 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_24 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_24;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_24 is

   component FA_93
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_94
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_95
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_96
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_96 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_95 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_94 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_93 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_23 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_23;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_23 is

   component FA_89
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_90
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_91
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_92
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_92 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_91 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_90 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_89 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_22 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_22;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_22 is

   component FA_85
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_86
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_87
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_88
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_88 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_87 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_86 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_85 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_21 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_21;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_21 is

   component FA_81
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_82
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_83
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_84
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_84 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_83 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_82 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_81 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_20 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_20;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_20 is

   component FA_77
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_78
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_79
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_80
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_80 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_79 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_78 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_77 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_19 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_19;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_19 is

   component FA_73
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_74
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_75
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_76
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_76 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_75 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_74 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_73 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_18 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_18;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_18 is

   component FA_69
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_70
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_71
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_72
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_72 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_71 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_70 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_69 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_17 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_17;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_17 is

   component FA_65
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_66
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_67
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_68
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_68 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_67 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_66 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_65 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_16 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_16;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_16 is

   component FA_61
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_62
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_63
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_64
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_64 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_63 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_62 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_61 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_15 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_15;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_15 is

   component FA_57
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_58
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_59
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_60
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_60 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_59 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_58 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_57 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_14 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_14;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_14 is

   component FA_53
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_54
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_55
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_56
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_56 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_55 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_54 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_53 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_13 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_13;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_13 is

   component FA_49
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_50
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_51
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_52
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_52 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_51 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_50 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_49 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_12 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_12;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_12 is

   component FA_45
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_46
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_47
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_48
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_48 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_47 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_46 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_45 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_11 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_11;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_11 is

   component FA_41
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_42
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_43
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_44
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_44 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_43 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_42 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_41 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_10 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_10;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_10 is

   component FA_37
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_38
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_39
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_40
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_40 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_39 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_38 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_37 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_9 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_9;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_9 is

   component FA_33
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_34
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_35
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_36
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_36 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_35 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_34 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_33 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_8 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_8;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_8 is

   component FA_29
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_30
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_31
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_32
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_32 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_31 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_30 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_29 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_7;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_7 is

   component FA_25
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_26
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_27
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_28
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_28 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_27 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_26 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_25 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_6;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_6 is

   component FA_21
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_22
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_23
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_24
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_24 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_23 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_22 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_21 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_5;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_5 is

   component FA_17
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_18
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_19
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_20
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_20 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_19 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_18 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_17 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_4;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_4 is

   component FA_13
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_14
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_15
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_16
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_16 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_15 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_14 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_13 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_3;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_3 is

   component FA_9
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_10
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_11
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_12
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_12 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_11 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_10 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_9 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_2;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_2 is

   component FA_5
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_6
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_7
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_8
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_8 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_7 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_6 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_5 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_1;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_1 is

   component FA_1
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_3
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_4
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_4 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_3 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   FAI_3 : FA_2 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   FAI_4 : FA_1 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity P4_ADDER_NBIT64_2 is

   port( A, B : in std_logic_vector (63 downto 0);  Cin : in std_logic;  S : 
         out std_logic_vector (63 downto 0);  Cout, ovf : out std_logic);

end P4_ADDER_NBIT64_2;

architecture SYN_STRUCTURAL of P4_ADDER_NBIT64_2 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component sum_generator_n_bit64_n_CSB16_2
      port( A, B : in std_logic_vector (63 downto 0);  C_in : in 
            std_logic_vector (15 downto 0);  S : out std_logic_vector (63 
            downto 0));
   end component;
   
   component CARRY_GENERATOR_NBIT64_NBIT_PER_BLOCK4_2
      port( A, B : in std_logic_vector (63 downto 0);  Cin : in std_logic;  Co 
            : out std_logic_vector (15 downto 0));
   end component;
   
   component my_xor_65
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_66
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_67
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_68
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_69
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_70
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_71
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_72
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_73
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_74
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_75
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_76
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_77
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_78
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_79
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_80
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_81
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_82
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_83
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_84
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_85
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_86
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_87
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_88
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_89
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_90
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_91
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_92
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_93
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_94
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_95
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_96
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_97
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_98
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_99
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_100
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_101
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_102
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_103
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_104
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_105
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_106
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_107
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_108
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_109
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_110
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_111
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_112
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_113
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_114
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_115
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_116
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_117
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_118
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_119
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_120
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_121
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_122
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_123
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_124
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_125
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_126
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_127
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_128
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal S_63_port, S_62_port, S_61_port, S_60_port, S_59_port, S_58_port, 
      S_57_port, S_56_port, S_55_port, S_54_port, S_53_port, S_52_port, 
      S_51_port, S_50_port, S_49_port, S_48_port, S_47_port, S_46_port, 
      S_45_port, S_44_port, S_43_port, S_42_port, S_41_port, S_40_port, 
      S_39_port, S_38_port, S_37_port, S_36_port, S_35_port, S_34_port, 
      S_33_port, S_32_port, S_31_port, S_30_port, S_29_port, S_28_port, 
      S_27_port, S_26_port, S_25_port, S_24_port, S_23_port, S_22_port, 
      S_21_port, S_20_port, S_19_port, S_18_port, S_17_port, S_16_port, 
      S_15_port, S_14_port, S_13_port, S_12_port, S_11_port, S_10_port, 
      S_9_port, S_8_port, S_7_port, S_6_port, S_5_port, S_4_port, S_3_port, 
      S_2_port, S_1_port, S_0_port, xor_b_63_port, xor_b_62_port, xor_b_61_port
      , xor_b_60_port, xor_b_59_port, xor_b_58_port, xor_b_57_port, 
      xor_b_56_port, xor_b_55_port, xor_b_54_port, xor_b_53_port, xor_b_52_port
      , xor_b_51_port, xor_b_50_port, xor_b_49_port, xor_b_48_port, 
      xor_b_47_port, xor_b_46_port, xor_b_45_port, xor_b_44_port, xor_b_43_port
      , xor_b_42_port, xor_b_41_port, xor_b_40_port, xor_b_39_port, 
      xor_b_38_port, xor_b_37_port, xor_b_36_port, xor_b_35_port, xor_b_34_port
      , xor_b_33_port, xor_b_32_port, xor_b_31_port, xor_b_30_port, 
      xor_b_29_port, xor_b_28_port, xor_b_27_port, xor_b_26_port, xor_b_25_port
      , xor_b_24_port, xor_b_23_port, xor_b_22_port, xor_b_21_port, 
      xor_b_20_port, xor_b_19_port, xor_b_18_port, xor_b_17_port, xor_b_16_port
      , xor_b_15_port, xor_b_14_port, xor_b_13_port, xor_b_12_port, 
      xor_b_11_port, xor_b_10_port, xor_b_9_port, xor_b_8_port, xor_b_7_port, 
      xor_b_6_port, xor_b_5_port, xor_b_4_port, xor_b_3_port, xor_b_2_port, 
      xor_b_1_port, xor_b_0_port, carry_14_port, carry_13_port, carry_12_port, 
      carry_11_port, carry_10_port, carry_9_port, carry_8_port, carry_7_port, 
      carry_6_port, carry_5_port, carry_4_port, carry_3_port, carry_2_port, 
      carry_1_port, carry_0_port, n3, n4 : std_logic;

begin
   S <= ( S_63_port, S_62_port, S_61_port, S_60_port, S_59_port, S_58_port, 
      S_57_port, S_56_port, S_55_port, S_54_port, S_53_port, S_52_port, 
      S_51_port, S_50_port, S_49_port, S_48_port, S_47_port, S_46_port, 
      S_45_port, S_44_port, S_43_port, S_42_port, S_41_port, S_40_port, 
      S_39_port, S_38_port, S_37_port, S_36_port, S_35_port, S_34_port, 
      S_33_port, S_32_port, S_31_port, S_30_port, S_29_port, S_28_port, 
      S_27_port, S_26_port, S_25_port, S_24_port, S_23_port, S_22_port, 
      S_21_port, S_20_port, S_19_port, S_18_port, S_17_port, S_16_port, 
      S_15_port, S_14_port, S_13_port, S_12_port, S_11_port, S_10_port, 
      S_9_port, S_8_port, S_7_port, S_6_port, S_5_port, S_4_port, S_3_port, 
      S_2_port, S_1_port, S_0_port );
   
   U3 : XOR2_X1 port map( A => xor_b_63_port, B => A(63), Z => n3);
   bc_xor_63 : my_xor_128 port map( A => B(63), B => Cin, xor_out => 
                           xor_b_63_port);
   bc_xor_62 : my_xor_127 port map( A => B(62), B => Cin, xor_out => 
                           xor_b_62_port);
   bc_xor_61 : my_xor_126 port map( A => B(61), B => Cin, xor_out => 
                           xor_b_61_port);
   bc_xor_60 : my_xor_125 port map( A => B(60), B => Cin, xor_out => 
                           xor_b_60_port);
   bc_xor_59 : my_xor_124 port map( A => B(59), B => Cin, xor_out => 
                           xor_b_59_port);
   bc_xor_58 : my_xor_123 port map( A => B(58), B => Cin, xor_out => 
                           xor_b_58_port);
   bc_xor_57 : my_xor_122 port map( A => B(57), B => Cin, xor_out => 
                           xor_b_57_port);
   bc_xor_56 : my_xor_121 port map( A => B(56), B => Cin, xor_out => 
                           xor_b_56_port);
   bc_xor_55 : my_xor_120 port map( A => B(55), B => Cin, xor_out => 
                           xor_b_55_port);
   bc_xor_54 : my_xor_119 port map( A => B(54), B => Cin, xor_out => 
                           xor_b_54_port);
   bc_xor_53 : my_xor_118 port map( A => B(53), B => Cin, xor_out => 
                           xor_b_53_port);
   bc_xor_52 : my_xor_117 port map( A => B(52), B => Cin, xor_out => 
                           xor_b_52_port);
   bc_xor_51 : my_xor_116 port map( A => B(51), B => Cin, xor_out => 
                           xor_b_51_port);
   bc_xor_50 : my_xor_115 port map( A => B(50), B => Cin, xor_out => 
                           xor_b_50_port);
   bc_xor_49 : my_xor_114 port map( A => B(49), B => Cin, xor_out => 
                           xor_b_49_port);
   bc_xor_48 : my_xor_113 port map( A => B(48), B => Cin, xor_out => 
                           xor_b_48_port);
   bc_xor_47 : my_xor_112 port map( A => B(47), B => Cin, xor_out => 
                           xor_b_47_port);
   bc_xor_46 : my_xor_111 port map( A => B(46), B => Cin, xor_out => 
                           xor_b_46_port);
   bc_xor_45 : my_xor_110 port map( A => B(45), B => Cin, xor_out => 
                           xor_b_45_port);
   bc_xor_44 : my_xor_109 port map( A => B(44), B => Cin, xor_out => 
                           xor_b_44_port);
   bc_xor_43 : my_xor_108 port map( A => B(43), B => Cin, xor_out => 
                           xor_b_43_port);
   bc_xor_42 : my_xor_107 port map( A => B(42), B => Cin, xor_out => 
                           xor_b_42_port);
   bc_xor_41 : my_xor_106 port map( A => B(41), B => Cin, xor_out => 
                           xor_b_41_port);
   bc_xor_40 : my_xor_105 port map( A => B(40), B => Cin, xor_out => 
                           xor_b_40_port);
   bc_xor_39 : my_xor_104 port map( A => B(39), B => Cin, xor_out => 
                           xor_b_39_port);
   bc_xor_38 : my_xor_103 port map( A => B(38), B => Cin, xor_out => 
                           xor_b_38_port);
   bc_xor_37 : my_xor_102 port map( A => B(37), B => Cin, xor_out => 
                           xor_b_37_port);
   bc_xor_36 : my_xor_101 port map( A => B(36), B => Cin, xor_out => 
                           xor_b_36_port);
   bc_xor_35 : my_xor_100 port map( A => B(35), B => Cin, xor_out => 
                           xor_b_35_port);
   bc_xor_34 : my_xor_99 port map( A => B(34), B => Cin, xor_out => 
                           xor_b_34_port);
   bc_xor_33 : my_xor_98 port map( A => B(33), B => Cin, xor_out => 
                           xor_b_33_port);
   bc_xor_32 : my_xor_97 port map( A => B(32), B => Cin, xor_out => 
                           xor_b_32_port);
   bc_xor_31 : my_xor_96 port map( A => B(31), B => Cin, xor_out => 
                           xor_b_31_port);
   bc_xor_30 : my_xor_95 port map( A => B(30), B => Cin, xor_out => 
                           xor_b_30_port);
   bc_xor_29 : my_xor_94 port map( A => B(29), B => Cin, xor_out => 
                           xor_b_29_port);
   bc_xor_28 : my_xor_93 port map( A => B(28), B => Cin, xor_out => 
                           xor_b_28_port);
   bc_xor_27 : my_xor_92 port map( A => B(27), B => Cin, xor_out => 
                           xor_b_27_port);
   bc_xor_26 : my_xor_91 port map( A => B(26), B => Cin, xor_out => 
                           xor_b_26_port);
   bc_xor_25 : my_xor_90 port map( A => B(25), B => Cin, xor_out => 
                           xor_b_25_port);
   bc_xor_24 : my_xor_89 port map( A => B(24), B => Cin, xor_out => 
                           xor_b_24_port);
   bc_xor_23 : my_xor_88 port map( A => B(23), B => Cin, xor_out => 
                           xor_b_23_port);
   bc_xor_22 : my_xor_87 port map( A => B(22), B => Cin, xor_out => 
                           xor_b_22_port);
   bc_xor_21 : my_xor_86 port map( A => B(21), B => Cin, xor_out => 
                           xor_b_21_port);
   bc_xor_20 : my_xor_85 port map( A => B(20), B => Cin, xor_out => 
                           xor_b_20_port);
   bc_xor_19 : my_xor_84 port map( A => B(19), B => Cin, xor_out => 
                           xor_b_19_port);
   bc_xor_18 : my_xor_83 port map( A => B(18), B => Cin, xor_out => 
                           xor_b_18_port);
   bc_xor_17 : my_xor_82 port map( A => B(17), B => Cin, xor_out => 
                           xor_b_17_port);
   bc_xor_16 : my_xor_81 port map( A => B(16), B => Cin, xor_out => 
                           xor_b_16_port);
   bc_xor_15 : my_xor_80 port map( A => B(15), B => Cin, xor_out => 
                           xor_b_15_port);
   bc_xor_14 : my_xor_79 port map( A => B(14), B => Cin, xor_out => 
                           xor_b_14_port);
   bc_xor_13 : my_xor_78 port map( A => B(13), B => Cin, xor_out => 
                           xor_b_13_port);
   bc_xor_12 : my_xor_77 port map( A => B(12), B => Cin, xor_out => 
                           xor_b_12_port);
   bc_xor_11 : my_xor_76 port map( A => B(11), B => Cin, xor_out => 
                           xor_b_11_port);
   bc_xor_10 : my_xor_75 port map( A => B(10), B => Cin, xor_out => 
                           xor_b_10_port);
   bc_xor_9 : my_xor_74 port map( A => B(9), B => Cin, xor_out => xor_b_9_port)
                           ;
   bc_xor_8 : my_xor_73 port map( A => B(8), B => Cin, xor_out => xor_b_8_port)
                           ;
   bc_xor_7 : my_xor_72 port map( A => B(7), B => Cin, xor_out => xor_b_7_port)
                           ;
   bc_xor_6 : my_xor_71 port map( A => B(6), B => Cin, xor_out => xor_b_6_port)
                           ;
   bc_xor_5 : my_xor_70 port map( A => B(5), B => Cin, xor_out => xor_b_5_port)
                           ;
   bc_xor_4 : my_xor_69 port map( A => B(4), B => Cin, xor_out => xor_b_4_port)
                           ;
   bc_xor_3 : my_xor_68 port map( A => B(3), B => Cin, xor_out => xor_b_3_port)
                           ;
   bc_xor_2 : my_xor_67 port map( A => B(2), B => Cin, xor_out => xor_b_2_port)
                           ;
   bc_xor_1 : my_xor_66 port map( A => B(1), B => Cin, xor_out => xor_b_1_port)
                           ;
   bc_xor_0 : my_xor_65 port map( A => B(0), B => Cin, xor_out => xor_b_0_port)
                           ;
   CG : CARRY_GENERATOR_NBIT64_NBIT_PER_BLOCK4_2 port map( A(63) => A(63), 
                           A(62) => A(62), A(61) => A(61), A(60) => A(60), 
                           A(59) => A(59), A(58) => A(58), A(57) => A(57), 
                           A(56) => A(56), A(55) => A(55), A(54) => A(54), 
                           A(53) => A(53), A(52) => A(52), A(51) => A(51), 
                           A(50) => A(50), A(49) => A(49), A(48) => A(48), 
                           A(47) => A(47), A(46) => A(46), A(45) => A(45), 
                           A(44) => A(44), A(43) => A(43), A(42) => A(42), 
                           A(41) => A(41), A(40) => A(40), A(39) => A(39), 
                           A(38) => A(38), A(37) => A(37), A(36) => A(36), 
                           A(35) => A(35), A(34) => A(34), A(33) => A(33), 
                           A(32) => A(32), A(31) => A(31), A(30) => A(30), 
                           A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(63) => xor_b_63_port, B(62) =>
                           xor_b_62_port, B(61) => xor_b_61_port, B(60) => 
                           xor_b_60_port, B(59) => xor_b_59_port, B(58) => 
                           xor_b_58_port, B(57) => xor_b_57_port, B(56) => 
                           xor_b_56_port, B(55) => xor_b_55_port, B(54) => 
                           xor_b_54_port, B(53) => xor_b_53_port, B(52) => 
                           xor_b_52_port, B(51) => xor_b_51_port, B(50) => 
                           xor_b_50_port, B(49) => xor_b_49_port, B(48) => 
                           xor_b_48_port, B(47) => xor_b_47_port, B(46) => 
                           xor_b_46_port, B(45) => xor_b_45_port, B(44) => 
                           xor_b_44_port, B(43) => xor_b_43_port, B(42) => 
                           xor_b_42_port, B(41) => xor_b_41_port, B(40) => 
                           xor_b_40_port, B(39) => xor_b_39_port, B(38) => 
                           xor_b_38_port, B(37) => xor_b_37_port, B(36) => 
                           xor_b_36_port, B(35) => xor_b_35_port, B(34) => 
                           xor_b_34_port, B(33) => xor_b_33_port, B(32) => 
                           xor_b_32_port, B(31) => xor_b_31_port, B(30) => 
                           xor_b_30_port, B(29) => xor_b_29_port, B(28) => 
                           xor_b_28_port, B(27) => xor_b_27_port, B(26) => 
                           xor_b_26_port, B(25) => xor_b_25_port, B(24) => 
                           xor_b_24_port, B(23) => xor_b_23_port, B(22) => 
                           xor_b_22_port, B(21) => xor_b_21_port, B(20) => 
                           xor_b_20_port, B(19) => xor_b_19_port, B(18) => 
                           xor_b_18_port, B(17) => xor_b_17_port, B(16) => 
                           xor_b_16_port, B(15) => xor_b_15_port, B(14) => 
                           xor_b_14_port, B(13) => xor_b_13_port, B(12) => 
                           xor_b_12_port, B(11) => xor_b_11_port, B(10) => 
                           xor_b_10_port, B(9) => xor_b_9_port, B(8) => 
                           xor_b_8_port, B(7) => xor_b_7_port, B(6) => 
                           xor_b_6_port, B(5) => xor_b_5_port, B(4) => 
                           xor_b_4_port, B(3) => xor_b_3_port, B(2) => 
                           xor_b_2_port, B(1) => xor_b_1_port, B(0) => 
                           xor_b_0_port, Cin => Cin, Co(15) => Cout, Co(14) => 
                           carry_14_port, Co(13) => carry_13_port, Co(12) => 
                           carry_12_port, Co(11) => carry_11_port, Co(10) => 
                           carry_10_port, Co(9) => carry_9_port, Co(8) => 
                           carry_8_port, Co(7) => carry_7_port, Co(6) => 
                           carry_6_port, Co(5) => carry_5_port, Co(4) => 
                           carry_4_port, Co(3) => carry_3_port, Co(2) => 
                           carry_2_port, Co(1) => carry_1_port, Co(0) => 
                           carry_0_port);
   SG : sum_generator_n_bit64_n_CSB16_2 port map( A(63) => A(63), A(62) => 
                           A(62), A(61) => A(61), A(60) => A(60), A(59) => 
                           A(59), A(58) => A(58), A(57) => A(57), A(56) => 
                           A(56), A(55) => A(55), A(54) => A(54), A(53) => 
                           A(53), A(52) => A(52), A(51) => A(51), A(50) => 
                           A(50), A(49) => A(49), A(48) => A(48), A(47) => 
                           A(47), A(46) => A(46), A(45) => A(45), A(44) => 
                           A(44), A(43) => A(43), A(42) => A(42), A(41) => 
                           A(41), A(40) => A(40), A(39) => A(39), A(38) => 
                           A(38), A(37) => A(37), A(36) => A(36), A(35) => 
                           A(35), A(34) => A(34), A(33) => A(33), A(32) => 
                           A(32), A(31) => A(31), A(30) => A(30), A(29) => 
                           A(29), A(28) => A(28), A(27) => A(27), A(26) => 
                           A(26), A(25) => A(25), A(24) => A(24), A(23) => 
                           A(23), A(22) => A(22), A(21) => A(21), A(20) => 
                           A(20), A(19) => A(19), A(18) => A(18), A(17) => 
                           A(17), A(16) => A(16), A(15) => A(15), A(14) => 
                           A(14), A(13) => A(13), A(12) => A(12), A(11) => 
                           A(11), A(10) => A(10), A(9) => A(9), A(8) => A(8), 
                           A(7) => A(7), A(6) => A(6), A(5) => A(5), A(4) => 
                           A(4), A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(63) => xor_b_63_port, B(62) => 
                           xor_b_62_port, B(61) => xor_b_61_port, B(60) => 
                           xor_b_60_port, B(59) => xor_b_59_port, B(58) => 
                           xor_b_58_port, B(57) => xor_b_57_port, B(56) => 
                           xor_b_56_port, B(55) => xor_b_55_port, B(54) => 
                           xor_b_54_port, B(53) => xor_b_53_port, B(52) => 
                           xor_b_52_port, B(51) => xor_b_51_port, B(50) => 
                           xor_b_50_port, B(49) => xor_b_49_port, B(48) => 
                           xor_b_48_port, B(47) => xor_b_47_port, B(46) => 
                           xor_b_46_port, B(45) => xor_b_45_port, B(44) => 
                           xor_b_44_port, B(43) => xor_b_43_port, B(42) => 
                           xor_b_42_port, B(41) => xor_b_41_port, B(40) => 
                           xor_b_40_port, B(39) => xor_b_39_port, B(38) => 
                           xor_b_38_port, B(37) => xor_b_37_port, B(36) => 
                           xor_b_36_port, B(35) => xor_b_35_port, B(34) => 
                           xor_b_34_port, B(33) => xor_b_33_port, B(32) => 
                           xor_b_32_port, B(31) => xor_b_31_port, B(30) => 
                           xor_b_30_port, B(29) => xor_b_29_port, B(28) => 
                           xor_b_28_port, B(27) => xor_b_27_port, B(26) => 
                           xor_b_26_port, B(25) => xor_b_25_port, B(24) => 
                           xor_b_24_port, B(23) => xor_b_23_port, B(22) => 
                           xor_b_22_port, B(21) => xor_b_21_port, B(20) => 
                           xor_b_20_port, B(19) => xor_b_19_port, B(18) => 
                           xor_b_18_port, B(17) => xor_b_17_port, B(16) => 
                           xor_b_16_port, B(15) => xor_b_15_port, B(14) => 
                           xor_b_14_port, B(13) => xor_b_13_port, B(12) => 
                           xor_b_12_port, B(11) => xor_b_11_port, B(10) => 
                           xor_b_10_port, B(9) => xor_b_9_port, B(8) => 
                           xor_b_8_port, B(7) => xor_b_7_port, B(6) => 
                           xor_b_6_port, B(5) => xor_b_5_port, B(4) => 
                           xor_b_4_port, B(3) => xor_b_3_port, B(2) => 
                           xor_b_2_port, B(1) => xor_b_1_port, B(0) => 
                           xor_b_0_port, C_in(15) => carry_14_port, C_in(14) =>
                           carry_13_port, C_in(13) => carry_12_port, C_in(12) 
                           => carry_11_port, C_in(11) => carry_10_port, 
                           C_in(10) => carry_9_port, C_in(9) => carry_8_port, 
                           C_in(8) => carry_7_port, C_in(7) => carry_6_port, 
                           C_in(6) => carry_5_port, C_in(5) => carry_4_port, 
                           C_in(4) => carry_3_port, C_in(3) => carry_2_port, 
                           C_in(2) => carry_1_port, C_in(1) => carry_0_port, 
                           C_in(0) => Cin, S(63) => S_63_port, S(62) => 
                           S_62_port, S(61) => S_61_port, S(60) => S_60_port, 
                           S(59) => S_59_port, S(58) => S_58_port, S(57) => 
                           S_57_port, S(56) => S_56_port, S(55) => S_55_port, 
                           S(54) => S_54_port, S(53) => S_53_port, S(52) => 
                           S_52_port, S(51) => S_51_port, S(50) => S_50_port, 
                           S(49) => S_49_port, S(48) => S_48_port, S(47) => 
                           S_47_port, S(46) => S_46_port, S(45) => S_45_port, 
                           S(44) => S_44_port, S(43) => S_43_port, S(42) => 
                           S_42_port, S(41) => S_41_port, S(40) => S_40_port, 
                           S(39) => S_39_port, S(38) => S_38_port, S(37) => 
                           S_37_port, S(36) => S_36_port, S(35) => S_35_port, 
                           S(34) => S_34_port, S(33) => S_33_port, S(32) => 
                           S_32_port, S(31) => S_31_port, S(30) => S_30_port, 
                           S(29) => S_29_port, S(28) => S_28_port, S(27) => 
                           S_27_port, S(26) => S_26_port, S(25) => S_25_port, 
                           S(24) => S_24_port, S(23) => S_23_port, S(22) => 
                           S_22_port, S(21) => S_21_port, S(20) => S_20_port, 
                           S(19) => S_19_port, S(18) => S_18_port, S(17) => 
                           S_17_port, S(16) => S_16_port, S(15) => S_15_port, 
                           S(14) => S_14_port, S(13) => S_13_port, S(12) => 
                           S_12_port, S(11) => S_11_port, S(10) => S_10_port, 
                           S(9) => S_9_port, S(8) => S_8_port, S(7) => S_7_port
                           , S(6) => S_6_port, S(5) => S_5_port, S(4) => 
                           S_4_port, S(3) => S_3_port, S(2) => S_2_port, S(1) 
                           => S_1_port, S(0) => S_0_port);
   U1 : NOR2_X1 port map( A1 => n4, A2 => n3, ZN => ovf);
   U2 : XNOR2_X1 port map( A => A(63), B => S_63_port, ZN => n4);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity P4_ADDER_NBIT64_1 is

   port( A, B : in std_logic_vector (63 downto 0);  Cin : in std_logic;  S : 
         out std_logic_vector (63 downto 0);  Cout, ovf : out std_logic);

end P4_ADDER_NBIT64_1;

architecture SYN_STRUCTURAL of P4_ADDER_NBIT64_1 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component sum_generator_n_bit64_n_CSB16_1
      port( A, B : in std_logic_vector (63 downto 0);  C_in : in 
            std_logic_vector (15 downto 0);  S : out std_logic_vector (63 
            downto 0));
   end component;
   
   component CARRY_GENERATOR_NBIT64_NBIT_PER_BLOCK4_1
      port( A, B : in std_logic_vector (63 downto 0);  Cin : in std_logic;  Co 
            : out std_logic_vector (15 downto 0));
   end component;
   
   component my_xor_1
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_2
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_3
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_4
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_5
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_6
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_7
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_8
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_9
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_10
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_11
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_12
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_13
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_14
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_15
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_16
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_17
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_18
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_19
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_20
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_21
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_22
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_23
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_24
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_25
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_26
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_27
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_28
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_29
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_30
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_31
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_32
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_33
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_34
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_35
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_36
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_37
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_38
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_39
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_40
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_41
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_42
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_43
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_44
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_45
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_46
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_47
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_48
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_49
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_50
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_51
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_52
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_53
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_54
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_55
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_56
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_57
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_58
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_59
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_60
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_61
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_62
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_63
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_64
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal S_63_port, S_62_port, S_61_port, S_60_port, S_59_port, S_58_port, 
      S_57_port, S_56_port, S_55_port, S_54_port, S_53_port, S_52_port, 
      S_51_port, S_50_port, S_49_port, S_48_port, S_47_port, S_46_port, 
      S_45_port, S_44_port, S_43_port, S_42_port, S_41_port, S_40_port, 
      S_39_port, S_38_port, S_37_port, S_36_port, S_35_port, S_34_port, 
      S_33_port, S_32_port, S_31_port, S_30_port, S_29_port, S_28_port, 
      S_27_port, S_26_port, S_25_port, S_24_port, S_23_port, S_22_port, 
      S_21_port, S_20_port, S_19_port, S_18_port, S_17_port, S_16_port, 
      S_15_port, S_14_port, S_13_port, S_12_port, S_11_port, S_10_port, 
      S_9_port, S_8_port, S_7_port, S_6_port, S_5_port, S_4_port, S_3_port, 
      S_2_port, S_1_port, S_0_port, xor_b_63_port, xor_b_62_port, xor_b_61_port
      , xor_b_60_port, xor_b_59_port, xor_b_58_port, xor_b_57_port, 
      xor_b_56_port, xor_b_55_port, xor_b_54_port, xor_b_53_port, xor_b_52_port
      , xor_b_51_port, xor_b_50_port, xor_b_49_port, xor_b_48_port, 
      xor_b_47_port, xor_b_46_port, xor_b_45_port, xor_b_44_port, xor_b_43_port
      , xor_b_42_port, xor_b_41_port, xor_b_40_port, xor_b_39_port, 
      xor_b_38_port, xor_b_37_port, xor_b_36_port, xor_b_35_port, xor_b_34_port
      , xor_b_33_port, xor_b_32_port, xor_b_31_port, xor_b_30_port, 
      xor_b_29_port, xor_b_28_port, xor_b_27_port, xor_b_26_port, xor_b_25_port
      , xor_b_24_port, xor_b_23_port, xor_b_22_port, xor_b_21_port, 
      xor_b_20_port, xor_b_19_port, xor_b_18_port, xor_b_17_port, xor_b_16_port
      , xor_b_15_port, xor_b_14_port, xor_b_13_port, xor_b_12_port, 
      xor_b_11_port, xor_b_10_port, xor_b_9_port, xor_b_8_port, xor_b_7_port, 
      xor_b_6_port, xor_b_5_port, xor_b_4_port, xor_b_3_port, xor_b_2_port, 
      xor_b_1_port, xor_b_0_port, carry_14_port, carry_13_port, carry_12_port, 
      carry_11_port, carry_10_port, carry_9_port, carry_8_port, carry_7_port, 
      carry_6_port, carry_5_port, carry_4_port, carry_3_port, carry_2_port, 
      carry_1_port, carry_0_port, n3, n4 : std_logic;

begin
   S <= ( S_63_port, S_62_port, S_61_port, S_60_port, S_59_port, S_58_port, 
      S_57_port, S_56_port, S_55_port, S_54_port, S_53_port, S_52_port, 
      S_51_port, S_50_port, S_49_port, S_48_port, S_47_port, S_46_port, 
      S_45_port, S_44_port, S_43_port, S_42_port, S_41_port, S_40_port, 
      S_39_port, S_38_port, S_37_port, S_36_port, S_35_port, S_34_port, 
      S_33_port, S_32_port, S_31_port, S_30_port, S_29_port, S_28_port, 
      S_27_port, S_26_port, S_25_port, S_24_port, S_23_port, S_22_port, 
      S_21_port, S_20_port, S_19_port, S_18_port, S_17_port, S_16_port, 
      S_15_port, S_14_port, S_13_port, S_12_port, S_11_port, S_10_port, 
      S_9_port, S_8_port, S_7_port, S_6_port, S_5_port, S_4_port, S_3_port, 
      S_2_port, S_1_port, S_0_port );
   
   U3 : XOR2_X1 port map( A => xor_b_63_port, B => A(63), Z => n3);
   bc_xor_63 : my_xor_64 port map( A => B(63), B => Cin, xor_out => 
                           xor_b_63_port);
   bc_xor_62 : my_xor_63 port map( A => B(62), B => Cin, xor_out => 
                           xor_b_62_port);
   bc_xor_61 : my_xor_62 port map( A => B(61), B => Cin, xor_out => 
                           xor_b_61_port);
   bc_xor_60 : my_xor_61 port map( A => B(60), B => Cin, xor_out => 
                           xor_b_60_port);
   bc_xor_59 : my_xor_60 port map( A => B(59), B => Cin, xor_out => 
                           xor_b_59_port);
   bc_xor_58 : my_xor_59 port map( A => B(58), B => Cin, xor_out => 
                           xor_b_58_port);
   bc_xor_57 : my_xor_58 port map( A => B(57), B => Cin, xor_out => 
                           xor_b_57_port);
   bc_xor_56 : my_xor_57 port map( A => B(56), B => Cin, xor_out => 
                           xor_b_56_port);
   bc_xor_55 : my_xor_56 port map( A => B(55), B => Cin, xor_out => 
                           xor_b_55_port);
   bc_xor_54 : my_xor_55 port map( A => B(54), B => Cin, xor_out => 
                           xor_b_54_port);
   bc_xor_53 : my_xor_54 port map( A => B(53), B => Cin, xor_out => 
                           xor_b_53_port);
   bc_xor_52 : my_xor_53 port map( A => B(52), B => Cin, xor_out => 
                           xor_b_52_port);
   bc_xor_51 : my_xor_52 port map( A => B(51), B => Cin, xor_out => 
                           xor_b_51_port);
   bc_xor_50 : my_xor_51 port map( A => B(50), B => Cin, xor_out => 
                           xor_b_50_port);
   bc_xor_49 : my_xor_50 port map( A => B(49), B => Cin, xor_out => 
                           xor_b_49_port);
   bc_xor_48 : my_xor_49 port map( A => B(48), B => Cin, xor_out => 
                           xor_b_48_port);
   bc_xor_47 : my_xor_48 port map( A => B(47), B => Cin, xor_out => 
                           xor_b_47_port);
   bc_xor_46 : my_xor_47 port map( A => B(46), B => Cin, xor_out => 
                           xor_b_46_port);
   bc_xor_45 : my_xor_46 port map( A => B(45), B => Cin, xor_out => 
                           xor_b_45_port);
   bc_xor_44 : my_xor_45 port map( A => B(44), B => Cin, xor_out => 
                           xor_b_44_port);
   bc_xor_43 : my_xor_44 port map( A => B(43), B => Cin, xor_out => 
                           xor_b_43_port);
   bc_xor_42 : my_xor_43 port map( A => B(42), B => Cin, xor_out => 
                           xor_b_42_port);
   bc_xor_41 : my_xor_42 port map( A => B(41), B => Cin, xor_out => 
                           xor_b_41_port);
   bc_xor_40 : my_xor_41 port map( A => B(40), B => Cin, xor_out => 
                           xor_b_40_port);
   bc_xor_39 : my_xor_40 port map( A => B(39), B => Cin, xor_out => 
                           xor_b_39_port);
   bc_xor_38 : my_xor_39 port map( A => B(38), B => Cin, xor_out => 
                           xor_b_38_port);
   bc_xor_37 : my_xor_38 port map( A => B(37), B => Cin, xor_out => 
                           xor_b_37_port);
   bc_xor_36 : my_xor_37 port map( A => B(36), B => Cin, xor_out => 
                           xor_b_36_port);
   bc_xor_35 : my_xor_36 port map( A => B(35), B => Cin, xor_out => 
                           xor_b_35_port);
   bc_xor_34 : my_xor_35 port map( A => B(34), B => Cin, xor_out => 
                           xor_b_34_port);
   bc_xor_33 : my_xor_34 port map( A => B(33), B => Cin, xor_out => 
                           xor_b_33_port);
   bc_xor_32 : my_xor_33 port map( A => B(32), B => Cin, xor_out => 
                           xor_b_32_port);
   bc_xor_31 : my_xor_32 port map( A => B(31), B => Cin, xor_out => 
                           xor_b_31_port);
   bc_xor_30 : my_xor_31 port map( A => B(30), B => Cin, xor_out => 
                           xor_b_30_port);
   bc_xor_29 : my_xor_30 port map( A => B(29), B => Cin, xor_out => 
                           xor_b_29_port);
   bc_xor_28 : my_xor_29 port map( A => B(28), B => Cin, xor_out => 
                           xor_b_28_port);
   bc_xor_27 : my_xor_28 port map( A => B(27), B => Cin, xor_out => 
                           xor_b_27_port);
   bc_xor_26 : my_xor_27 port map( A => B(26), B => Cin, xor_out => 
                           xor_b_26_port);
   bc_xor_25 : my_xor_26 port map( A => B(25), B => Cin, xor_out => 
                           xor_b_25_port);
   bc_xor_24 : my_xor_25 port map( A => B(24), B => Cin, xor_out => 
                           xor_b_24_port);
   bc_xor_23 : my_xor_24 port map( A => B(23), B => Cin, xor_out => 
                           xor_b_23_port);
   bc_xor_22 : my_xor_23 port map( A => B(22), B => Cin, xor_out => 
                           xor_b_22_port);
   bc_xor_21 : my_xor_22 port map( A => B(21), B => Cin, xor_out => 
                           xor_b_21_port);
   bc_xor_20 : my_xor_21 port map( A => B(20), B => Cin, xor_out => 
                           xor_b_20_port);
   bc_xor_19 : my_xor_20 port map( A => B(19), B => Cin, xor_out => 
                           xor_b_19_port);
   bc_xor_18 : my_xor_19 port map( A => B(18), B => Cin, xor_out => 
                           xor_b_18_port);
   bc_xor_17 : my_xor_18 port map( A => B(17), B => Cin, xor_out => 
                           xor_b_17_port);
   bc_xor_16 : my_xor_17 port map( A => B(16), B => Cin, xor_out => 
                           xor_b_16_port);
   bc_xor_15 : my_xor_16 port map( A => B(15), B => Cin, xor_out => 
                           xor_b_15_port);
   bc_xor_14 : my_xor_15 port map( A => B(14), B => Cin, xor_out => 
                           xor_b_14_port);
   bc_xor_13 : my_xor_14 port map( A => B(13), B => Cin, xor_out => 
                           xor_b_13_port);
   bc_xor_12 : my_xor_13 port map( A => B(12), B => Cin, xor_out => 
                           xor_b_12_port);
   bc_xor_11 : my_xor_12 port map( A => B(11), B => Cin, xor_out => 
                           xor_b_11_port);
   bc_xor_10 : my_xor_11 port map( A => B(10), B => Cin, xor_out => 
                           xor_b_10_port);
   bc_xor_9 : my_xor_10 port map( A => B(9), B => Cin, xor_out => xor_b_9_port)
                           ;
   bc_xor_8 : my_xor_9 port map( A => B(8), B => Cin, xor_out => xor_b_8_port);
   bc_xor_7 : my_xor_8 port map( A => B(7), B => Cin, xor_out => xor_b_7_port);
   bc_xor_6 : my_xor_7 port map( A => B(6), B => Cin, xor_out => xor_b_6_port);
   bc_xor_5 : my_xor_6 port map( A => B(5), B => Cin, xor_out => xor_b_5_port);
   bc_xor_4 : my_xor_5 port map( A => B(4), B => Cin, xor_out => xor_b_4_port);
   bc_xor_3 : my_xor_4 port map( A => B(3), B => Cin, xor_out => xor_b_3_port);
   bc_xor_2 : my_xor_3 port map( A => B(2), B => Cin, xor_out => xor_b_2_port);
   bc_xor_1 : my_xor_2 port map( A => B(1), B => Cin, xor_out => xor_b_1_port);
   bc_xor_0 : my_xor_1 port map( A => B(0), B => Cin, xor_out => xor_b_0_port);
   CG : CARRY_GENERATOR_NBIT64_NBIT_PER_BLOCK4_1 port map( A(63) => A(63), 
                           A(62) => A(62), A(61) => A(61), A(60) => A(60), 
                           A(59) => A(59), A(58) => A(58), A(57) => A(57), 
                           A(56) => A(56), A(55) => A(55), A(54) => A(54), 
                           A(53) => A(53), A(52) => A(52), A(51) => A(51), 
                           A(50) => A(50), A(49) => A(49), A(48) => A(48), 
                           A(47) => A(47), A(46) => A(46), A(45) => A(45), 
                           A(44) => A(44), A(43) => A(43), A(42) => A(42), 
                           A(41) => A(41), A(40) => A(40), A(39) => A(39), 
                           A(38) => A(38), A(37) => A(37), A(36) => A(36), 
                           A(35) => A(35), A(34) => A(34), A(33) => A(33), 
                           A(32) => A(32), A(31) => A(31), A(30) => A(30), 
                           A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(63) => xor_b_63_port, B(62) =>
                           xor_b_62_port, B(61) => xor_b_61_port, B(60) => 
                           xor_b_60_port, B(59) => xor_b_59_port, B(58) => 
                           xor_b_58_port, B(57) => xor_b_57_port, B(56) => 
                           xor_b_56_port, B(55) => xor_b_55_port, B(54) => 
                           xor_b_54_port, B(53) => xor_b_53_port, B(52) => 
                           xor_b_52_port, B(51) => xor_b_51_port, B(50) => 
                           xor_b_50_port, B(49) => xor_b_49_port, B(48) => 
                           xor_b_48_port, B(47) => xor_b_47_port, B(46) => 
                           xor_b_46_port, B(45) => xor_b_45_port, B(44) => 
                           xor_b_44_port, B(43) => xor_b_43_port, B(42) => 
                           xor_b_42_port, B(41) => xor_b_41_port, B(40) => 
                           xor_b_40_port, B(39) => xor_b_39_port, B(38) => 
                           xor_b_38_port, B(37) => xor_b_37_port, B(36) => 
                           xor_b_36_port, B(35) => xor_b_35_port, B(34) => 
                           xor_b_34_port, B(33) => xor_b_33_port, B(32) => 
                           xor_b_32_port, B(31) => xor_b_31_port, B(30) => 
                           xor_b_30_port, B(29) => xor_b_29_port, B(28) => 
                           xor_b_28_port, B(27) => xor_b_27_port, B(26) => 
                           xor_b_26_port, B(25) => xor_b_25_port, B(24) => 
                           xor_b_24_port, B(23) => xor_b_23_port, B(22) => 
                           xor_b_22_port, B(21) => xor_b_21_port, B(20) => 
                           xor_b_20_port, B(19) => xor_b_19_port, B(18) => 
                           xor_b_18_port, B(17) => xor_b_17_port, B(16) => 
                           xor_b_16_port, B(15) => xor_b_15_port, B(14) => 
                           xor_b_14_port, B(13) => xor_b_13_port, B(12) => 
                           xor_b_12_port, B(11) => xor_b_11_port, B(10) => 
                           xor_b_10_port, B(9) => xor_b_9_port, B(8) => 
                           xor_b_8_port, B(7) => xor_b_7_port, B(6) => 
                           xor_b_6_port, B(5) => xor_b_5_port, B(4) => 
                           xor_b_4_port, B(3) => xor_b_3_port, B(2) => 
                           xor_b_2_port, B(1) => xor_b_1_port, B(0) => 
                           xor_b_0_port, Cin => Cin, Co(15) => Cout, Co(14) => 
                           carry_14_port, Co(13) => carry_13_port, Co(12) => 
                           carry_12_port, Co(11) => carry_11_port, Co(10) => 
                           carry_10_port, Co(9) => carry_9_port, Co(8) => 
                           carry_8_port, Co(7) => carry_7_port, Co(6) => 
                           carry_6_port, Co(5) => carry_5_port, Co(4) => 
                           carry_4_port, Co(3) => carry_3_port, Co(2) => 
                           carry_2_port, Co(1) => carry_1_port, Co(0) => 
                           carry_0_port);
   SG : sum_generator_n_bit64_n_CSB16_1 port map( A(63) => A(63), A(62) => 
                           A(62), A(61) => A(61), A(60) => A(60), A(59) => 
                           A(59), A(58) => A(58), A(57) => A(57), A(56) => 
                           A(56), A(55) => A(55), A(54) => A(54), A(53) => 
                           A(53), A(52) => A(52), A(51) => A(51), A(50) => 
                           A(50), A(49) => A(49), A(48) => A(48), A(47) => 
                           A(47), A(46) => A(46), A(45) => A(45), A(44) => 
                           A(44), A(43) => A(43), A(42) => A(42), A(41) => 
                           A(41), A(40) => A(40), A(39) => A(39), A(38) => 
                           A(38), A(37) => A(37), A(36) => A(36), A(35) => 
                           A(35), A(34) => A(34), A(33) => A(33), A(32) => 
                           A(32), A(31) => A(31), A(30) => A(30), A(29) => 
                           A(29), A(28) => A(28), A(27) => A(27), A(26) => 
                           A(26), A(25) => A(25), A(24) => A(24), A(23) => 
                           A(23), A(22) => A(22), A(21) => A(21), A(20) => 
                           A(20), A(19) => A(19), A(18) => A(18), A(17) => 
                           A(17), A(16) => A(16), A(15) => A(15), A(14) => 
                           A(14), A(13) => A(13), A(12) => A(12), A(11) => 
                           A(11), A(10) => A(10), A(9) => A(9), A(8) => A(8), 
                           A(7) => A(7), A(6) => A(6), A(5) => A(5), A(4) => 
                           A(4), A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(63) => xor_b_63_port, B(62) => 
                           xor_b_62_port, B(61) => xor_b_61_port, B(60) => 
                           xor_b_60_port, B(59) => xor_b_59_port, B(58) => 
                           xor_b_58_port, B(57) => xor_b_57_port, B(56) => 
                           xor_b_56_port, B(55) => xor_b_55_port, B(54) => 
                           xor_b_54_port, B(53) => xor_b_53_port, B(52) => 
                           xor_b_52_port, B(51) => xor_b_51_port, B(50) => 
                           xor_b_50_port, B(49) => xor_b_49_port, B(48) => 
                           xor_b_48_port, B(47) => xor_b_47_port, B(46) => 
                           xor_b_46_port, B(45) => xor_b_45_port, B(44) => 
                           xor_b_44_port, B(43) => xor_b_43_port, B(42) => 
                           xor_b_42_port, B(41) => xor_b_41_port, B(40) => 
                           xor_b_40_port, B(39) => xor_b_39_port, B(38) => 
                           xor_b_38_port, B(37) => xor_b_37_port, B(36) => 
                           xor_b_36_port, B(35) => xor_b_35_port, B(34) => 
                           xor_b_34_port, B(33) => xor_b_33_port, B(32) => 
                           xor_b_32_port, B(31) => xor_b_31_port, B(30) => 
                           xor_b_30_port, B(29) => xor_b_29_port, B(28) => 
                           xor_b_28_port, B(27) => xor_b_27_port, B(26) => 
                           xor_b_26_port, B(25) => xor_b_25_port, B(24) => 
                           xor_b_24_port, B(23) => xor_b_23_port, B(22) => 
                           xor_b_22_port, B(21) => xor_b_21_port, B(20) => 
                           xor_b_20_port, B(19) => xor_b_19_port, B(18) => 
                           xor_b_18_port, B(17) => xor_b_17_port, B(16) => 
                           xor_b_16_port, B(15) => xor_b_15_port, B(14) => 
                           xor_b_14_port, B(13) => xor_b_13_port, B(12) => 
                           xor_b_12_port, B(11) => xor_b_11_port, B(10) => 
                           xor_b_10_port, B(9) => xor_b_9_port, B(8) => 
                           xor_b_8_port, B(7) => xor_b_7_port, B(6) => 
                           xor_b_6_port, B(5) => xor_b_5_port, B(4) => 
                           xor_b_4_port, B(3) => xor_b_3_port, B(2) => 
                           xor_b_2_port, B(1) => xor_b_1_port, B(0) => 
                           xor_b_0_port, C_in(15) => carry_14_port, C_in(14) =>
                           carry_13_port, C_in(13) => carry_12_port, C_in(12) 
                           => carry_11_port, C_in(11) => carry_10_port, 
                           C_in(10) => carry_9_port, C_in(9) => carry_8_port, 
                           C_in(8) => carry_7_port, C_in(7) => carry_6_port, 
                           C_in(6) => carry_5_port, C_in(5) => carry_4_port, 
                           C_in(4) => carry_3_port, C_in(3) => carry_2_port, 
                           C_in(2) => carry_1_port, C_in(1) => carry_0_port, 
                           C_in(0) => Cin, S(63) => S_63_port, S(62) => 
                           S_62_port, S(61) => S_61_port, S(60) => S_60_port, 
                           S(59) => S_59_port, S(58) => S_58_port, S(57) => 
                           S_57_port, S(56) => S_56_port, S(55) => S_55_port, 
                           S(54) => S_54_port, S(53) => S_53_port, S(52) => 
                           S_52_port, S(51) => S_51_port, S(50) => S_50_port, 
                           S(49) => S_49_port, S(48) => S_48_port, S(47) => 
                           S_47_port, S(46) => S_46_port, S(45) => S_45_port, 
                           S(44) => S_44_port, S(43) => S_43_port, S(42) => 
                           S_42_port, S(41) => S_41_port, S(40) => S_40_port, 
                           S(39) => S_39_port, S(38) => S_38_port, S(37) => 
                           S_37_port, S(36) => S_36_port, S(35) => S_35_port, 
                           S(34) => S_34_port, S(33) => S_33_port, S(32) => 
                           S_32_port, S(31) => S_31_port, S(30) => S_30_port, 
                           S(29) => S_29_port, S(28) => S_28_port, S(27) => 
                           S_27_port, S(26) => S_26_port, S(25) => S_25_port, 
                           S(24) => S_24_port, S(23) => S_23_port, S(22) => 
                           S_22_port, S(21) => S_21_port, S(20) => S_20_port, 
                           S(19) => S_19_port, S(18) => S_18_port, S(17) => 
                           S_17_port, S(16) => S_16_port, S(15) => S_15_port, 
                           S(14) => S_14_port, S(13) => S_13_port, S(12) => 
                           S_12_port, S(11) => S_11_port, S(10) => S_10_port, 
                           S(9) => S_9_port, S(8) => S_8_port, S(7) => S_7_port
                           , S(6) => S_6_port, S(5) => S_5_port, S(4) => 
                           S_4_port, S(3) => S_3_port, S(2) => S_2_port, S(1) 
                           => S_1_port, S(0) => S_0_port);
   U1 : NOR2_X1 port map( A1 => n4, A2 => n3, ZN => ovf);
   U2 : XNOR2_X1 port map( A => A(63), B => S_63_port, ZN => n4);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity mux51_gen_NBIT32_3 is

   port( A0, A1, A2, A3, A4 : in std_logic_vector (31 downto 0);  SEL : in 
         std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end mux51_gen_NBIT32_3;

architecture SYN_data_fl of mux51_gen_NBIT32_3 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, 
      n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98
      , n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, 
      n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, 
      n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, 
      n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, 
      n147, n148, n149, n150, n151, n152, n153, n154, n155 : std_logic;

begin
   
   U2 : BUF_X1 port map( A => n150, Z => n73);
   U3 : BUF_X1 port map( A => n150, Z => n74);
   U4 : BUF_X1 port map( A => n149, Z => n1);
   U5 : BUF_X1 port map( A => n153, Z => n82);
   U6 : BUF_X1 port map( A => n153, Z => n83);
   U7 : BUF_X1 port map( A => n153, Z => n84);
   U8 : BUF_X1 port map( A => n152, Z => n79);
   U9 : BUF_X1 port map( A => n152, Z => n80);
   U10 : BUF_X1 port map( A => n151, Z => n76);
   U11 : BUF_X1 port map( A => n151, Z => n77);
   U12 : BUF_X1 port map( A => n150, Z => n75);
   U13 : BUF_X1 port map( A => n152, Z => n81);
   U14 : BUF_X1 port map( A => n151, Z => n78);
   U15 : INV_X1 port map( A => SEL(2), ZN => n86);
   U16 : INV_X1 port map( A => SEL(1), ZN => n85);
   U17 : BUF_X1 port map( A => n149, Z => n2);
   U18 : BUF_X1 port map( A => n149, Z => n72);
   U19 : NOR3_X1 port map( A1 => SEL(0), A2 => SEL(2), A3 => n85, ZN => n153);
   U20 : NOR3_X1 port map( A1 => SEL(0), A2 => SEL(1), A3 => n1, ZN => n150);
   U21 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => SEL(0), ZN => n149
                           );
   U22 : AND3_X1 port map( A1 => SEL(0), A2 => n86, A3 => SEL(1), ZN => n151);
   U23 : AND3_X1 port map( A1 => n85, A2 => n86, A3 => SEL(0), ZN => n152);
   U24 : NAND2_X1 port map( A1 => n126, A2 => n125, ZN => Y(27));
   U25 : AOI22_X1 port map( A1 => A4(27), A2 => n74, B1 => A0(27), B2 => n2, ZN
                           => n126);
   U26 : AOI222_X1 port map( A1 => A2(27), A2 => n83, B1 => A1(27), B2 => n80, 
                           C1 => A3(27), C2 => n77, ZN => n125);
   U27 : NAND2_X1 port map( A1 => n128, A2 => n127, ZN => Y(28));
   U28 : AOI22_X1 port map( A1 => A4(28), A2 => n74, B1 => A0(28), B2 => n2, ZN
                           => n128);
   U29 : AOI222_X1 port map( A1 => A2(28), A2 => n83, B1 => A1(28), B2 => n80, 
                           C1 => A3(28), C2 => n77, ZN => n127);
   U30 : NAND2_X1 port map( A1 => n130, A2 => n129, ZN => Y(29));
   U31 : AOI22_X1 port map( A1 => A4(29), A2 => n74, B1 => A0(29), B2 => n2, ZN
                           => n130);
   U32 : AOI222_X1 port map( A1 => A2(29), A2 => n83, B1 => A1(29), B2 => n80, 
                           C1 => A3(29), C2 => n77, ZN => n129);
   U33 : NAND2_X1 port map( A1 => n134, A2 => n133, ZN => Y(30));
   U34 : AOI22_X1 port map( A1 => A4(30), A2 => n74, B1 => A0(30), B2 => n72, 
                           ZN => n134);
   U35 : AOI222_X1 port map( A1 => A2(30), A2 => n84, B1 => A1(30), B2 => n80, 
                           C1 => A3(30), C2 => n77, ZN => n133);
   U36 : NAND2_X1 port map( A1 => n136, A2 => n135, ZN => Y(31));
   U37 : AOI22_X1 port map( A1 => A4(31), A2 => n75, B1 => A0(31), B2 => n72, 
                           ZN => n136);
   U38 : AOI222_X1 port map( A1 => A2(31), A2 => n84, B1 => A1(31), B2 => n81, 
                           C1 => A3(31), C2 => n78, ZN => n135);
   U39 : NAND2_X1 port map( A1 => n120, A2 => n119, ZN => Y(24));
   U40 : AOI22_X1 port map( A1 => A4(24), A2 => n74, B1 => A0(24), B2 => n2, ZN
                           => n120);
   U41 : AOI222_X1 port map( A1 => A2(24), A2 => n83, B1 => A1(24), B2 => n80, 
                           C1 => A3(24), C2 => n77, ZN => n119);
   U42 : NAND2_X1 port map( A1 => n122, A2 => n121, ZN => Y(25));
   U43 : AOI22_X1 port map( A1 => A4(25), A2 => n74, B1 => A0(25), B2 => n2, ZN
                           => n122);
   U44 : AOI222_X1 port map( A1 => A2(25), A2 => n83, B1 => A1(25), B2 => n80, 
                           C1 => A3(25), C2 => n77, ZN => n121);
   U45 : NAND2_X1 port map( A1 => n124, A2 => n123, ZN => Y(26));
   U46 : AOI22_X1 port map( A1 => A4(26), A2 => n74, B1 => A0(26), B2 => n2, ZN
                           => n124);
   U47 : AOI222_X1 port map( A1 => A2(26), A2 => n83, B1 => A1(26), B2 => n80, 
                           C1 => A3(26), C2 => n77, ZN => n123);
   U48 : NAND2_X1 port map( A1 => n96, A2 => n95, ZN => Y(13));
   U49 : AOI22_X1 port map( A1 => A4(13), A2 => n73, B1 => A0(13), B2 => n1, ZN
                           => n96);
   U50 : AOI222_X1 port map( A1 => A2(13), A2 => n82, B1 => A1(13), B2 => n79, 
                           C1 => A3(13), C2 => n76, ZN => n95);
   U51 : NAND2_X1 port map( A1 => n98, A2 => n97, ZN => Y(14));
   U52 : AOI22_X1 port map( A1 => A4(14), A2 => n73, B1 => A0(14), B2 => n1, ZN
                           => n98);
   U53 : AOI222_X1 port map( A1 => A2(14), A2 => n82, B1 => A1(14), B2 => n79, 
                           C1 => A3(14), C2 => n76, ZN => n97);
   U54 : NAND2_X1 port map( A1 => n100, A2 => n99, ZN => Y(15));
   U55 : AOI22_X1 port map( A1 => A4(15), A2 => n73, B1 => A0(15), B2 => n1, ZN
                           => n100);
   U56 : AOI222_X1 port map( A1 => A2(15), A2 => n82, B1 => A1(15), B2 => n79, 
                           C1 => A3(15), C2 => n76, ZN => n99);
   U57 : NAND2_X1 port map( A1 => n102, A2 => n101, ZN => Y(16));
   U58 : AOI22_X1 port map( A1 => A4(16), A2 => n73, B1 => A0(16), B2 => n1, ZN
                           => n102);
   U59 : AOI222_X1 port map( A1 => A2(16), A2 => n82, B1 => A1(16), B2 => n79, 
                           C1 => A3(16), C2 => n76, ZN => n101);
   U60 : NAND2_X1 port map( A1 => n104, A2 => n103, ZN => Y(17));
   U61 : AOI22_X1 port map( A1 => A4(17), A2 => n73, B1 => A0(17), B2 => n1, ZN
                           => n104);
   U62 : AOI222_X1 port map( A1 => A2(17), A2 => n82, B1 => A1(17), B2 => n79, 
                           C1 => A3(17), C2 => n76, ZN => n103);
   U63 : NAND2_X1 port map( A1 => n106, A2 => n105, ZN => Y(18));
   U64 : AOI22_X1 port map( A1 => A4(18), A2 => n73, B1 => A0(18), B2 => n1, ZN
                           => n106);
   U65 : AOI222_X1 port map( A1 => A2(18), A2 => n82, B1 => A1(18), B2 => n79, 
                           C1 => A3(18), C2 => n76, ZN => n105);
   U66 : NAND2_X1 port map( A1 => n108, A2 => n107, ZN => Y(19));
   U67 : AOI22_X1 port map( A1 => A4(19), A2 => n73, B1 => A0(19), B2 => n1, ZN
                           => n108);
   U68 : AOI222_X1 port map( A1 => A2(19), A2 => n82, B1 => A1(19), B2 => n79, 
                           C1 => A3(19), C2 => n76, ZN => n107);
   U69 : NAND2_X1 port map( A1 => n112, A2 => n111, ZN => Y(20));
   U70 : AOI22_X1 port map( A1 => A4(20), A2 => n74, B1 => A0(20), B2 => n2, ZN
                           => n112);
   U71 : AOI222_X1 port map( A1 => A2(20), A2 => n83, B1 => A1(20), B2 => n80, 
                           C1 => A3(20), C2 => n77, ZN => n111);
   U72 : NAND2_X1 port map( A1 => n114, A2 => n113, ZN => Y(21));
   U73 : AOI22_X1 port map( A1 => A4(21), A2 => n74, B1 => A0(21), B2 => n2, ZN
                           => n114);
   U74 : AOI222_X1 port map( A1 => A2(21), A2 => n83, B1 => A1(21), B2 => n80, 
                           C1 => A3(21), C2 => n77, ZN => n113);
   U75 : NAND2_X1 port map( A1 => n116, A2 => n115, ZN => Y(22));
   U76 : AOI22_X1 port map( A1 => A4(22), A2 => n74, B1 => A0(22), B2 => n2, ZN
                           => n116);
   U77 : AOI222_X1 port map( A1 => A2(22), A2 => n83, B1 => A1(22), B2 => n80, 
                           C1 => A3(22), C2 => n77, ZN => n115);
   U78 : NAND2_X1 port map( A1 => n118, A2 => n117, ZN => Y(23));
   U79 : AOI22_X1 port map( A1 => A4(23), A2 => n74, B1 => A0(23), B2 => n2, ZN
                           => n118);
   U80 : AOI222_X1 port map( A1 => A2(23), A2 => n83, B1 => A1(23), B2 => n80, 
                           C1 => A3(23), C2 => n77, ZN => n117);
   U81 : NAND2_X1 port map( A1 => n90, A2 => n89, ZN => Y(10));
   U82 : AOI22_X1 port map( A1 => A4(10), A2 => n73, B1 => A0(10), B2 => n1, ZN
                           => n90);
   U83 : AOI222_X1 port map( A1 => A2(10), A2 => n82, B1 => A1(10), B2 => n79, 
                           C1 => A3(10), C2 => n76, ZN => n89);
   U84 : NAND2_X1 port map( A1 => n92, A2 => n91, ZN => Y(11));
   U85 : AOI22_X1 port map( A1 => A4(11), A2 => n73, B1 => A0(11), B2 => n1, ZN
                           => n92);
   U86 : AOI222_X1 port map( A1 => A2(11), A2 => n82, B1 => A1(11), B2 => n79, 
                           C1 => A3(11), C2 => n76, ZN => n91);
   U87 : NAND2_X1 port map( A1 => n94, A2 => n93, ZN => Y(12));
   U88 : AOI22_X1 port map( A1 => A4(12), A2 => n73, B1 => A0(12), B2 => n1, ZN
                           => n94);
   U89 : AOI222_X1 port map( A1 => A2(12), A2 => n82, B1 => A1(12), B2 => n79, 
                           C1 => A3(12), C2 => n76, ZN => n93);
   U90 : NAND2_X1 port map( A1 => n138, A2 => n137, ZN => Y(3));
   U91 : AOI222_X1 port map( A1 => A2(3), A2 => n84, B1 => A1(3), B2 => n81, C1
                           => A3(3), C2 => n78, ZN => n137);
   U92 : AOI22_X1 port map( A1 => A4(3), A2 => n75, B1 => A0(3), B2 => n72, ZN 
                           => n138);
   U93 : NAND2_X1 port map( A1 => n140, A2 => n139, ZN => Y(4));
   U94 : AOI222_X1 port map( A1 => A2(4), A2 => n84, B1 => A1(4), B2 => n81, C1
                           => A3(4), C2 => n78, ZN => n139);
   U95 : AOI22_X1 port map( A1 => A4(4), A2 => n75, B1 => A0(4), B2 => n72, ZN 
                           => n140);
   U96 : NAND2_X1 port map( A1 => n142, A2 => n141, ZN => Y(5));
   U97 : AOI222_X1 port map( A1 => A2(5), A2 => n84, B1 => A1(5), B2 => n81, C1
                           => A3(5), C2 => n78, ZN => n141);
   U98 : AOI22_X1 port map( A1 => A4(5), A2 => n75, B1 => A0(5), B2 => n72, ZN 
                           => n142);
   U99 : NAND2_X1 port map( A1 => n144, A2 => n143, ZN => Y(6));
   U100 : AOI22_X1 port map( A1 => A4(6), A2 => n75, B1 => A0(6), B2 => n72, ZN
                           => n144);
   U101 : AOI222_X1 port map( A1 => A2(6), A2 => n84, B1 => A1(6), B2 => n81, 
                           C1 => A3(6), C2 => n78, ZN => n143);
   U102 : NAND2_X1 port map( A1 => n146, A2 => n145, ZN => Y(7));
   U103 : AOI22_X1 port map( A1 => A4(7), A2 => n75, B1 => A0(7), B2 => n72, ZN
                           => n146);
   U104 : AOI222_X1 port map( A1 => A2(7), A2 => n84, B1 => A1(7), B2 => n81, 
                           C1 => A3(7), C2 => n78, ZN => n145);
   U105 : NAND2_X1 port map( A1 => n148, A2 => n147, ZN => Y(8));
   U106 : AOI22_X1 port map( A1 => A4(8), A2 => n75, B1 => A0(8), B2 => n72, ZN
                           => n148);
   U107 : AOI222_X1 port map( A1 => A2(8), A2 => n84, B1 => A1(8), B2 => n81, 
                           C1 => A3(8), C2 => n78, ZN => n147);
   U108 : NAND2_X1 port map( A1 => n155, A2 => n154, ZN => Y(9));
   U109 : AOI22_X1 port map( A1 => A4(9), A2 => n75, B1 => A0(9), B2 => n72, ZN
                           => n155);
   U110 : AOI222_X1 port map( A1 => A2(9), A2 => n84, B1 => A1(9), B2 => n81, 
                           C1 => A3(9), C2 => n78, ZN => n154);
   U111 : NAND2_X1 port map( A1 => n132, A2 => n131, ZN => Y(2));
   U112 : AOI22_X1 port map( A1 => A4(2), A2 => n74, B1 => A0(2), B2 => n2, ZN 
                           => n132);
   U113 : AOI222_X1 port map( A1 => A2(2), A2 => n84, B1 => A1(2), B2 => n80, 
                           C1 => A3(2), C2 => n77, ZN => n131);
   U114 : NAND2_X1 port map( A1 => n110, A2 => n109, ZN => Y(1));
   U115 : AOI22_X1 port map( A1 => A4(1), A2 => n73, B1 => A0(1), B2 => n2, ZN 
                           => n110);
   U116 : AOI222_X1 port map( A1 => A2(1), A2 => n83, B1 => A1(1), B2 => n79, 
                           C1 => A3(1), C2 => n76, ZN => n109);
   U117 : NAND2_X1 port map( A1 => n88, A2 => n87, ZN => Y(0));
   U118 : AOI22_X1 port map( A1 => A4(0), A2 => n73, B1 => A0(0), B2 => n1, ZN 
                           => n88);
   U119 : AOI222_X1 port map( A1 => A2(0), A2 => n82, B1 => A1(0), B2 => n79, 
                           C1 => A3(0), C2 => n76, ZN => n87);

end SYN_data_fl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity mux51_gen_NBIT32_2 is

   port( A0, A1, A2, A3, A4 : in std_logic_vector (31 downto 0);  SEL : in 
         std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end mux51_gen_NBIT32_2;

architecture SYN_data_fl of mux51_gen_NBIT32_2 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, 
      n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98
      , n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, 
      n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, 
      n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, 
      n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, 
      n147, n148, n149, n150, n151, n152, n153, n154, n155 : std_logic;

begin
   
   U2 : BUF_X1 port map( A => n150, Z => n74);
   U3 : BUF_X1 port map( A => n150, Z => n73);
   U4 : BUF_X1 port map( A => n149, Z => n1);
   U5 : BUF_X1 port map( A => n153, Z => n83);
   U6 : BUF_X1 port map( A => n153, Z => n82);
   U7 : BUF_X1 port map( A => n153, Z => n84);
   U8 : BUF_X1 port map( A => n152, Z => n80);
   U9 : BUF_X1 port map( A => n152, Z => n79);
   U10 : BUF_X1 port map( A => n151, Z => n77);
   U11 : BUF_X1 port map( A => n151, Z => n76);
   U12 : BUF_X1 port map( A => n150, Z => n75);
   U13 : BUF_X1 port map( A => n152, Z => n81);
   U14 : BUF_X1 port map( A => n151, Z => n78);
   U15 : BUF_X1 port map( A => n149, Z => n2);
   U16 : BUF_X1 port map( A => n149, Z => n72);
   U17 : NAND2_X1 port map( A1 => n134, A2 => n133, ZN => Y(30));
   U18 : AOI22_X1 port map( A1 => A4(30), A2 => n74, B1 => A0(30), B2 => n72, 
                           ZN => n134);
   U19 : AOI222_X1 port map( A1 => A2(30), A2 => n84, B1 => A1(30), B2 => n80, 
                           C1 => A3(30), C2 => n77, ZN => n133);
   U20 : NAND2_X1 port map( A1 => n130, A2 => n129, ZN => Y(29));
   U21 : AOI22_X1 port map( A1 => A4(29), A2 => n74, B1 => A0(29), B2 => n2, ZN
                           => n130);
   U22 : AOI222_X1 port map( A1 => A2(29), A2 => n83, B1 => A1(29), B2 => n80, 
                           C1 => A3(29), C2 => n77, ZN => n129);
   U23 : NAND2_X1 port map( A1 => n128, A2 => n127, ZN => Y(28));
   U24 : AOI22_X1 port map( A1 => A4(28), A2 => n74, B1 => A0(28), B2 => n2, ZN
                           => n128);
   U25 : AOI222_X1 port map( A1 => A2(28), A2 => n83, B1 => A1(28), B2 => n80, 
                           C1 => A3(28), C2 => n77, ZN => n127);
   U26 : NAND2_X1 port map( A1 => n126, A2 => n125, ZN => Y(27));
   U27 : AOI22_X1 port map( A1 => A4(27), A2 => n74, B1 => A0(27), B2 => n2, ZN
                           => n126);
   U28 : AOI222_X1 port map( A1 => A2(27), A2 => n83, B1 => A1(27), B2 => n80, 
                           C1 => A3(27), C2 => n77, ZN => n125);
   U29 : NAND2_X1 port map( A1 => n124, A2 => n123, ZN => Y(26));
   U30 : AOI22_X1 port map( A1 => A4(26), A2 => n74, B1 => A0(26), B2 => n2, ZN
                           => n124);
   U31 : AOI222_X1 port map( A1 => A2(26), A2 => n83, B1 => A1(26), B2 => n80, 
                           C1 => A3(26), C2 => n77, ZN => n123);
   U32 : NAND2_X1 port map( A1 => n122, A2 => n121, ZN => Y(25));
   U33 : AOI22_X1 port map( A1 => A4(25), A2 => n74, B1 => A0(25), B2 => n2, ZN
                           => n122);
   U34 : AOI222_X1 port map( A1 => A2(25), A2 => n83, B1 => A1(25), B2 => n80, 
                           C1 => A3(25), C2 => n77, ZN => n121);
   U35 : NAND2_X1 port map( A1 => n120, A2 => n119, ZN => Y(24));
   U36 : AOI22_X1 port map( A1 => A4(24), A2 => n74, B1 => A0(24), B2 => n2, ZN
                           => n120);
   U37 : AOI222_X1 port map( A1 => A2(24), A2 => n83, B1 => A1(24), B2 => n80, 
                           C1 => A3(24), C2 => n77, ZN => n119);
   U38 : NAND2_X1 port map( A1 => n118, A2 => n117, ZN => Y(23));
   U39 : AOI22_X1 port map( A1 => A4(23), A2 => n74, B1 => A0(23), B2 => n2, ZN
                           => n118);
   U40 : AOI222_X1 port map( A1 => A2(23), A2 => n83, B1 => A1(23), B2 => n80, 
                           C1 => A3(23), C2 => n77, ZN => n117);
   U41 : NAND2_X1 port map( A1 => n116, A2 => n115, ZN => Y(22));
   U42 : AOI22_X1 port map( A1 => A4(22), A2 => n74, B1 => A0(22), B2 => n2, ZN
                           => n116);
   U43 : AOI222_X1 port map( A1 => A2(22), A2 => n83, B1 => A1(22), B2 => n80, 
                           C1 => A3(22), C2 => n77, ZN => n115);
   U44 : NAND2_X1 port map( A1 => n136, A2 => n135, ZN => Y(31));
   U45 : AOI22_X1 port map( A1 => A4(31), A2 => n75, B1 => A0(31), B2 => n72, 
                           ZN => n136);
   U46 : AOI222_X1 port map( A1 => A2(31), A2 => n84, B1 => A1(31), B2 => n81, 
                           C1 => A3(31), C2 => n78, ZN => n135);
   U47 : NAND2_X1 port map( A1 => n114, A2 => n113, ZN => Y(21));
   U48 : AOI22_X1 port map( A1 => A4(21), A2 => n74, B1 => A0(21), B2 => n2, ZN
                           => n114);
   U49 : AOI222_X1 port map( A1 => A2(21), A2 => n83, B1 => A1(21), B2 => n80, 
                           C1 => A3(21), C2 => n77, ZN => n113);
   U50 : NAND2_X1 port map( A1 => n112, A2 => n111, ZN => Y(20));
   U51 : AOI22_X1 port map( A1 => A4(20), A2 => n74, B1 => A0(20), B2 => n2, ZN
                           => n112);
   U52 : AOI222_X1 port map( A1 => A2(20), A2 => n83, B1 => A1(20), B2 => n80, 
                           C1 => A3(20), C2 => n77, ZN => n111);
   U53 : NAND2_X1 port map( A1 => n108, A2 => n107, ZN => Y(19));
   U54 : AOI22_X1 port map( A1 => A4(19), A2 => n73, B1 => A0(19), B2 => n1, ZN
                           => n108);
   U55 : AOI222_X1 port map( A1 => A2(19), A2 => n82, B1 => A1(19), B2 => n79, 
                           C1 => A3(19), C2 => n76, ZN => n107);
   U56 : NAND2_X1 port map( A1 => n106, A2 => n105, ZN => Y(18));
   U57 : AOI22_X1 port map( A1 => A4(18), A2 => n73, B1 => A0(18), B2 => n1, ZN
                           => n106);
   U58 : AOI222_X1 port map( A1 => A2(18), A2 => n82, B1 => A1(18), B2 => n79, 
                           C1 => A3(18), C2 => n76, ZN => n105);
   U59 : NAND2_X1 port map( A1 => n104, A2 => n103, ZN => Y(17));
   U60 : AOI22_X1 port map( A1 => A4(17), A2 => n73, B1 => A0(17), B2 => n1, ZN
                           => n104);
   U61 : AOI222_X1 port map( A1 => A2(17), A2 => n82, B1 => A1(17), B2 => n79, 
                           C1 => A3(17), C2 => n76, ZN => n103);
   U62 : NAND2_X1 port map( A1 => n102, A2 => n101, ZN => Y(16));
   U63 : AOI22_X1 port map( A1 => A4(16), A2 => n73, B1 => A0(16), B2 => n1, ZN
                           => n102);
   U64 : AOI222_X1 port map( A1 => A2(16), A2 => n82, B1 => A1(16), B2 => n79, 
                           C1 => A3(16), C2 => n76, ZN => n101);
   U65 : NAND2_X1 port map( A1 => n100, A2 => n99, ZN => Y(15));
   U66 : AOI22_X1 port map( A1 => A4(15), A2 => n73, B1 => A0(15), B2 => n1, ZN
                           => n100);
   U67 : AOI222_X1 port map( A1 => A2(15), A2 => n82, B1 => A1(15), B2 => n79, 
                           C1 => A3(15), C2 => n76, ZN => n99);
   U68 : NAND2_X1 port map( A1 => n98, A2 => n97, ZN => Y(14));
   U69 : AOI22_X1 port map( A1 => A4(14), A2 => n73, B1 => A0(14), B2 => n1, ZN
                           => n98);
   U70 : AOI222_X1 port map( A1 => A2(14), A2 => n82, B1 => A1(14), B2 => n79, 
                           C1 => A3(14), C2 => n76, ZN => n97);
   U71 : NAND2_X1 port map( A1 => n96, A2 => n95, ZN => Y(13));
   U72 : AOI22_X1 port map( A1 => A4(13), A2 => n73, B1 => A0(13), B2 => n1, ZN
                           => n96);
   U73 : AOI222_X1 port map( A1 => A2(13), A2 => n82, B1 => A1(13), B2 => n79, 
                           C1 => A3(13), C2 => n76, ZN => n95);
   U74 : NAND2_X1 port map( A1 => n94, A2 => n93, ZN => Y(12));
   U75 : AOI22_X1 port map( A1 => A4(12), A2 => n73, B1 => A0(12), B2 => n1, ZN
                           => n94);
   U76 : AOI222_X1 port map( A1 => A2(12), A2 => n82, B1 => A1(12), B2 => n79, 
                           C1 => A3(12), C2 => n76, ZN => n93);
   U77 : NAND2_X1 port map( A1 => n92, A2 => n91, ZN => Y(11));
   U78 : AOI22_X1 port map( A1 => A4(11), A2 => n73, B1 => A0(11), B2 => n1, ZN
                           => n92);
   U79 : AOI222_X1 port map( A1 => A2(11), A2 => n82, B1 => A1(11), B2 => n79, 
                           C1 => A3(11), C2 => n76, ZN => n91);
   U80 : NAND2_X1 port map( A1 => n155, A2 => n154, ZN => Y(9));
   U81 : AOI22_X1 port map( A1 => A4(9), A2 => n75, B1 => A0(9), B2 => n72, ZN 
                           => n155);
   U82 : AOI222_X1 port map( A1 => A2(9), A2 => n84, B1 => A1(9), B2 => n81, C1
                           => A3(9), C2 => n78, ZN => n154);
   U83 : NAND2_X1 port map( A1 => n148, A2 => n147, ZN => Y(8));
   U84 : AOI22_X1 port map( A1 => A4(8), A2 => n75, B1 => A0(8), B2 => n72, ZN 
                           => n148);
   U85 : AOI222_X1 port map( A1 => A2(8), A2 => n84, B1 => A1(8), B2 => n81, C1
                           => A3(8), C2 => n78, ZN => n147);
   U86 : NAND2_X1 port map( A1 => n90, A2 => n89, ZN => Y(10));
   U87 : AOI22_X1 port map( A1 => A4(10), A2 => n73, B1 => A0(10), B2 => n1, ZN
                           => n90);
   U88 : AOI222_X1 port map( A1 => A2(10), A2 => n82, B1 => A1(10), B2 => n79, 
                           C1 => A3(10), C2 => n76, ZN => n89);
   U89 : NAND2_X1 port map( A1 => n140, A2 => n139, ZN => Y(4));
   U90 : AOI22_X1 port map( A1 => A4(4), A2 => n75, B1 => A0(4), B2 => n72, ZN 
                           => n140);
   U91 : AOI222_X1 port map( A1 => A2(4), A2 => n84, B1 => A1(4), B2 => n81, C1
                           => A3(4), C2 => n78, ZN => n139);
   U92 : NOR3_X1 port map( A1 => SEL(0), A2 => SEL(1), A3 => n1, ZN => n150);
   U93 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => SEL(0), ZN => n149
                           );
   U94 : NOR3_X1 port map( A1 => SEL(0), A2 => SEL(2), A3 => n86, ZN => n153);
   U95 : NAND2_X1 port map( A1 => n144, A2 => n143, ZN => Y(6));
   U96 : AOI222_X1 port map( A1 => A2(6), A2 => n84, B1 => A1(6), B2 => n81, C1
                           => A3(6), C2 => n78, ZN => n143);
   U97 : AOI22_X1 port map( A1 => A4(6), A2 => n75, B1 => A0(6), B2 => n72, ZN 
                           => n144);
   U98 : NAND2_X1 port map( A1 => n142, A2 => n141, ZN => Y(5));
   U99 : AOI222_X1 port map( A1 => A2(5), A2 => n84, B1 => A1(5), B2 => n81, C1
                           => A3(5), C2 => n78, ZN => n141);
   U100 : AOI22_X1 port map( A1 => A4(5), A2 => n75, B1 => A0(5), B2 => n72, ZN
                           => n142);
   U101 : AND3_X1 port map( A1 => SEL(0), A2 => n85, A3 => SEL(1), ZN => n151);
   U102 : AND3_X1 port map( A1 => n86, A2 => n85, A3 => SEL(0), ZN => n152);
   U103 : INV_X1 port map( A => SEL(1), ZN => n86);
   U104 : NAND2_X1 port map( A1 => n146, A2 => n145, ZN => Y(7));
   U105 : AOI22_X1 port map( A1 => A4(7), A2 => n75, B1 => A0(7), B2 => n72, ZN
                           => n146);
   U106 : AOI222_X1 port map( A1 => A2(7), A2 => n84, B1 => A1(7), B2 => n81, 
                           C1 => A3(7), C2 => n78, ZN => n145);
   U107 : INV_X1 port map( A => SEL(2), ZN => n85);
   U108 : NAND2_X1 port map( A1 => n110, A2 => n109, ZN => Y(1));
   U109 : AOI22_X1 port map( A1 => A4(1), A2 => n73, B1 => A0(1), B2 => n2, ZN 
                           => n110);
   U110 : AOI222_X1 port map( A1 => A2(1), A2 => n83, B1 => A1(1), B2 => n79, 
                           C1 => A3(1), C2 => n76, ZN => n109);
   U111 : NAND2_X1 port map( A1 => n138, A2 => n137, ZN => Y(3));
   U112 : AOI22_X1 port map( A1 => A4(3), A2 => n75, B1 => A0(3), B2 => n72, ZN
                           => n138);
   U113 : AOI222_X1 port map( A1 => A2(3), A2 => n84, B1 => A1(3), B2 => n81, 
                           C1 => A3(3), C2 => n78, ZN => n137);
   U114 : NAND2_X1 port map( A1 => n132, A2 => n131, ZN => Y(2));
   U115 : AOI22_X1 port map( A1 => A4(2), A2 => n74, B1 => A0(2), B2 => n2, ZN 
                           => n132);
   U116 : AOI222_X1 port map( A1 => A2(2), A2 => n84, B1 => A1(2), B2 => n80, 
                           C1 => A3(2), C2 => n77, ZN => n131);
   U117 : NAND2_X1 port map( A1 => n88, A2 => n87, ZN => Y(0));
   U118 : AOI22_X1 port map( A1 => A4(0), A2 => n73, B1 => A0(0), B2 => n1, ZN 
                           => n88);
   U119 : AOI222_X1 port map( A1 => A2(0), A2 => n82, B1 => A1(0), B2 => n79, 
                           C1 => A3(0), C2 => n76, ZN => n87);

end SYN_data_fl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity mux51_gen_NBIT32_1 is

   port( A0, A1, A2, A3, A4 : in std_logic_vector (31 downto 0);  SEL : in 
         std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end mux51_gen_NBIT32_1;

architecture SYN_data_fl of mux51_gen_NBIT32_1 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, 
      n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98
      , n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, 
      n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, 
      n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, 
      n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, 
      n147, n148, n149, n150, n151, n152, n153, n154, n155 : std_logic;

begin
   
   U2 : BUF_X1 port map( A => n150, Z => n74);
   U3 : BUF_X1 port map( A => n150, Z => n73);
   U4 : BUF_X1 port map( A => n149, Z => n1);
   U5 : BUF_X1 port map( A => n153, Z => n83);
   U6 : BUF_X1 port map( A => n153, Z => n82);
   U7 : BUF_X1 port map( A => n153, Z => n84);
   U8 : BUF_X1 port map( A => n152, Z => n80);
   U9 : BUF_X1 port map( A => n152, Z => n79);
   U10 : BUF_X1 port map( A => n151, Z => n77);
   U11 : BUF_X1 port map( A => n151, Z => n76);
   U12 : BUF_X1 port map( A => n150, Z => n75);
   U13 : BUF_X1 port map( A => n152, Z => n81);
   U14 : BUF_X1 port map( A => n151, Z => n78);
   U15 : BUF_X1 port map( A => n149, Z => n2);
   U16 : BUF_X1 port map( A => n149, Z => n72);
   U17 : NAND2_X1 port map( A1 => n134, A2 => n133, ZN => Y(30));
   U18 : AOI22_X1 port map( A1 => A4(30), A2 => n74, B1 => A0(30), B2 => n72, 
                           ZN => n134);
   U19 : AOI222_X1 port map( A1 => A2(30), A2 => n84, B1 => A1(30), B2 => n80, 
                           C1 => A3(30), C2 => n77, ZN => n133);
   U20 : NAND2_X1 port map( A1 => n130, A2 => n129, ZN => Y(29));
   U21 : AOI22_X1 port map( A1 => A4(29), A2 => n74, B1 => A0(29), B2 => n2, ZN
                           => n130);
   U22 : AOI222_X1 port map( A1 => A2(29), A2 => n83, B1 => A1(29), B2 => n80, 
                           C1 => A3(29), C2 => n77, ZN => n129);
   U23 : NAND2_X1 port map( A1 => n128, A2 => n127, ZN => Y(28));
   U24 : AOI22_X1 port map( A1 => A4(28), A2 => n74, B1 => A0(28), B2 => n2, ZN
                           => n128);
   U25 : AOI222_X1 port map( A1 => A2(28), A2 => n83, B1 => A1(28), B2 => n80, 
                           C1 => A3(28), C2 => n77, ZN => n127);
   U26 : NAND2_X1 port map( A1 => n126, A2 => n125, ZN => Y(27));
   U27 : AOI22_X1 port map( A1 => A4(27), A2 => n74, B1 => A0(27), B2 => n2, ZN
                           => n126);
   U28 : AOI222_X1 port map( A1 => A2(27), A2 => n83, B1 => A1(27), B2 => n80, 
                           C1 => A3(27), C2 => n77, ZN => n125);
   U29 : NAND2_X1 port map( A1 => n124, A2 => n123, ZN => Y(26));
   U30 : AOI22_X1 port map( A1 => A4(26), A2 => n74, B1 => A0(26), B2 => n2, ZN
                           => n124);
   U31 : AOI222_X1 port map( A1 => A2(26), A2 => n83, B1 => A1(26), B2 => n80, 
                           C1 => A3(26), C2 => n77, ZN => n123);
   U32 : NAND2_X1 port map( A1 => n122, A2 => n121, ZN => Y(25));
   U33 : AOI22_X1 port map( A1 => A4(25), A2 => n74, B1 => A0(25), B2 => n2, ZN
                           => n122);
   U34 : AOI222_X1 port map( A1 => A2(25), A2 => n83, B1 => A1(25), B2 => n80, 
                           C1 => A3(25), C2 => n77, ZN => n121);
   U35 : NAND2_X1 port map( A1 => n120, A2 => n119, ZN => Y(24));
   U36 : AOI22_X1 port map( A1 => A4(24), A2 => n74, B1 => A0(24), B2 => n2, ZN
                           => n120);
   U37 : AOI222_X1 port map( A1 => A2(24), A2 => n83, B1 => A1(24), B2 => n80, 
                           C1 => A3(24), C2 => n77, ZN => n119);
   U38 : NAND2_X1 port map( A1 => n118, A2 => n117, ZN => Y(23));
   U39 : AOI22_X1 port map( A1 => A4(23), A2 => n74, B1 => A0(23), B2 => n2, ZN
                           => n118);
   U40 : AOI222_X1 port map( A1 => A2(23), A2 => n83, B1 => A1(23), B2 => n80, 
                           C1 => A3(23), C2 => n77, ZN => n117);
   U41 : NAND2_X1 port map( A1 => n116, A2 => n115, ZN => Y(22));
   U42 : AOI22_X1 port map( A1 => A4(22), A2 => n74, B1 => A0(22), B2 => n2, ZN
                           => n116);
   U43 : AOI222_X1 port map( A1 => A2(22), A2 => n83, B1 => A1(22), B2 => n80, 
                           C1 => A3(22), C2 => n77, ZN => n115);
   U44 : NAND2_X1 port map( A1 => n114, A2 => n113, ZN => Y(21));
   U45 : AOI22_X1 port map( A1 => A4(21), A2 => n74, B1 => A0(21), B2 => n2, ZN
                           => n114);
   U46 : AOI222_X1 port map( A1 => A2(21), A2 => n83, B1 => A1(21), B2 => n80, 
                           C1 => A3(21), C2 => n77, ZN => n113);
   U47 : NAND2_X1 port map( A1 => n136, A2 => n135, ZN => Y(31));
   U48 : AOI22_X1 port map( A1 => A4(31), A2 => n75, B1 => A0(31), B2 => n72, 
                           ZN => n136);
   U49 : AOI222_X1 port map( A1 => A2(31), A2 => n84, B1 => A1(31), B2 => n81, 
                           C1 => A3(31), C2 => n78, ZN => n135);
   U50 : NAND2_X1 port map( A1 => n112, A2 => n111, ZN => Y(20));
   U51 : AOI22_X1 port map( A1 => A4(20), A2 => n74, B1 => A0(20), B2 => n2, ZN
                           => n112);
   U52 : AOI222_X1 port map( A1 => A2(20), A2 => n83, B1 => A1(20), B2 => n80, 
                           C1 => A3(20), C2 => n77, ZN => n111);
   U53 : NAND2_X1 port map( A1 => n108, A2 => n107, ZN => Y(19));
   U54 : AOI22_X1 port map( A1 => A4(19), A2 => n73, B1 => A0(19), B2 => n1, ZN
                           => n108);
   U55 : AOI222_X1 port map( A1 => A2(19), A2 => n82, B1 => A1(19), B2 => n79, 
                           C1 => A3(19), C2 => n76, ZN => n107);
   U56 : NAND2_X1 port map( A1 => n106, A2 => n105, ZN => Y(18));
   U57 : AOI22_X1 port map( A1 => A4(18), A2 => n73, B1 => A0(18), B2 => n1, ZN
                           => n106);
   U58 : AOI222_X1 port map( A1 => A2(18), A2 => n82, B1 => A1(18), B2 => n79, 
                           C1 => A3(18), C2 => n76, ZN => n105);
   U59 : NAND2_X1 port map( A1 => n104, A2 => n103, ZN => Y(17));
   U60 : AOI22_X1 port map( A1 => A4(17), A2 => n73, B1 => A0(17), B2 => n1, ZN
                           => n104);
   U61 : AOI222_X1 port map( A1 => A2(17), A2 => n82, B1 => A1(17), B2 => n79, 
                           C1 => A3(17), C2 => n76, ZN => n103);
   U62 : NAND2_X1 port map( A1 => n102, A2 => n101, ZN => Y(16));
   U63 : AOI22_X1 port map( A1 => A4(16), A2 => n73, B1 => A0(16), B2 => n1, ZN
                           => n102);
   U64 : AOI222_X1 port map( A1 => A2(16), A2 => n82, B1 => A1(16), B2 => n79, 
                           C1 => A3(16), C2 => n76, ZN => n101);
   U65 : NAND2_X1 port map( A1 => n100, A2 => n99, ZN => Y(15));
   U66 : AOI22_X1 port map( A1 => A4(15), A2 => n73, B1 => A0(15), B2 => n1, ZN
                           => n100);
   U67 : AOI222_X1 port map( A1 => A2(15), A2 => n82, B1 => A1(15), B2 => n79, 
                           C1 => A3(15), C2 => n76, ZN => n99);
   U68 : NAND2_X1 port map( A1 => n98, A2 => n97, ZN => Y(14));
   U69 : AOI22_X1 port map( A1 => A4(14), A2 => n73, B1 => A0(14), B2 => n1, ZN
                           => n98);
   U70 : AOI222_X1 port map( A1 => A2(14), A2 => n82, B1 => A1(14), B2 => n79, 
                           C1 => A3(14), C2 => n76, ZN => n97);
   U71 : NAND2_X1 port map( A1 => n96, A2 => n95, ZN => Y(13));
   U72 : AOI22_X1 port map( A1 => A4(13), A2 => n73, B1 => A0(13), B2 => n1, ZN
                           => n96);
   U73 : AOI222_X1 port map( A1 => A2(13), A2 => n82, B1 => A1(13), B2 => n79, 
                           C1 => A3(13), C2 => n76, ZN => n95);
   U74 : NAND2_X1 port map( A1 => n94, A2 => n93, ZN => Y(12));
   U75 : AOI22_X1 port map( A1 => A4(12), A2 => n73, B1 => A0(12), B2 => n1, ZN
                           => n94);
   U76 : AOI222_X1 port map( A1 => A2(12), A2 => n82, B1 => A1(12), B2 => n79, 
                           C1 => A3(12), C2 => n76, ZN => n93);
   U77 : NAND2_X1 port map( A1 => n92, A2 => n91, ZN => Y(11));
   U78 : AOI22_X1 port map( A1 => A4(11), A2 => n73, B1 => A0(11), B2 => n1, ZN
                           => n92);
   U79 : AOI222_X1 port map( A1 => A2(11), A2 => n82, B1 => A1(11), B2 => n79, 
                           C1 => A3(11), C2 => n76, ZN => n91);
   U80 : NAND2_X1 port map( A1 => n90, A2 => n89, ZN => Y(10));
   U81 : AOI22_X1 port map( A1 => A4(10), A2 => n73, B1 => A0(10), B2 => n1, ZN
                           => n90);
   U82 : AOI222_X1 port map( A1 => A2(10), A2 => n82, B1 => A1(10), B2 => n79, 
                           C1 => A3(10), C2 => n76, ZN => n89);
   U83 : NAND2_X1 port map( A1 => n155, A2 => n154, ZN => Y(9));
   U84 : AOI22_X1 port map( A1 => A4(9), A2 => n75, B1 => A0(9), B2 => n72, ZN 
                           => n155);
   U85 : AOI222_X1 port map( A1 => A2(9), A2 => n84, B1 => A1(9), B2 => n81, C1
                           => A3(9), C2 => n78, ZN => n154);
   U86 : NAND2_X1 port map( A1 => n148, A2 => n147, ZN => Y(8));
   U87 : AOI22_X1 port map( A1 => A4(8), A2 => n75, B1 => A0(8), B2 => n72, ZN 
                           => n148);
   U88 : AOI222_X1 port map( A1 => A2(8), A2 => n84, B1 => A1(8), B2 => n81, C1
                           => A3(8), C2 => n78, ZN => n147);
   U89 : NAND2_X1 port map( A1 => n146, A2 => n145, ZN => Y(7));
   U90 : AOI22_X1 port map( A1 => A4(7), A2 => n75, B1 => A0(7), B2 => n72, ZN 
                           => n146);
   U91 : AOI222_X1 port map( A1 => A2(7), A2 => n84, B1 => A1(7), B2 => n81, C1
                           => A3(7), C2 => n78, ZN => n145);
   U92 : NAND2_X1 port map( A1 => n138, A2 => n137, ZN => Y(3));
   U93 : AOI22_X1 port map( A1 => A4(3), A2 => n75, B1 => A0(3), B2 => n72, ZN 
                           => n138);
   U94 : AOI222_X1 port map( A1 => A2(3), A2 => n84, B1 => A1(3), B2 => n81, C1
                           => A3(3), C2 => n78, ZN => n137);
   U95 : NOR3_X1 port map( A1 => SEL(0), A2 => SEL(1), A3 => n1, ZN => n150);
   U96 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => SEL(0), ZN => n149
                           );
   U97 : NOR3_X1 port map( A1 => SEL(0), A2 => SEL(2), A3 => n86, ZN => n153);
   U98 : NAND2_X1 port map( A1 => n142, A2 => n141, ZN => Y(5));
   U99 : AOI222_X1 port map( A1 => A2(5), A2 => n84, B1 => A1(5), B2 => n81, C1
                           => A3(5), C2 => n78, ZN => n141);
   U100 : AOI22_X1 port map( A1 => A4(5), A2 => n75, B1 => A0(5), B2 => n72, ZN
                           => n142);
   U101 : NAND2_X1 port map( A1 => n140, A2 => n139, ZN => Y(4));
   U102 : AOI222_X1 port map( A1 => A2(4), A2 => n84, B1 => A1(4), B2 => n81, 
                           C1 => A3(4), C2 => n78, ZN => n139);
   U103 : AOI22_X1 port map( A1 => A4(4), A2 => n75, B1 => A0(4), B2 => n72, ZN
                           => n140);
   U104 : AND3_X1 port map( A1 => SEL(0), A2 => n85, A3 => SEL(1), ZN => n151);
   U105 : AND3_X1 port map( A1 => n86, A2 => n85, A3 => SEL(0), ZN => n152);
   U106 : INV_X1 port map( A => SEL(1), ZN => n86);
   U107 : NAND2_X1 port map( A1 => n144, A2 => n143, ZN => Y(6));
   U108 : AOI22_X1 port map( A1 => A4(6), A2 => n75, B1 => A0(6), B2 => n72, ZN
                           => n144);
   U109 : AOI222_X1 port map( A1 => A2(6), A2 => n84, B1 => A1(6), B2 => n81, 
                           C1 => A3(6), C2 => n78, ZN => n143);
   U110 : INV_X1 port map( A => SEL(2), ZN => n85);
   U111 : NAND2_X1 port map( A1 => n110, A2 => n109, ZN => Y(1));
   U112 : AOI22_X1 port map( A1 => A4(1), A2 => n73, B1 => A0(1), B2 => n2, ZN 
                           => n110);
   U113 : AOI222_X1 port map( A1 => A2(1), A2 => n83, B1 => A1(1), B2 => n79, 
                           C1 => A3(1), C2 => n76, ZN => n109);
   U114 : NAND2_X1 port map( A1 => n132, A2 => n131, ZN => Y(2));
   U115 : AOI22_X1 port map( A1 => A4(2), A2 => n74, B1 => A0(2), B2 => n2, ZN 
                           => n132);
   U116 : AOI222_X1 port map( A1 => A2(2), A2 => n84, B1 => A1(2), B2 => n80, 
                           C1 => A3(2), C2 => n77, ZN => n131);
   U117 : NAND2_X1 port map( A1 => n88, A2 => n87, ZN => Y(0));
   U118 : AOI22_X1 port map( A1 => A4(0), A2 => n73, B1 => A0(0), B2 => n1, ZN 
                           => n88);
   U119 : AOI222_X1 port map( A1 => A2(0), A2 => n82, B1 => A1(0), B2 => n79, 
                           C1 => A3(0), C2 => n76, ZN => n87);

end SYN_data_fl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity negate_NBIT32_7 is

   port( A : in std_logic_vector (31 downto 0);  Y : out std_logic_vector (31 
         downto 0));

end negate_NBIT32_7;

architecture SYN_data_fl of negate_NBIT32_7 is

   component negate_NBIT32_7_DW01_sub_0
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  DIFF
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   signal n3, n4, n_1439 : std_logic;

begin
   
   n4 <= '0';
   n3 <= '0';
   sub_add_14_b0 : negate_NBIT32_7_DW01_sub_0 port map( A(31) => n4, A(30) => 
                           n4, A(29) => n4, A(28) => n4, A(27) => n4, A(26) => 
                           n4, A(25) => n4, A(24) => n4, A(23) => n4, A(22) => 
                           n4, A(21) => n4, A(20) => n4, A(19) => n4, A(18) => 
                           n4, A(17) => n4, A(16) => n4, A(15) => n4, A(14) => 
                           n4, A(13) => n4, A(12) => n4, A(11) => n4, A(10) => 
                           n4, A(9) => n4, A(8) => n4, A(7) => n4, A(6) => n4, 
                           A(5) => n4, A(4) => n4, A(3) => n4, A(2) => n4, A(1)
                           => n4, A(0) => n4, B(31) => A(31), B(30) => A(30), 
                           B(29) => A(29), B(28) => A(28), B(27) => A(27), 
                           B(26) => A(26), B(25) => A(25), B(24) => A(24), 
                           B(23) => A(23), B(22) => A(22), B(21) => A(21), 
                           B(20) => A(20), B(19) => A(19), B(18) => A(18), 
                           B(17) => A(17), B(16) => A(16), B(15) => A(15), 
                           B(14) => A(14), B(13) => A(13), B(12) => A(12), 
                           B(11) => A(11), B(10) => A(10), B(9) => A(9), B(8) 
                           => A(8), B(7) => A(7), B(6) => A(6), B(5) => A(5), 
                           B(4) => A(4), B(3) => A(3), B(2) => A(2), B(1) => 
                           A(1), B(0) => A(0), CI => n3, DIFF(31) => Y(31), 
                           DIFF(30) => Y(30), DIFF(29) => Y(29), DIFF(28) => 
                           Y(28), DIFF(27) => Y(27), DIFF(26) => Y(26), 
                           DIFF(25) => Y(25), DIFF(24) => Y(24), DIFF(23) => 
                           Y(23), DIFF(22) => Y(22), DIFF(21) => Y(21), 
                           DIFF(20) => Y(20), DIFF(19) => Y(19), DIFF(18) => 
                           Y(18), DIFF(17) => Y(17), DIFF(16) => Y(16), 
                           DIFF(15) => Y(15), DIFF(14) => Y(14), DIFF(13) => 
                           Y(13), DIFF(12) => Y(12), DIFF(11) => Y(11), 
                           DIFF(10) => Y(10), DIFF(9) => Y(9), DIFF(8) => Y(8),
                           DIFF(7) => Y(7), DIFF(6) => Y(6), DIFF(5) => Y(5), 
                           DIFF(4) => Y(4), DIFF(3) => Y(3), DIFF(2) => Y(2), 
                           DIFF(1) => Y(1), DIFF(0) => Y(0), CO => n_1439);

end SYN_data_fl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity negate_NBIT32_6 is

   port( A : in std_logic_vector (31 downto 0);  Y : out std_logic_vector (31 
         downto 0));

end negate_NBIT32_6;

architecture SYN_data_fl of negate_NBIT32_6 is

   component negate_NBIT32_6_DW01_sub_0
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  DIFF
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   signal n3, n4, n_1440 : std_logic;

begin
   
   n4 <= '0';
   n3 <= '0';
   sub_add_14_b0 : negate_NBIT32_6_DW01_sub_0 port map( A(31) => n4, A(30) => 
                           n4, A(29) => n4, A(28) => n4, A(27) => n4, A(26) => 
                           n4, A(25) => n4, A(24) => n4, A(23) => n4, A(22) => 
                           n4, A(21) => n4, A(20) => n4, A(19) => n4, A(18) => 
                           n4, A(17) => n4, A(16) => n4, A(15) => n4, A(14) => 
                           n4, A(13) => n4, A(12) => n4, A(11) => n4, A(10) => 
                           n4, A(9) => n4, A(8) => n4, A(7) => n4, A(6) => n4, 
                           A(5) => n4, A(4) => n4, A(3) => n4, A(2) => n4, A(1)
                           => n4, A(0) => n4, B(31) => A(31), B(30) => A(30), 
                           B(29) => A(29), B(28) => A(28), B(27) => A(27), 
                           B(26) => A(26), B(25) => A(25), B(24) => A(24), 
                           B(23) => A(23), B(22) => A(22), B(21) => A(21), 
                           B(20) => A(20), B(19) => A(19), B(18) => A(18), 
                           B(17) => A(17), B(16) => A(16), B(15) => A(15), 
                           B(14) => A(14), B(13) => A(13), B(12) => A(12), 
                           B(11) => A(11), B(10) => A(10), B(9) => A(9), B(8) 
                           => A(8), B(7) => A(7), B(6) => A(6), B(5) => A(5), 
                           B(4) => A(4), B(3) => A(3), B(2) => A(2), B(1) => 
                           A(1), B(0) => A(0), CI => n3, DIFF(31) => Y(31), 
                           DIFF(30) => Y(30), DIFF(29) => Y(29), DIFF(28) => 
                           Y(28), DIFF(27) => Y(27), DIFF(26) => Y(26), 
                           DIFF(25) => Y(25), DIFF(24) => Y(24), DIFF(23) => 
                           Y(23), DIFF(22) => Y(22), DIFF(21) => Y(21), 
                           DIFF(20) => Y(20), DIFF(19) => Y(19), DIFF(18) => 
                           Y(18), DIFF(17) => Y(17), DIFF(16) => Y(16), 
                           DIFF(15) => Y(15), DIFF(14) => Y(14), DIFF(13) => 
                           Y(13), DIFF(12) => Y(12), DIFF(11) => Y(11), 
                           DIFF(10) => Y(10), DIFF(9) => Y(9), DIFF(8) => Y(8),
                           DIFF(7) => Y(7), DIFF(6) => Y(6), DIFF(5) => Y(5), 
                           DIFF(4) => Y(4), DIFF(3) => Y(3), DIFF(2) => Y(2), 
                           DIFF(1) => Y(1), DIFF(0) => Y(0), CO => n_1440);

end SYN_data_fl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity negate_NBIT32_5 is

   port( A : in std_logic_vector (31 downto 0);  Y : out std_logic_vector (31 
         downto 0));

end negate_NBIT32_5;

architecture SYN_data_fl of negate_NBIT32_5 is

   component negate_NBIT32_5_DW01_sub_0
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  DIFF
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   signal n3, n4, n_1441 : std_logic;

begin
   
   n4 <= '0';
   n3 <= '0';
   sub_add_14_b0 : negate_NBIT32_5_DW01_sub_0 port map( A(31) => n4, A(30) => 
                           n4, A(29) => n4, A(28) => n4, A(27) => n4, A(26) => 
                           n4, A(25) => n4, A(24) => n4, A(23) => n4, A(22) => 
                           n4, A(21) => n4, A(20) => n4, A(19) => n4, A(18) => 
                           n4, A(17) => n4, A(16) => n4, A(15) => n4, A(14) => 
                           n4, A(13) => n4, A(12) => n4, A(11) => n4, A(10) => 
                           n4, A(9) => n4, A(8) => n4, A(7) => n4, A(6) => n4, 
                           A(5) => n4, A(4) => n4, A(3) => n4, A(2) => n4, A(1)
                           => n4, A(0) => n4, B(31) => A(31), B(30) => A(30), 
                           B(29) => A(29), B(28) => A(28), B(27) => A(27), 
                           B(26) => A(26), B(25) => A(25), B(24) => A(24), 
                           B(23) => A(23), B(22) => A(22), B(21) => A(21), 
                           B(20) => A(20), B(19) => A(19), B(18) => A(18), 
                           B(17) => A(17), B(16) => A(16), B(15) => A(15), 
                           B(14) => A(14), B(13) => A(13), B(12) => A(12), 
                           B(11) => A(11), B(10) => A(10), B(9) => A(9), B(8) 
                           => A(8), B(7) => A(7), B(6) => A(6), B(5) => A(5), 
                           B(4) => A(4), B(3) => A(3), B(2) => A(2), B(1) => 
                           A(1), B(0) => A(0), CI => n3, DIFF(31) => Y(31), 
                           DIFF(30) => Y(30), DIFF(29) => Y(29), DIFF(28) => 
                           Y(28), DIFF(27) => Y(27), DIFF(26) => Y(26), 
                           DIFF(25) => Y(25), DIFF(24) => Y(24), DIFF(23) => 
                           Y(23), DIFF(22) => Y(22), DIFF(21) => Y(21), 
                           DIFF(20) => Y(20), DIFF(19) => Y(19), DIFF(18) => 
                           Y(18), DIFF(17) => Y(17), DIFF(16) => Y(16), 
                           DIFF(15) => Y(15), DIFF(14) => Y(14), DIFF(13) => 
                           Y(13), DIFF(12) => Y(12), DIFF(11) => Y(11), 
                           DIFF(10) => Y(10), DIFF(9) => Y(9), DIFF(8) => Y(8),
                           DIFF(7) => Y(7), DIFF(6) => Y(6), DIFF(5) => Y(5), 
                           DIFF(4) => Y(4), DIFF(3) => Y(3), DIFF(2) => Y(2), 
                           DIFF(1) => Y(1), DIFF(0) => Y(0), CO => n_1441);

end SYN_data_fl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity negate_NBIT32_4 is

   port( A : in std_logic_vector (31 downto 0);  Y : out std_logic_vector (31 
         downto 0));

end negate_NBIT32_4;

architecture SYN_data_fl of negate_NBIT32_4 is

   component negate_NBIT32_4_DW01_sub_0
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  DIFF
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   signal n3, n4, n_1442 : std_logic;

begin
   
   n4 <= '0';
   n3 <= '0';
   sub_add_14_b0 : negate_NBIT32_4_DW01_sub_0 port map( A(31) => n4, A(30) => 
                           n4, A(29) => n4, A(28) => n4, A(27) => n4, A(26) => 
                           n4, A(25) => n4, A(24) => n4, A(23) => n4, A(22) => 
                           n4, A(21) => n4, A(20) => n4, A(19) => n4, A(18) => 
                           n4, A(17) => n4, A(16) => n4, A(15) => n4, A(14) => 
                           n4, A(13) => n4, A(12) => n4, A(11) => n4, A(10) => 
                           n4, A(9) => n4, A(8) => n4, A(7) => n4, A(6) => n4, 
                           A(5) => n4, A(4) => n4, A(3) => n4, A(2) => n4, A(1)
                           => n4, A(0) => n4, B(31) => A(31), B(30) => A(30), 
                           B(29) => A(29), B(28) => A(28), B(27) => A(27), 
                           B(26) => A(26), B(25) => A(25), B(24) => A(24), 
                           B(23) => A(23), B(22) => A(22), B(21) => A(21), 
                           B(20) => A(20), B(19) => A(19), B(18) => A(18), 
                           B(17) => A(17), B(16) => A(16), B(15) => A(15), 
                           B(14) => A(14), B(13) => A(13), B(12) => A(12), 
                           B(11) => A(11), B(10) => A(10), B(9) => A(9), B(8) 
                           => A(8), B(7) => A(7), B(6) => A(6), B(5) => A(5), 
                           B(4) => A(4), B(3) => A(3), B(2) => A(2), B(1) => 
                           A(1), B(0) => A(0), CI => n3, DIFF(31) => Y(31), 
                           DIFF(30) => Y(30), DIFF(29) => Y(29), DIFF(28) => 
                           Y(28), DIFF(27) => Y(27), DIFF(26) => Y(26), 
                           DIFF(25) => Y(25), DIFF(24) => Y(24), DIFF(23) => 
                           Y(23), DIFF(22) => Y(22), DIFF(21) => Y(21), 
                           DIFF(20) => Y(20), DIFF(19) => Y(19), DIFF(18) => 
                           Y(18), DIFF(17) => Y(17), DIFF(16) => Y(16), 
                           DIFF(15) => Y(15), DIFF(14) => Y(14), DIFF(13) => 
                           Y(13), DIFF(12) => Y(12), DIFF(11) => Y(11), 
                           DIFF(10) => Y(10), DIFF(9) => Y(9), DIFF(8) => Y(8),
                           DIFF(7) => Y(7), DIFF(6) => Y(6), DIFF(5) => Y(5), 
                           DIFF(4) => Y(4), DIFF(3) => Y(3), DIFF(2) => Y(2), 
                           DIFF(1) => Y(1), DIFF(0) => Y(0), CO => n_1442);

end SYN_data_fl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity negate_NBIT32_3 is

   port( A : in std_logic_vector (31 downto 0);  Y : out std_logic_vector (31 
         downto 0));

end negate_NBIT32_3;

architecture SYN_data_fl of negate_NBIT32_3 is

   component negate_NBIT32_3_DW01_sub_0
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  DIFF
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   signal n3, n4, n_1443 : std_logic;

begin
   
   n4 <= '0';
   n3 <= '0';
   sub_add_14_b0 : negate_NBIT32_3_DW01_sub_0 port map( A(31) => n4, A(30) => 
                           n4, A(29) => n4, A(28) => n4, A(27) => n4, A(26) => 
                           n4, A(25) => n4, A(24) => n4, A(23) => n4, A(22) => 
                           n4, A(21) => n4, A(20) => n4, A(19) => n4, A(18) => 
                           n4, A(17) => n4, A(16) => n4, A(15) => n4, A(14) => 
                           n4, A(13) => n4, A(12) => n4, A(11) => n4, A(10) => 
                           n4, A(9) => n4, A(8) => n4, A(7) => n4, A(6) => n4, 
                           A(5) => n4, A(4) => n4, A(3) => n4, A(2) => n4, A(1)
                           => n4, A(0) => n4, B(31) => A(31), B(30) => A(30), 
                           B(29) => A(29), B(28) => A(28), B(27) => A(27), 
                           B(26) => A(26), B(25) => A(25), B(24) => A(24), 
                           B(23) => A(23), B(22) => A(22), B(21) => A(21), 
                           B(20) => A(20), B(19) => A(19), B(18) => A(18), 
                           B(17) => A(17), B(16) => A(16), B(15) => A(15), 
                           B(14) => A(14), B(13) => A(13), B(12) => A(12), 
                           B(11) => A(11), B(10) => A(10), B(9) => A(9), B(8) 
                           => A(8), B(7) => A(7), B(6) => A(6), B(5) => A(5), 
                           B(4) => A(4), B(3) => A(3), B(2) => A(2), B(1) => 
                           A(1), B(0) => A(0), CI => n3, DIFF(31) => Y(31), 
                           DIFF(30) => Y(30), DIFF(29) => Y(29), DIFF(28) => 
                           Y(28), DIFF(27) => Y(27), DIFF(26) => Y(26), 
                           DIFF(25) => Y(25), DIFF(24) => Y(24), DIFF(23) => 
                           Y(23), DIFF(22) => Y(22), DIFF(21) => Y(21), 
                           DIFF(20) => Y(20), DIFF(19) => Y(19), DIFF(18) => 
                           Y(18), DIFF(17) => Y(17), DIFF(16) => Y(16), 
                           DIFF(15) => Y(15), DIFF(14) => Y(14), DIFF(13) => 
                           Y(13), DIFF(12) => Y(12), DIFF(11) => Y(11), 
                           DIFF(10) => Y(10), DIFF(9) => Y(9), DIFF(8) => Y(8),
                           DIFF(7) => Y(7), DIFF(6) => Y(6), DIFF(5) => Y(5), 
                           DIFF(4) => Y(4), DIFF(3) => Y(3), DIFF(2) => Y(2), 
                           DIFF(1) => Y(1), DIFF(0) => Y(0), CO => n_1443);

end SYN_data_fl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity negate_NBIT32_2 is

   port( A : in std_logic_vector (31 downto 0);  Y : out std_logic_vector (31 
         downto 0));

end negate_NBIT32_2;

architecture SYN_data_fl of negate_NBIT32_2 is

   component negate_NBIT32_2_DW01_sub_0
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  DIFF
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   signal n3, n4, n_1444 : std_logic;

begin
   
   n4 <= '0';
   n3 <= '0';
   sub_add_14_b0 : negate_NBIT32_2_DW01_sub_0 port map( A(31) => n4, A(30) => 
                           n4, A(29) => n4, A(28) => n4, A(27) => n4, A(26) => 
                           n4, A(25) => n4, A(24) => n4, A(23) => n4, A(22) => 
                           n4, A(21) => n4, A(20) => n4, A(19) => n4, A(18) => 
                           n4, A(17) => n4, A(16) => n4, A(15) => n4, A(14) => 
                           n4, A(13) => n4, A(12) => n4, A(11) => n4, A(10) => 
                           n4, A(9) => n4, A(8) => n4, A(7) => n4, A(6) => n4, 
                           A(5) => n4, A(4) => n4, A(3) => n4, A(2) => n4, A(1)
                           => n4, A(0) => n4, B(31) => A(31), B(30) => A(30), 
                           B(29) => A(29), B(28) => A(28), B(27) => A(27), 
                           B(26) => A(26), B(25) => A(25), B(24) => A(24), 
                           B(23) => A(23), B(22) => A(22), B(21) => A(21), 
                           B(20) => A(20), B(19) => A(19), B(18) => A(18), 
                           B(17) => A(17), B(16) => A(16), B(15) => A(15), 
                           B(14) => A(14), B(13) => A(13), B(12) => A(12), 
                           B(11) => A(11), B(10) => A(10), B(9) => A(9), B(8) 
                           => A(8), B(7) => A(7), B(6) => A(6), B(5) => A(5), 
                           B(4) => A(4), B(3) => A(3), B(2) => A(2), B(1) => 
                           A(1), B(0) => A(0), CI => n3, DIFF(31) => Y(31), 
                           DIFF(30) => Y(30), DIFF(29) => Y(29), DIFF(28) => 
                           Y(28), DIFF(27) => Y(27), DIFF(26) => Y(26), 
                           DIFF(25) => Y(25), DIFF(24) => Y(24), DIFF(23) => 
                           Y(23), DIFF(22) => Y(22), DIFF(21) => Y(21), 
                           DIFF(20) => Y(20), DIFF(19) => Y(19), DIFF(18) => 
                           Y(18), DIFF(17) => Y(17), DIFF(16) => Y(16), 
                           DIFF(15) => Y(15), DIFF(14) => Y(14), DIFF(13) => 
                           Y(13), DIFF(12) => Y(12), DIFF(11) => Y(11), 
                           DIFF(10) => Y(10), DIFF(9) => Y(9), DIFF(8) => Y(8),
                           DIFF(7) => Y(7), DIFF(6) => Y(6), DIFF(5) => Y(5), 
                           DIFF(4) => Y(4), DIFF(3) => Y(3), DIFF(2) => Y(2), 
                           DIFF(1) => Y(1), DIFF(0) => Y(0), CO => n_1444);

end SYN_data_fl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity negate_NBIT32_1 is

   port( A : in std_logic_vector (31 downto 0);  Y : out std_logic_vector (31 
         downto 0));

end negate_NBIT32_1;

architecture SYN_data_fl of negate_NBIT32_1 is

   component negate_NBIT32_1_DW01_sub_0
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  DIFF
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   signal n3, n4, n_1445 : std_logic;

begin
   
   n4 <= '0';
   n3 <= '0';
   sub_add_14_b0 : negate_NBIT32_1_DW01_sub_0 port map( A(31) => n4, A(30) => 
                           n4, A(29) => n4, A(28) => n4, A(27) => n4, A(26) => 
                           n4, A(25) => n4, A(24) => n4, A(23) => n4, A(22) => 
                           n4, A(21) => n4, A(20) => n4, A(19) => n4, A(18) => 
                           n4, A(17) => n4, A(16) => n4, A(15) => n4, A(14) => 
                           n4, A(13) => n4, A(12) => n4, A(11) => n4, A(10) => 
                           n4, A(9) => n4, A(8) => n4, A(7) => n4, A(6) => n4, 
                           A(5) => n4, A(4) => n4, A(3) => n4, A(2) => n4, A(1)
                           => n4, A(0) => n4, B(31) => A(31), B(30) => A(30), 
                           B(29) => A(29), B(28) => A(28), B(27) => A(27), 
                           B(26) => A(26), B(25) => A(25), B(24) => A(24), 
                           B(23) => A(23), B(22) => A(22), B(21) => A(21), 
                           B(20) => A(20), B(19) => A(19), B(18) => A(18), 
                           B(17) => A(17), B(16) => A(16), B(15) => A(15), 
                           B(14) => A(14), B(13) => A(13), B(12) => A(12), 
                           B(11) => A(11), B(10) => A(10), B(9) => A(9), B(8) 
                           => A(8), B(7) => A(7), B(6) => A(6), B(5) => A(5), 
                           B(4) => A(4), B(3) => A(3), B(2) => A(2), B(1) => 
                           A(1), B(0) => A(0), CI => n3, DIFF(31) => Y(31), 
                           DIFF(30) => Y(30), DIFF(29) => Y(29), DIFF(28) => 
                           Y(28), DIFF(27) => Y(27), DIFF(26) => Y(26), 
                           DIFF(25) => Y(25), DIFF(24) => Y(24), DIFF(23) => 
                           Y(23), DIFF(22) => Y(22), DIFF(21) => Y(21), 
                           DIFF(20) => Y(20), DIFF(19) => Y(19), DIFF(18) => 
                           Y(18), DIFF(17) => Y(17), DIFF(16) => Y(16), 
                           DIFF(15) => Y(15), DIFF(14) => Y(14), DIFF(13) => 
                           Y(13), DIFF(12) => Y(12), DIFF(11) => Y(11), 
                           DIFF(10) => Y(10), DIFF(9) => Y(9), DIFF(8) => Y(8),
                           DIFF(7) => Y(7), DIFF(6) => Y(6), DIFF(5) => Y(5), 
                           DIFF(4) => Y(4), DIFF(3) => Y(3), DIFF(2) => Y(2), 
                           DIFF(1) => Y(1), DIFF(0) => Y(0), CO => n_1445);

end SYN_data_fl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity shl2_NBIT32_2 is

   port( A : in std_logic_vector (31 downto 0);  Y : out std_logic_vector (31 
         downto 0));

end shl2_NBIT32_2;

architecture SYN_behavioral of shl2_NBIT32_2 is

signal X_Logic0_port : std_logic;

begin
   Y <= ( A(29), A(28), A(27), A(26), A(25), A(24), A(23), A(22), A(21), A(20),
      A(19), A(18), A(17), A(16), A(15), A(14), A(13), A(12), A(11), A(10), 
      A(9), A(8), A(7), A(6), A(5), A(4), A(3), A(2), A(1), A(0), X_Logic0_port
      , X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity shl2_NBIT32_1 is

   port( A : in std_logic_vector (31 downto 0);  Y : out std_logic_vector (31 
         downto 0));

end shl2_NBIT32_1;

architecture SYN_behavioral of shl2_NBIT32_1 is

signal X_Logic0_port : std_logic;

begin
   Y <= ( A(29), A(28), A(27), A(26), A(25), A(24), A(23), A(22), A(21), A(20),
      A(19), A(18), A(17), A(16), A(15), A(14), A(13), A(12), A(11), A(10), 
      A(9), A(8), A(7), A(6), A(5), A(4), A(3), A(2), A(1), A(0), X_Logic0_port
      , X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity shl1_NBIT32_2 is

   port( A : in std_logic_vector (31 downto 0);  Y : out std_logic_vector (31 
         downto 0));

end shl1_NBIT32_2;

architecture SYN_datafl of shl1_NBIT32_2 is

signal X_Logic0_port : std_logic;

begin
   Y <= ( A(30), A(29), A(28), A(27), A(26), A(25), A(24), A(23), A(22), A(21),
      A(20), A(19), A(18), A(17), A(16), A(15), A(14), A(13), A(12), A(11), 
      A(10), A(9), A(8), A(7), A(6), A(5), A(4), A(3), A(2), A(1), A(0), 
      X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_datafl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity shl1_NBIT32_1 is

   port( A : in std_logic_vector (31 downto 0);  Y : out std_logic_vector (31 
         downto 0));

end shl1_NBIT32_1;

architecture SYN_datafl of shl1_NBIT32_1 is

signal X_Logic0_port : std_logic;

begin
   Y <= ( A(30), A(29), A(28), A(27), A(26), A(25), A(24), A(23), A(22), A(21),
      A(20), A(19), A(18), A(17), A(16), A(15), A(14), A(13), A(12), A(11), 
      A(10), A(9), A(8), A(7), A(6), A(5), A(4), A(3), A(2), A(1), A(0), 
      X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_datafl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity enc33_3 is

   port( A : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (2 
         downto 0));

end enc33_3;

architecture SYN_behavioral of enc33_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n7, n8, n9 : std_logic;

begin
   
   U8 : XOR2_X1 port map( A => A(0), B => A(1), Z => n8);
   U1 : NOR3_X1 port map( A1 => n1, A2 => n9, A3 => n8, ZN => Y(2));
   U2 : OAI21_X1 port map( B1 => n2, B2 => n1, A => n7, ZN => Y(1));
   U3 : NAND2_X1 port map( A1 => n9, A2 => n1, ZN => n7);
   U4 : INV_X1 port map( A => n8, ZN => n2);
   U5 : OAI21_X1 port map( B1 => A(2), B2 => n2, A => n7, ZN => Y(0));
   U6 : AND2_X1 port map( A1 => A(1), A2 => A(0), ZN => n9);
   U7 : INV_X1 port map( A => A(2), ZN => n1);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity enc33_2 is

   port( A : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (2 
         downto 0));

end enc33_2;

architecture SYN_behavioral of enc33_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n7, n8, n9 : std_logic;

begin
   
   U8 : XOR2_X1 port map( A => A(0), B => A(1), Z => n8);
   U1 : NOR3_X1 port map( A1 => n2, A2 => n9, A3 => n8, ZN => Y(2));
   U2 : INV_X1 port map( A => n8, ZN => n1);
   U3 : NAND2_X1 port map( A1 => n9, A2 => n2, ZN => n7);
   U4 : OAI21_X1 port map( B1 => n1, B2 => n2, A => n7, ZN => Y(1));
   U5 : INV_X1 port map( A => A(2), ZN => n2);
   U6 : OAI21_X1 port map( B1 => A(2), B2 => n1, A => n7, ZN => Y(0));
   U7 : AND2_X1 port map( A1 => A(1), A2 => A(0), ZN => n9);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity enc33_1 is

   port( A : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (2 
         downto 0));

end enc33_1;

architecture SYN_behavioral of enc33_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n7, n8, n9 : std_logic;

begin
   
   U8 : XOR2_X1 port map( A => A(0), B => A(1), Z => n8);
   U1 : NOR3_X1 port map( A1 => n2, A2 => n9, A3 => n8, ZN => Y(2));
   U2 : INV_X1 port map( A => n8, ZN => n1);
   U3 : OAI21_X1 port map( B1 => n1, B2 => n2, A => n7, ZN => Y(1));
   U4 : NAND2_X1 port map( A1 => n9, A2 => n2, ZN => n7);
   U5 : INV_X1 port map( A => A(2), ZN => n2);
   U6 : OAI21_X1 port map( B1 => A(2), B2 => n1, A => n7, ZN => Y(0));
   U7 : AND2_X1 port map( A1 => A(1), A2 => A(0), ZN => n9);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_63 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_63;

architecture SYN_STRUCTURAL of carry_select_block_n4_63 is

   component MUX21_GENERIC_NBIT4_63
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_125
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_126
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1446, 
      n_1447 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_126 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1446);
   RCA1 : RCA_GEN_NBIT4_125 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1447);
   mux : MUX21_GENERIC_NBIT4_63 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_62 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_62;

architecture SYN_STRUCTURAL of carry_select_block_n4_62 is

   component MUX21_GENERIC_NBIT4_62
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_123
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_124
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1448, 
      n_1449 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_124 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1448);
   RCA1 : RCA_GEN_NBIT4_123 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1449);
   mux : MUX21_GENERIC_NBIT4_62 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_61 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_61;

architecture SYN_STRUCTURAL of carry_select_block_n4_61 is

   component MUX21_GENERIC_NBIT4_61
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_121
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_122
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1450, 
      n_1451 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_122 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1450);
   RCA1 : RCA_GEN_NBIT4_121 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1451);
   mux : MUX21_GENERIC_NBIT4_61 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_60 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_60;

architecture SYN_STRUCTURAL of carry_select_block_n4_60 is

   component MUX21_GENERIC_NBIT4_60
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_119
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_120
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1452, 
      n_1453 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_120 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1452);
   RCA1 : RCA_GEN_NBIT4_119 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1453);
   mux : MUX21_GENERIC_NBIT4_60 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_59 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_59;

architecture SYN_STRUCTURAL of carry_select_block_n4_59 is

   component MUX21_GENERIC_NBIT4_59
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_117
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_118
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1454, 
      n_1455 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_118 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1454);
   RCA1 : RCA_GEN_NBIT4_117 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1455);
   mux : MUX21_GENERIC_NBIT4_59 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_58 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_58;

architecture SYN_STRUCTURAL of carry_select_block_n4_58 is

   component MUX21_GENERIC_NBIT4_58
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_115
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_116
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1456, 
      n_1457 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_116 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1456);
   RCA1 : RCA_GEN_NBIT4_115 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1457);
   mux : MUX21_GENERIC_NBIT4_58 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_57 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_57;

architecture SYN_STRUCTURAL of carry_select_block_n4_57 is

   component MUX21_GENERIC_NBIT4_57
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_113
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_114
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1458, 
      n_1459 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_114 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1458);
   RCA1 : RCA_GEN_NBIT4_113 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1459);
   mux : MUX21_GENERIC_NBIT4_57 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_56 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_56;

architecture SYN_STRUCTURAL of carry_select_block_n4_56 is

   component MUX21_GENERIC_NBIT4_56
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_111
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_112
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1460, 
      n_1461 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_112 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1460);
   RCA1 : RCA_GEN_NBIT4_111 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1461);
   mux : MUX21_GENERIC_NBIT4_56 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_55 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_55;

architecture SYN_STRUCTURAL of carry_select_block_n4_55 is

   component MUX21_GENERIC_NBIT4_55
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_109
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_110
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1462, 
      n_1463 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_110 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1462);
   RCA1 : RCA_GEN_NBIT4_109 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1463);
   mux : MUX21_GENERIC_NBIT4_55 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_54 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_54;

architecture SYN_STRUCTURAL of carry_select_block_n4_54 is

   component MUX21_GENERIC_NBIT4_54
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_107
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_108
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1464, 
      n_1465 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_108 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1464);
   RCA1 : RCA_GEN_NBIT4_107 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1465);
   mux : MUX21_GENERIC_NBIT4_54 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_53 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_53;

architecture SYN_STRUCTURAL of carry_select_block_n4_53 is

   component MUX21_GENERIC_NBIT4_53
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_105
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_106
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1466, 
      n_1467 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_106 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1466);
   RCA1 : RCA_GEN_NBIT4_105 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1467);
   mux : MUX21_GENERIC_NBIT4_53 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_52 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_52;

architecture SYN_STRUCTURAL of carry_select_block_n4_52 is

   component MUX21_GENERIC_NBIT4_52
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_103
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_104
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1468, 
      n_1469 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_104 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1468);
   RCA1 : RCA_GEN_NBIT4_103 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1469);
   mux : MUX21_GENERIC_NBIT4_52 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_51 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_51;

architecture SYN_STRUCTURAL of carry_select_block_n4_51 is

   component MUX21_GENERIC_NBIT4_51
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_101
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_102
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1470, 
      n_1471 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_102 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1470);
   RCA1 : RCA_GEN_NBIT4_101 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1471);
   mux : MUX21_GENERIC_NBIT4_51 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_50 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_50;

architecture SYN_STRUCTURAL of carry_select_block_n4_50 is

   component MUX21_GENERIC_NBIT4_50
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_99
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_100
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1472, 
      n_1473 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_100 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1472);
   RCA1 : RCA_GEN_NBIT4_99 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1473);
   mux : MUX21_GENERIC_NBIT4_50 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_49 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_49;

architecture SYN_STRUCTURAL of carry_select_block_n4_49 is

   component MUX21_GENERIC_NBIT4_49
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_97
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_98
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1474, 
      n_1475 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_98 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1474);
   RCA1 : RCA_GEN_NBIT4_97 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1475);
   mux : MUX21_GENERIC_NBIT4_49 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_48 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_48;

architecture SYN_STRUCTURAL of carry_select_block_n4_48 is

   component MUX21_GENERIC_NBIT4_48
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_95
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_96
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1476, 
      n_1477 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_96 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1476);
   RCA1 : RCA_GEN_NBIT4_95 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1477);
   mux : MUX21_GENERIC_NBIT4_48 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_47 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_47;

architecture SYN_STRUCTURAL of carry_select_block_n4_47 is

   component MUX21_GENERIC_NBIT4_47
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_93
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_94
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1478, 
      n_1479 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_94 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1478);
   RCA1 : RCA_GEN_NBIT4_93 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1479);
   mux : MUX21_GENERIC_NBIT4_47 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_46 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_46;

architecture SYN_STRUCTURAL of carry_select_block_n4_46 is

   component MUX21_GENERIC_NBIT4_46
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_91
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_92
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1480, 
      n_1481 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_92 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1480);
   RCA1 : RCA_GEN_NBIT4_91 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1481);
   mux : MUX21_GENERIC_NBIT4_46 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_45 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_45;

architecture SYN_STRUCTURAL of carry_select_block_n4_45 is

   component MUX21_GENERIC_NBIT4_45
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_89
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_90
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1482, 
      n_1483 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_90 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1482);
   RCA1 : RCA_GEN_NBIT4_89 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1483);
   mux : MUX21_GENERIC_NBIT4_45 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_44 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_44;

architecture SYN_STRUCTURAL of carry_select_block_n4_44 is

   component MUX21_GENERIC_NBIT4_44
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_87
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_88
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1484, 
      n_1485 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_88 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1484);
   RCA1 : RCA_GEN_NBIT4_87 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1485);
   mux : MUX21_GENERIC_NBIT4_44 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_43 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_43;

architecture SYN_STRUCTURAL of carry_select_block_n4_43 is

   component MUX21_GENERIC_NBIT4_43
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_85
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_86
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1486, 
      n_1487 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_86 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1486);
   RCA1 : RCA_GEN_NBIT4_85 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1487);
   mux : MUX21_GENERIC_NBIT4_43 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_42 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_42;

architecture SYN_STRUCTURAL of carry_select_block_n4_42 is

   component MUX21_GENERIC_NBIT4_42
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_83
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_84
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1488, 
      n_1489 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_84 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1488);
   RCA1 : RCA_GEN_NBIT4_83 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1489);
   mux : MUX21_GENERIC_NBIT4_42 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_41 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_41;

architecture SYN_STRUCTURAL of carry_select_block_n4_41 is

   component MUX21_GENERIC_NBIT4_41
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_81
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_82
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1490, 
      n_1491 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_82 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1490);
   RCA1 : RCA_GEN_NBIT4_81 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1491);
   mux : MUX21_GENERIC_NBIT4_41 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_40 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_40;

architecture SYN_STRUCTURAL of carry_select_block_n4_40 is

   component MUX21_GENERIC_NBIT4_40
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_79
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_80
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1492, 
      n_1493 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_80 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1492);
   RCA1 : RCA_GEN_NBIT4_79 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1493);
   mux : MUX21_GENERIC_NBIT4_40 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_39 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_39;

architecture SYN_STRUCTURAL of carry_select_block_n4_39 is

   component MUX21_GENERIC_NBIT4_39
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_77
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_78
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1494, 
      n_1495 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_78 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1494);
   RCA1 : RCA_GEN_NBIT4_77 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1495);
   mux : MUX21_GENERIC_NBIT4_39 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_38 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_38;

architecture SYN_STRUCTURAL of carry_select_block_n4_38 is

   component MUX21_GENERIC_NBIT4_38
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_75
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_76
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1496, 
      n_1497 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_76 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1496);
   RCA1 : RCA_GEN_NBIT4_75 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1497);
   mux : MUX21_GENERIC_NBIT4_38 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_37 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_37;

architecture SYN_STRUCTURAL of carry_select_block_n4_37 is

   component MUX21_GENERIC_NBIT4_37
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_73
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_74
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1498, 
      n_1499 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_74 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1498);
   RCA1 : RCA_GEN_NBIT4_73 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1499);
   mux : MUX21_GENERIC_NBIT4_37 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_36 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_36;

architecture SYN_STRUCTURAL of carry_select_block_n4_36 is

   component MUX21_GENERIC_NBIT4_36
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_71
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_72
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1500, 
      n_1501 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_72 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1500);
   RCA1 : RCA_GEN_NBIT4_71 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1501);
   mux : MUX21_GENERIC_NBIT4_36 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_35 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_35;

architecture SYN_STRUCTURAL of carry_select_block_n4_35 is

   component MUX21_GENERIC_NBIT4_35
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_69
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_70
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1502, 
      n_1503 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_70 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1502);
   RCA1 : RCA_GEN_NBIT4_69 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1503);
   mux : MUX21_GENERIC_NBIT4_35 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_34 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_34;

architecture SYN_STRUCTURAL of carry_select_block_n4_34 is

   component MUX21_GENERIC_NBIT4_34
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_67
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_68
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1504, 
      n_1505 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_68 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1504);
   RCA1 : RCA_GEN_NBIT4_67 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1505);
   mux : MUX21_GENERIC_NBIT4_34 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_33 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_33;

architecture SYN_STRUCTURAL of carry_select_block_n4_33 is

   component MUX21_GENERIC_NBIT4_33
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_65
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_66
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1506, 
      n_1507 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_66 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1506);
   RCA1 : RCA_GEN_NBIT4_65 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1507);
   mux : MUX21_GENERIC_NBIT4_33 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_32 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_32;

architecture SYN_STRUCTURAL_architecture of carry_select_block_n4_32 is

   component MUX21_GENERIC_NBIT4_32
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_63
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_64
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1508, 
      n_1509 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_64 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1508);
   RCA1 : RCA_GEN_NBIT4_63 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1509);
   mux : MUX21_GENERIC_NBIT4_32 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_31 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_31;

architecture SYN_STRUCTURAL_architecture2 of carry_select_block_n4_31 is

   component MUX21_GENERIC_NBIT4_31
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_61
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_62
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1510, 
      n_1511 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_62 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1510);
   RCA1 : RCA_GEN_NBIT4_61 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1511);
   mux : MUX21_GENERIC_NBIT4_31 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_30 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_30;

architecture SYN_STRUCTURAL_architecture3 of carry_select_block_n4_30 is

   component MUX21_GENERIC_NBIT4_30
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_59
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_60
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1512, 
      n_1513 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_60 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1512);
   RCA1 : RCA_GEN_NBIT4_59 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1513);
   mux : MUX21_GENERIC_NBIT4_30 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_29 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_29;

architecture SYN_STRUCTURAL_architecture4 of carry_select_block_n4_29 is

   component MUX21_GENERIC_NBIT4_29
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_57
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_58
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1514, 
      n_1515 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_58 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1514);
   RCA1 : RCA_GEN_NBIT4_57 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1515);
   mux : MUX21_GENERIC_NBIT4_29 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_28 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_28;

architecture SYN_STRUCTURAL_architecture5 of carry_select_block_n4_28 is

   component MUX21_GENERIC_NBIT4_28
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_55
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_56
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1516, 
      n_1517 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_56 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1516);
   RCA1 : RCA_GEN_NBIT4_55 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1517);
   mux : MUX21_GENERIC_NBIT4_28 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL_architecture5;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_27 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_27;

architecture SYN_STRUCTURAL_architecture6 of carry_select_block_n4_27 is

   component MUX21_GENERIC_NBIT4_27
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_53
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_54
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1518, 
      n_1519 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_54 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1518);
   RCA1 : RCA_GEN_NBIT4_53 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1519);
   mux : MUX21_GENERIC_NBIT4_27 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL_architecture6;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_26 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_26;

architecture SYN_STRUCTURAL_architecture7 of carry_select_block_n4_26 is

   component MUX21_GENERIC_NBIT4_26
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_51
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_52
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1520, 
      n_1521 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_52 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1520);
   RCA1 : RCA_GEN_NBIT4_51 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1521);
   mux : MUX21_GENERIC_NBIT4_26 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL_architecture7;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_25 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_25;

architecture SYN_STRUCTURAL_architecture8 of carry_select_block_n4_25 is

   component MUX21_GENERIC_NBIT4_25
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_49
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_50
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1522, 
      n_1523 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_50 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1522);
   RCA1 : RCA_GEN_NBIT4_49 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1523);
   mux : MUX21_GENERIC_NBIT4_25 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL_architecture8;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_24 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_24;

architecture SYN_STRUCTURAL_architecture9 of carry_select_block_n4_24 is

   component MUX21_GENERIC_NBIT4_24
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_47
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_48
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1524, 
      n_1525 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_48 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1524);
   RCA1 : RCA_GEN_NBIT4_47 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1525);
   mux : MUX21_GENERIC_NBIT4_24 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL_architecture9;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_23 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_23;

architecture SYN_STRUCTURAL_architecture10 of carry_select_block_n4_23 is

   component MUX21_GENERIC_NBIT4_23
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_45
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_46
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1526, 
      n_1527 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_46 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1526);
   RCA1 : RCA_GEN_NBIT4_45 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1527);
   mux : MUX21_GENERIC_NBIT4_23 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL_architecture10;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_22 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_22;

architecture SYN_STRUCTURAL_architecture11 of carry_select_block_n4_22 is

   component MUX21_GENERIC_NBIT4_22
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_43
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_44
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1528, 
      n_1529 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_44 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1528);
   RCA1 : RCA_GEN_NBIT4_43 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1529);
   mux : MUX21_GENERIC_NBIT4_22 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL_architecture11;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_21 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_21;

architecture SYN_STRUCTURAL_architecture12 of carry_select_block_n4_21 is

   component MUX21_GENERIC_NBIT4_21
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_41
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_42
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1530, 
      n_1531 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_42 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1530);
   RCA1 : RCA_GEN_NBIT4_41 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1531);
   mux : MUX21_GENERIC_NBIT4_21 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL_architecture12;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_20 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_20;

architecture SYN_STRUCTURAL_architecture13 of carry_select_block_n4_20 is

   component MUX21_GENERIC_NBIT4_20
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_39
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_40
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1532, 
      n_1533 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_40 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1532);
   RCA1 : RCA_GEN_NBIT4_39 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1533);
   mux : MUX21_GENERIC_NBIT4_20 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL_architecture13;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_19 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_19;

architecture SYN_STRUCTURAL_architecture14 of carry_select_block_n4_19 is

   component MUX21_GENERIC_NBIT4_19
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_37
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_38
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1534, 
      n_1535 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_38 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1534);
   RCA1 : RCA_GEN_NBIT4_37 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1535);
   mux : MUX21_GENERIC_NBIT4_19 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL_architecture14;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_18 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_18;

architecture SYN_STRUCTURAL_architecture15 of carry_select_block_n4_18 is

   component MUX21_GENERIC_NBIT4_18
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_35
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_36
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1536, 
      n_1537 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_36 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1536);
   RCA1 : RCA_GEN_NBIT4_35 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1537);
   mux : MUX21_GENERIC_NBIT4_18 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL_architecture15;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_17 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_17;

architecture SYN_STRUCTURAL_architecture16 of carry_select_block_n4_17 is

   component MUX21_GENERIC_NBIT4_17
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_33
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_34
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1538, 
      n_1539 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_34 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1538);
   RCA1 : RCA_GEN_NBIT4_33 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1539);
   mux : MUX21_GENERIC_NBIT4_17 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL_architecture16;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_16 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_16;

architecture SYN_STRUCTURAL_architecture of carry_select_block_n4_16 is

   component MUX21_GENERIC_NBIT4_16
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_31
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_32
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1540, 
      n_1541 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_32 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1540);
   RCA1 : RCA_GEN_NBIT4_31 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1541);
   mux : MUX21_GENERIC_NBIT4_16 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_15 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_15;

architecture SYN_STRUCTURAL_architecture2 of carry_select_block_n4_15 is

   component MUX21_GENERIC_NBIT4_15
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_29
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_30
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1542, 
      n_1543 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_30 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1542);
   RCA1 : RCA_GEN_NBIT4_29 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1543);
   mux : MUX21_GENERIC_NBIT4_15 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_14 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_14;

architecture SYN_STRUCTURAL_architecture3 of carry_select_block_n4_14 is

   component MUX21_GENERIC_NBIT4_14
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_27
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_28
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1544, 
      n_1545 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_28 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1544);
   RCA1 : RCA_GEN_NBIT4_27 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1545);
   mux : MUX21_GENERIC_NBIT4_14 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_13 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_13;

architecture SYN_STRUCTURAL_architecture4 of carry_select_block_n4_13 is

   component MUX21_GENERIC_NBIT4_13
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_25
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_26
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1546, 
      n_1547 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_26 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1546);
   RCA1 : RCA_GEN_NBIT4_25 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1547);
   mux : MUX21_GENERIC_NBIT4_13 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_12 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_12;

architecture SYN_STRUCTURAL_architecture5 of carry_select_block_n4_12 is

   component MUX21_GENERIC_NBIT4_12
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_23
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_24
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1548, 
      n_1549 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_24 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1548);
   RCA1 : RCA_GEN_NBIT4_23 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1549);
   mux : MUX21_GENERIC_NBIT4_12 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL_architecture5;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_11 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_11;

architecture SYN_STRUCTURAL_architecture6 of carry_select_block_n4_11 is

   component MUX21_GENERIC_NBIT4_11
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_21
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_22
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1550, 
      n_1551 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_22 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1550);
   RCA1 : RCA_GEN_NBIT4_21 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1551);
   mux : MUX21_GENERIC_NBIT4_11 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL_architecture6;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_10 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_10;

architecture SYN_STRUCTURAL_architecture7 of carry_select_block_n4_10 is

   component MUX21_GENERIC_NBIT4_10
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_19
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_20
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1552, 
      n_1553 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_20 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1552);
   RCA1 : RCA_GEN_NBIT4_19 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1553);
   mux : MUX21_GENERIC_NBIT4_10 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL_architecture7;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_9 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_9;

architecture SYN_STRUCTURAL_architecture8 of carry_select_block_n4_9 is

   component MUX21_GENERIC_NBIT4_9
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_17
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_18
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1554, 
      n_1555 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_18 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1554);
   RCA1 : RCA_GEN_NBIT4_17 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1555);
   mux : MUX21_GENERIC_NBIT4_9 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL_architecture8;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_8 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_8;

architecture SYN_STRUCTURAL_architecture9 of carry_select_block_n4_8 is

   component MUX21_GENERIC_NBIT4_8
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_15
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_16
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1556, 
      n_1557 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_16 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1556);
   RCA1 : RCA_GEN_NBIT4_15 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1557);
   mux : MUX21_GENERIC_NBIT4_8 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL_architecture9;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_7;

architecture SYN_STRUCTURAL_architecture10 of carry_select_block_n4_7 is

   component MUX21_GENERIC_NBIT4_7
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_13
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_14
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1558, 
      n_1559 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_14 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1558);
   RCA1 : RCA_GEN_NBIT4_13 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1559);
   mux : MUX21_GENERIC_NBIT4_7 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL_architecture10;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_6;

architecture SYN_STRUCTURAL_architecture11 of carry_select_block_n4_6 is

   component MUX21_GENERIC_NBIT4_6
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_11
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_12
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1560, 
      n_1561 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_12 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1560);
   RCA1 : RCA_GEN_NBIT4_11 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1561);
   mux : MUX21_GENERIC_NBIT4_6 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL_architecture11;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_5;

architecture SYN_STRUCTURAL_architecture12 of carry_select_block_n4_5 is

   component MUX21_GENERIC_NBIT4_5
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_9
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_10
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1562, 
      n_1563 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_10 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1562);
   RCA1 : RCA_GEN_NBIT4_9 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1563);
   mux : MUX21_GENERIC_NBIT4_5 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL_architecture12;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_4;

architecture SYN_STRUCTURAL_architecture13 of carry_select_block_n4_4 is

   component MUX21_GENERIC_NBIT4_4
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_7
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_8
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1564, 
      n_1565 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_8 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1564);
   RCA1 : RCA_GEN_NBIT4_7 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1565);
   mux : MUX21_GENERIC_NBIT4_4 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL_architecture13;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_3;

architecture SYN_STRUCTURAL_architecture14 of carry_select_block_n4_3 is

   component MUX21_GENERIC_NBIT4_3
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_5
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_6
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1566, 
      n_1567 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_6 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1566);
   RCA1 : RCA_GEN_NBIT4_5 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1567);
   mux : MUX21_GENERIC_NBIT4_3 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL_architecture14;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_2;

architecture SYN_STRUCTURAL_architecture15 of carry_select_block_n4_2 is

   component MUX21_GENERIC_NBIT4_2
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_3
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_4
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1568, 
      n_1569 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_4 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1568);
   RCA1 : RCA_GEN_NBIT4_3 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1569);
   mux : MUX21_GENERIC_NBIT4_2 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL_architecture15;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_1;

architecture SYN_STRUCTURAL_architecture16 of carry_select_block_n4_1 is

   component MUX21_GENERIC_NBIT4_1
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_1
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_2
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1570, 
      n_1571 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_2 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1570);
   RCA1 : RCA_GEN_NBIT4_1 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1571);
   mux : MUX21_GENERIC_NBIT4_1 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL_architecture16;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_68 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_68;

architecture SYN_behavioral of G_BLOCK_68 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_67 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_67;

architecture SYN_behavioral of G_BLOCK_67 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_66 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_66;

architecture SYN_behavioral of G_BLOCK_66 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_65 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_65;

architecture SYN_behavioral of G_BLOCK_65 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_64 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_64;

architecture SYN_behavioral of G_BLOCK_64 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_63 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_63;

architecture SYN_behavioral of G_BLOCK_63 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_62 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_62;

architecture SYN_behavioral of G_BLOCK_62 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_61 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_61;

architecture SYN_behavioral of G_BLOCK_61 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_60 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_60;

architecture SYN_behavioral of G_BLOCK_60 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_59 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_59;

architecture SYN_behavioral of G_BLOCK_59 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_58 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_58;

architecture SYN_behavioral of G_BLOCK_58 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_57 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_57;

architecture SYN_behavioral of G_BLOCK_57 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_56 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_56;

architecture SYN_behavioral of G_BLOCK_56 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_55 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_55;

architecture SYN_behavioral of G_BLOCK_55 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_54 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_54;

architecture SYN_behavioral of G_BLOCK_54 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_53 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_53;

architecture SYN_behavioral of G_BLOCK_53 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_52 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_52;

architecture SYN_behavioral of G_BLOCK_52 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_51 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_51;

architecture SYN_behavioral of G_BLOCK_51 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_50 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_50;

architecture SYN_behavioral of G_BLOCK_50 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_49 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_49;

architecture SYN_behavioral of G_BLOCK_49 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_48 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_48;

architecture SYN_behavioral of G_BLOCK_48 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_47 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_47;

architecture SYN_behavioral of G_BLOCK_47 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_46 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_46;

architecture SYN_behavioral of G_BLOCK_46 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_45 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_45;

architecture SYN_behavioral of G_BLOCK_45 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_44 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_44;

architecture SYN_behavioral of G_BLOCK_44 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_43 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_43;

architecture SYN_behavioral of G_BLOCK_43 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_42 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_42;

architecture SYN_behavioral of G_BLOCK_42 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_41 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_41;

architecture SYN_behavioral of G_BLOCK_41 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_40 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_40;

architecture SYN_behavioral of G_BLOCK_40 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_39 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_39;

architecture SYN_behavioral of G_BLOCK_39 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_38 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_38;

architecture SYN_behavioral of G_BLOCK_38 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_37 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_37;

architecture SYN_behavioral of G_BLOCK_37 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_36 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_36;

architecture SYN_behavioral of G_BLOCK_36 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_35 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_35;

architecture SYN_behavioral of G_BLOCK_35 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_34 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_34;

architecture SYN_behavioral of G_BLOCK_34 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_33 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_33;

architecture SYN_behavioral_architecture of G_BLOCK_33 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_32 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_32;

architecture SYN_behavioral_architecture2 of G_BLOCK_32 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_31 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_31;

architecture SYN_behavioral_architecture3 of G_BLOCK_31 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_30 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_30;

architecture SYN_behavioral_architecture4 of G_BLOCK_30 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_29 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_29;

architecture SYN_behavioral_architecture5 of G_BLOCK_29 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral_architecture5;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_28 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_28;

architecture SYN_behavioral_architecture6 of G_BLOCK_28 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral_architecture6;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_27 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_27;

architecture SYN_behavioral_architecture7 of G_BLOCK_27 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral_architecture7;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_26 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_26;

architecture SYN_behavioral_architecture8 of G_BLOCK_26 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral_architecture8;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_25 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_25;

architecture SYN_behavioral_architecture9 of G_BLOCK_25 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral_architecture9;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_24 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_24;

architecture SYN_behavioral_architecture10 of G_BLOCK_24 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral_architecture10;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_23 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_23;

architecture SYN_behavioral_architecture11 of G_BLOCK_23 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral_architecture11;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_22 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_22;

architecture SYN_behavioral_architecture12 of G_BLOCK_22 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral_architecture12;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_21 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_21;

architecture SYN_behavioral_architecture13 of G_BLOCK_21 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral_architecture13;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_20 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_20;

architecture SYN_behavioral_architecture14 of G_BLOCK_20 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral_architecture14;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_19 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_19;

architecture SYN_behavioral_architecture15 of G_BLOCK_19 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral_architecture15;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_18 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_18;

architecture SYN_behavioral_architecture16 of G_BLOCK_18 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral_architecture16;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_17 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_17;

architecture SYN_behavioral of G_BLOCK_17 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_16 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_16;

architecture SYN_behavioral_architecture of G_BLOCK_16 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_15 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_15;

architecture SYN_behavioral_architecture2 of G_BLOCK_15 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_14 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_14;

architecture SYN_behavioral_architecture3 of G_BLOCK_14 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_13 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_13;

architecture SYN_behavioral_architecture4 of G_BLOCK_13 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_12 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_12;

architecture SYN_behavioral_architecture5 of G_BLOCK_12 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral_architecture5;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_11 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_11;

architecture SYN_behavioral_architecture6 of G_BLOCK_11 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral_architecture6;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_10 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_10;

architecture SYN_behavioral_architecture7 of G_BLOCK_10 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral_architecture7;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_9 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_9;

architecture SYN_behavioral_architecture8 of G_BLOCK_9 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral_architecture8;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_8 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_8;

architecture SYN_behavioral_architecture9 of G_BLOCK_8 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral_architecture9;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_7 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_7;

architecture SYN_behavioral_architecture10 of G_BLOCK_7 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral_architecture10;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_6 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_6;

architecture SYN_behavioral_architecture11 of G_BLOCK_6 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral_architecture11;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_5 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_5;

architecture SYN_behavioral_architecture12 of G_BLOCK_5 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral_architecture12;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_4 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_4;

architecture SYN_behavioral_architecture13 of G_BLOCK_4 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral_architecture13;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_3 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_3;

architecture SYN_behavioral_architecture14 of G_BLOCK_3 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral_architecture14;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_2 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_2;

architecture SYN_behavioral_architecture15 of G_BLOCK_2 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral_architecture15;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_1 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_1;

architecture SYN_behavioral_architecture16 of G_BLOCK_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n3);

end SYN_behavioral_architecture16;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_242 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_242;

architecture SYN_behavioral of PG_BLOCK_242 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_241 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_241;

architecture SYN_behavioral of PG_BLOCK_241 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U2 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U3 : INV_X1 port map( A => n3, ZN => PG_G);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_240 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_240;

architecture SYN_behavioral of PG_BLOCK_240 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_239 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_239;

architecture SYN_behavioral of PG_BLOCK_239 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_238 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_238;

architecture SYN_behavioral of PG_BLOCK_238 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_237 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_237;

architecture SYN_behavioral of PG_BLOCK_237 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_236 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_236;

architecture SYN_behavioral of PG_BLOCK_236 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_235 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_235;

architecture SYN_behavioral of PG_BLOCK_235 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_234 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_234;

architecture SYN_behavioral of PG_BLOCK_234 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_233 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_233;

architecture SYN_behavioral of PG_BLOCK_233 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_232 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_232;

architecture SYN_behavioral of PG_BLOCK_232 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_231 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_231;

architecture SYN_behavioral of PG_BLOCK_231 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_230 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_230;

architecture SYN_behavioral of PG_BLOCK_230 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_229 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_229;

architecture SYN_behavioral of PG_BLOCK_229 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_228 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_228;

architecture SYN_behavioral of PG_BLOCK_228 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_227 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_227;

architecture SYN_behavioral of PG_BLOCK_227 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_226 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_226;

architecture SYN_behavioral of PG_BLOCK_226 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_225 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_225;

architecture SYN_behavioral of PG_BLOCK_225 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_224 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_224;

architecture SYN_behavioral of PG_BLOCK_224 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_223 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_223;

architecture SYN_behavioral of PG_BLOCK_223 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_222 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_222;

architecture SYN_behavioral of PG_BLOCK_222 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_221 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_221;

architecture SYN_behavioral of PG_BLOCK_221 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_220 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_220;

architecture SYN_behavioral of PG_BLOCK_220 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_219 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_219;

architecture SYN_behavioral of PG_BLOCK_219 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_218 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_218;

architecture SYN_behavioral of PG_BLOCK_218 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_217 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_217;

architecture SYN_behavioral of PG_BLOCK_217 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_216 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_216;

architecture SYN_behavioral of PG_BLOCK_216 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_215 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_215;

architecture SYN_behavioral of PG_BLOCK_215 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_214 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_214;

architecture SYN_behavioral of PG_BLOCK_214 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_213 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_213;

architecture SYN_behavioral of PG_BLOCK_213 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_212 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_212;

architecture SYN_behavioral of PG_BLOCK_212 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_211 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_211;

architecture SYN_behavioral of PG_BLOCK_211 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_210 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_210;

architecture SYN_behavioral of PG_BLOCK_210 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_209 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_209;

architecture SYN_behavioral of PG_BLOCK_209 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_208 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_208;

architecture SYN_behavioral of PG_BLOCK_208 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_207 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_207;

architecture SYN_behavioral of PG_BLOCK_207 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_206 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_206;

architecture SYN_behavioral of PG_BLOCK_206 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_205 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_205;

architecture SYN_behavioral of PG_BLOCK_205 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_204 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_204;

architecture SYN_behavioral of PG_BLOCK_204 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_203 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_203;

architecture SYN_behavioral of PG_BLOCK_203 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_202 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_202;

architecture SYN_behavioral of PG_BLOCK_202 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_201 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_201;

architecture SYN_behavioral of PG_BLOCK_201 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_200 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_200;

architecture SYN_behavioral of PG_BLOCK_200 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_199 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_199;

architecture SYN_behavioral of PG_BLOCK_199 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_198 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_198;

architecture SYN_behavioral of PG_BLOCK_198 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_197 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_197;

architecture SYN_behavioral of PG_BLOCK_197 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_196 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_196;

architecture SYN_behavioral of PG_BLOCK_196 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_195 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_195;

architecture SYN_behavioral of PG_BLOCK_195 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_194 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_194;

architecture SYN_behavioral of PG_BLOCK_194 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_193 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_193;

architecture SYN_behavioral of PG_BLOCK_193 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_192 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_192;

architecture SYN_behavioral of PG_BLOCK_192 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_191 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_191;

architecture SYN_behavioral of PG_BLOCK_191 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_190 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_190;

architecture SYN_behavioral of PG_BLOCK_190 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_189 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_189;

architecture SYN_behavioral of PG_BLOCK_189 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_188 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_188;

architecture SYN_behavioral of PG_BLOCK_188 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_187 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_187;

architecture SYN_behavioral of PG_BLOCK_187 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_186 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_186;

architecture SYN_behavioral of PG_BLOCK_186 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_185 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_185;

architecture SYN_behavioral of PG_BLOCK_185 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_184 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_184;

architecture SYN_behavioral of PG_BLOCK_184 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_183 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_183;

architecture SYN_behavioral of PG_BLOCK_183 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_182 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_182;

architecture SYN_behavioral of PG_BLOCK_182 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_181 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_181;

architecture SYN_behavioral of PG_BLOCK_181 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_180 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_180;

architecture SYN_behavioral of PG_BLOCK_180 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_179 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_179;

architecture SYN_behavioral of PG_BLOCK_179 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_178 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_178;

architecture SYN_behavioral of PG_BLOCK_178 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_177 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_177;

architecture SYN_behavioral of PG_BLOCK_177 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_176 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_176;

architecture SYN_behavioral of PG_BLOCK_176 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_175 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_175;

architecture SYN_behavioral of PG_BLOCK_175 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_174 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_174;

architecture SYN_behavioral of PG_BLOCK_174 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_173 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_173;

architecture SYN_behavioral of PG_BLOCK_173 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_172 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_172;

architecture SYN_behavioral of PG_BLOCK_172 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_171 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_171;

architecture SYN_behavioral of PG_BLOCK_171 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_170 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_170;

architecture SYN_behavioral of PG_BLOCK_170 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_169 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_169;

architecture SYN_behavioral of PG_BLOCK_169 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_168 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_168;

architecture SYN_behavioral of PG_BLOCK_168 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_167 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_167;

architecture SYN_behavioral of PG_BLOCK_167 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_166 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_166;

architecture SYN_behavioral of PG_BLOCK_166 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_165 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_165;

architecture SYN_behavioral of PG_BLOCK_165 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_164 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_164;

architecture SYN_behavioral of PG_BLOCK_164 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_163 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_163;

architecture SYN_behavioral of PG_BLOCK_163 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_162 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_162;

architecture SYN_behavioral of PG_BLOCK_162 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_161 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_161;

architecture SYN_behavioral of PG_BLOCK_161 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_160 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_160;

architecture SYN_behavioral of PG_BLOCK_160 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_159 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_159;

architecture SYN_behavioral of PG_BLOCK_159 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_158 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_158;

architecture SYN_behavioral of PG_BLOCK_158 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_157 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_157;

architecture SYN_behavioral of PG_BLOCK_157 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_156 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_156;

architecture SYN_behavioral of PG_BLOCK_156 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_155 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_155;

architecture SYN_behavioral of PG_BLOCK_155 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_154 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_154;

architecture SYN_behavioral of PG_BLOCK_154 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_153 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_153;

architecture SYN_behavioral of PG_BLOCK_153 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_152 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_152;

architecture SYN_behavioral of PG_BLOCK_152 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_151 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_151;

architecture SYN_behavioral of PG_BLOCK_151 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_150 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_150;

architecture SYN_behavioral of PG_BLOCK_150 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_149 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_149;

architecture SYN_behavioral of PG_BLOCK_149 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_148 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_148;

architecture SYN_behavioral of PG_BLOCK_148 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_147 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_147;

architecture SYN_behavioral of PG_BLOCK_147 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_146 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_146;

architecture SYN_behavioral of PG_BLOCK_146 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_145 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_145;

architecture SYN_behavioral of PG_BLOCK_145 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_144 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_144;

architecture SYN_behavioral of PG_BLOCK_144 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_143 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_143;

architecture SYN_behavioral of PG_BLOCK_143 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_142 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_142;

architecture SYN_behavioral of PG_BLOCK_142 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_141 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_141;

architecture SYN_behavioral of PG_BLOCK_141 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_140 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_140;

architecture SYN_behavioral of PG_BLOCK_140 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_139 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_139;

architecture SYN_behavioral of PG_BLOCK_139 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_138 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_138;

architecture SYN_behavioral of PG_BLOCK_138 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_137 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_137;

architecture SYN_behavioral of PG_BLOCK_137 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_136 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_136;

architecture SYN_behavioral of PG_BLOCK_136 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_135 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_135;

architecture SYN_behavioral of PG_BLOCK_135 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_134 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_134;

architecture SYN_behavioral of PG_BLOCK_134 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_133 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_133;

architecture SYN_behavioral of PG_BLOCK_133 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_132 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_132;

architecture SYN_behavioral of PG_BLOCK_132 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_131 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_131;

architecture SYN_behavioral of PG_BLOCK_131 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_130 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_130;

architecture SYN_behavioral of PG_BLOCK_130 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_129 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_129;

architecture SYN_behavioral of PG_BLOCK_129 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_128 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_128;

architecture SYN_behavioral of PG_BLOCK_128 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_127 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_127;

architecture SYN_behavioral of PG_BLOCK_127 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_126 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_126;

architecture SYN_behavioral_architecture17 of PG_BLOCK_126 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture17;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_125 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_125;

architecture SYN_behavioral_architecture18 of PG_BLOCK_125 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture18;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_124 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_124;

architecture SYN_behavioral_architecture19 of PG_BLOCK_124 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture19;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_123 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_123;

architecture SYN_behavioral_architecture20 of PG_BLOCK_123 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture20;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_122 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_122;

architecture SYN_behavioral_architecture21 of PG_BLOCK_122 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral_architecture21;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_121 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_121;

architecture SYN_behavioral_architecture22 of PG_BLOCK_121 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral_architecture22;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_120 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_120;

architecture SYN_behavioral_architecture23 of PG_BLOCK_120 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture23;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_119 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_119;

architecture SYN_behavioral_architecture24 of PG_BLOCK_119 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture24;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_118 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_118;

architecture SYN_behavioral_architecture25 of PG_BLOCK_118 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture25;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_117 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_117;

architecture SYN_behavioral_architecture26 of PG_BLOCK_117 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture26;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_116 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_116;

architecture SYN_behavioral_architecture27 of PG_BLOCK_116 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture27;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_115 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_115;

architecture SYN_behavioral_architecture28 of PG_BLOCK_115 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture28;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_114 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_114;

architecture SYN_behavioral_architecture29 of PG_BLOCK_114 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral_architecture29;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_113 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_113;

architecture SYN_behavioral_architecture30 of PG_BLOCK_113 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral_architecture30;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_112 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_112;

architecture SYN_behavioral_architecture31 of PG_BLOCK_112 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture31;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_111 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_111;

architecture SYN_behavioral_architecture32 of PG_BLOCK_111 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture32;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_110 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_110;

architecture SYN_behavioral_architecture33 of PG_BLOCK_110 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture33;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_109 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_109;

architecture SYN_behavioral_architecture34 of PG_BLOCK_109 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture34;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_108 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_108;

architecture SYN_behavioral_architecture35 of PG_BLOCK_108 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture35;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_107 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_107;

architecture SYN_behavioral_architecture36 of PG_BLOCK_107 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture36;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_106 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_106;

architecture SYN_behavioral_architecture37 of PG_BLOCK_106 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral_architecture37;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_105 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_105;

architecture SYN_behavioral_architecture38 of PG_BLOCK_105 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral_architecture38;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_104 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_104;

architecture SYN_behavioral_architecture39 of PG_BLOCK_104 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture39;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_103 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_103;

architecture SYN_behavioral_architecture40 of PG_BLOCK_103 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture40;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_102 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_102;

architecture SYN_behavioral_architecture41 of PG_BLOCK_102 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture41;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_101 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_101;

architecture SYN_behavioral_architecture42 of PG_BLOCK_101 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral_architecture42;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_100 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_100;

architecture SYN_behavioral_architecture43 of PG_BLOCK_100 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture43;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_99 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_99;

architecture SYN_behavioral_architecture44 of PG_BLOCK_99 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture44;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_98 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_98;

architecture SYN_behavioral_architecture45 of PG_BLOCK_98 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture45;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_97 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_97;

architecture SYN_behavioral_architecture46 of PG_BLOCK_97 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture46;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_96 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_96;

architecture SYN_behavioral_architecture47 of PG_BLOCK_96 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral_architecture47;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_95 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_95;

architecture SYN_behavioral_architecture48 of PG_BLOCK_95 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture48;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_94 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_94;

architecture SYN_behavioral_architecture49 of PG_BLOCK_94 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture49;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_93 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_93;

architecture SYN_behavioral_architecture50 of PG_BLOCK_93 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture50;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_92 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_92;

architecture SYN_behavioral_architecture51 of PG_BLOCK_92 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture51;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_91 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_91;

architecture SYN_behavioral_architecture52 of PG_BLOCK_91 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture52;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_90 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_90;

architecture SYN_behavioral_architecture53 of PG_BLOCK_90 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture53;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_89 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_89;

architecture SYN_behavioral_architecture54 of PG_BLOCK_89 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture54;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_88 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_88;

architecture SYN_behavioral_architecture55 of PG_BLOCK_88 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture55;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_87 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_87;

architecture SYN_behavioral_architecture56 of PG_BLOCK_87 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture56;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_86 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_86;

architecture SYN_behavioral_architecture57 of PG_BLOCK_86 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture57;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_85 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_85;

architecture SYN_behavioral_architecture58 of PG_BLOCK_85 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture58;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_84 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_84;

architecture SYN_behavioral_architecture59 of PG_BLOCK_84 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture59;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_83 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_83;

architecture SYN_behavioral_architecture60 of PG_BLOCK_83 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture60;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_82 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_82;

architecture SYN_behavioral_architecture61 of PG_BLOCK_82 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture61;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_81 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_81;

architecture SYN_behavioral_architecture62 of PG_BLOCK_81 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral_architecture62;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_80 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_80;

architecture SYN_behavioral_architecture63 of PG_BLOCK_80 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral_architecture63;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_79 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_79;

architecture SYN_behavioral_architecture64 of PG_BLOCK_79 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture64;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_78 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_78;

architecture SYN_behavioral_architecture65 of PG_BLOCK_78 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture65;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_77 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_77;

architecture SYN_behavioral_architecture66 of PG_BLOCK_77 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture66;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_76 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_76;

architecture SYN_behavioral_architecture67 of PG_BLOCK_76 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture67;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_75 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_75;

architecture SYN_behavioral_architecture68 of PG_BLOCK_75 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture68;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_74 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_74;

architecture SYN_behavioral_architecture69 of PG_BLOCK_74 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral_architecture69;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_73 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_73;

architecture SYN_behavioral_architecture70 of PG_BLOCK_73 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral_architecture70;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_72 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_72;

architecture SYN_behavioral_architecture71 of PG_BLOCK_72 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture71;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_71 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_71;

architecture SYN_behavioral_architecture72 of PG_BLOCK_71 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral_architecture72;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_70 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_70;

architecture SYN_behavioral_architecture73 of PG_BLOCK_70 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral_architecture73;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_69 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_69;

architecture SYN_behavioral_architecture74 of PG_BLOCK_69 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral_architecture74;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_68 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_68;

architecture SYN_behavioral_architecture75 of PG_BLOCK_68 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral_architecture75;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_67 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_67;

architecture SYN_behavioral_architecture76 of PG_BLOCK_67 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral_architecture76;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_66 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_66;

architecture SYN_behavioral_architecture77 of PG_BLOCK_66 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral_architecture77;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_65 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_65;

architecture SYN_behavioral_architecture78 of PG_BLOCK_65 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral_architecture78;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_64 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_64;

architecture SYN_behavioral_architecture79 of PG_BLOCK_64 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral_architecture79;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_63 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_63;

architecture SYN_behavioral_architecture17 of PG_BLOCK_63 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture17;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_62 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_62;

architecture SYN_behavioral_architecture18 of PG_BLOCK_62 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture18;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_61 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_61;

architecture SYN_behavioral_architecture19 of PG_BLOCK_61 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture19;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_60 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_60;

architecture SYN_behavioral_architecture20 of PG_BLOCK_60 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture20;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_59 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_59;

architecture SYN_behavioral_architecture21 of PG_BLOCK_59 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral_architecture21;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_58 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_58;

architecture SYN_behavioral_architecture22 of PG_BLOCK_58 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral_architecture22;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_57 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_57;

architecture SYN_behavioral_architecture23 of PG_BLOCK_57 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture23;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_56 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_56;

architecture SYN_behavioral_architecture24 of PG_BLOCK_56 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture24;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_55 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_55;

architecture SYN_behavioral_architecture25 of PG_BLOCK_55 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture25;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_54 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_54;

architecture SYN_behavioral_architecture26 of PG_BLOCK_54 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture26;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_53 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_53;

architecture SYN_behavioral_architecture27 of PG_BLOCK_53 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture27;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_52 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_52;

architecture SYN_behavioral_architecture28 of PG_BLOCK_52 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture28;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_51 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_51;

architecture SYN_behavioral_architecture29 of PG_BLOCK_51 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral_architecture29;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_50 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_50;

architecture SYN_behavioral_architecture30 of PG_BLOCK_50 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral_architecture30;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_49 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_49;

architecture SYN_behavioral_architecture31 of PG_BLOCK_49 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture31;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_48 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_48;

architecture SYN_behavioral_architecture32 of PG_BLOCK_48 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture32;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_47 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_47;

architecture SYN_behavioral_architecture33 of PG_BLOCK_47 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture33;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_46 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_46;

architecture SYN_behavioral_architecture34 of PG_BLOCK_46 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture34;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_45 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_45;

architecture SYN_behavioral_architecture35 of PG_BLOCK_45 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture35;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_44 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_44;

architecture SYN_behavioral_architecture36 of PG_BLOCK_44 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture36;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_43 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_43;

architecture SYN_behavioral_architecture37 of PG_BLOCK_43 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral_architecture37;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_42 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_42;

architecture SYN_behavioral_architecture38 of PG_BLOCK_42 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral_architecture38;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_41 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_41;

architecture SYN_behavioral_architecture39 of PG_BLOCK_41 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture39;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_40 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_40;

architecture SYN_behavioral_architecture40 of PG_BLOCK_40 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture40;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_39 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_39;

architecture SYN_behavioral_architecture41 of PG_BLOCK_39 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture41;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_38 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_38;

architecture SYN_behavioral_architecture42 of PG_BLOCK_38 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral_architecture42;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_37 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_37;

architecture SYN_behavioral_architecture43 of PG_BLOCK_37 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture43;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_36 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_36;

architecture SYN_behavioral_architecture44 of PG_BLOCK_36 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture44;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_35 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_35;

architecture SYN_behavioral_architecture45 of PG_BLOCK_35 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture45;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_34 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_34;

architecture SYN_behavioral_architecture46 of PG_BLOCK_34 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture46;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_33 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_33;

architecture SYN_behavioral_architecture47 of PG_BLOCK_33 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral_architecture47;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_32 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_32;

architecture SYN_behavioral_architecture48 of PG_BLOCK_32 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture48;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_31 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_31;

architecture SYN_behavioral_architecture49 of PG_BLOCK_31 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture49;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_30 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_30;

architecture SYN_behavioral_architecture50 of PG_BLOCK_30 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture50;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_29 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_29;

architecture SYN_behavioral_architecture51 of PG_BLOCK_29 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture51;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_28 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_28;

architecture SYN_behavioral_architecture52 of PG_BLOCK_28 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture52;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_27 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_27;

architecture SYN_behavioral_architecture53 of PG_BLOCK_27 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture53;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_26 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_26;

architecture SYN_behavioral_architecture54 of PG_BLOCK_26 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture54;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_25 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_25;

architecture SYN_behavioral_architecture55 of PG_BLOCK_25 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture55;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_24 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_24;

architecture SYN_behavioral_architecture56 of PG_BLOCK_24 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture56;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_23 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_23;

architecture SYN_behavioral_architecture57 of PG_BLOCK_23 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture57;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_22 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_22;

architecture SYN_behavioral_architecture58 of PG_BLOCK_22 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture58;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_21 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_21;

architecture SYN_behavioral_architecture59 of PG_BLOCK_21 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture59;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_20 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_20;

architecture SYN_behavioral_architecture60 of PG_BLOCK_20 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture60;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_19 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_19;

architecture SYN_behavioral_architecture61 of PG_BLOCK_19 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture61;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_18 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_18;

architecture SYN_behavioral_architecture62 of PG_BLOCK_18 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral_architecture62;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_17 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_17;

architecture SYN_behavioral_architecture63 of PG_BLOCK_17 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral_architecture63;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_16 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_16;

architecture SYN_behavioral_architecture64 of PG_BLOCK_16 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral_architecture64;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_15 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_15;

architecture SYN_behavioral_architecture65 of PG_BLOCK_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture65;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_14 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_14;

architecture SYN_behavioral_architecture66 of PG_BLOCK_14 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture66;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_13 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_13;

architecture SYN_behavioral_architecture67 of PG_BLOCK_13 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture67;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_12 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_12;

architecture SYN_behavioral_architecture68 of PG_BLOCK_12 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture68;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_11 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_11;

architecture SYN_behavioral_architecture69 of PG_BLOCK_11 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral_architecture69;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_10 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_10;

architecture SYN_behavioral_architecture70 of PG_BLOCK_10 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral_architecture70;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_9 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_9;

architecture SYN_behavioral_architecture71 of PG_BLOCK_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);
   U3 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);

end SYN_behavioral_architecture71;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_8 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_8;

architecture SYN_behavioral_architecture72 of PG_BLOCK_8 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral_architecture72;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_7 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_7;

architecture SYN_behavioral_architecture73 of PG_BLOCK_7 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral_architecture73;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_6 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_6;

architecture SYN_behavioral_architecture74 of PG_BLOCK_6 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral_architecture74;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_5 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_5;

architecture SYN_behavioral_architecture75 of PG_BLOCK_5 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n3, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral_architecture75;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_4 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_4;

architecture SYN_behavioral_architecture76 of PG_BLOCK_4 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral_architecture76;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_3 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_3;

architecture SYN_behavioral_architecture77 of PG_BLOCK_3 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral_architecture77;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_2 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_2;

architecture SYN_behavioral_architecture78 of PG_BLOCK_2 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral_architecture78;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_1 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_1;

architecture SYN_behavioral_architecture79 of PG_BLOCK_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => PG_G);
   U2 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n3);

end SYN_behavioral_architecture79;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_250 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_250;

architecture SYN_behavioral of pg_net_250 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_249 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_249;

architecture SYN_behavioral of pg_net_249 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_248 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_248;

architecture SYN_behavioral of pg_net_248 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_247 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_247;

architecture SYN_behavioral of pg_net_247 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_246 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_246;

architecture SYN_behavioral of pg_net_246 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_245 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_245;

architecture SYN_behavioral of pg_net_245 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_244 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_244;

architecture SYN_behavioral of pg_net_244 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_243 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_243;

architecture SYN_behavioral of pg_net_243 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_242 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_242;

architecture SYN_behavioral of pg_net_242 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_241 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_241;

architecture SYN_behavioral of pg_net_241 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_240 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_240;

architecture SYN_behavioral of pg_net_240 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_239 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_239;

architecture SYN_behavioral of pg_net_239 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_238 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_238;

architecture SYN_behavioral of pg_net_238 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_237 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_237;

architecture SYN_behavioral of pg_net_237 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_236 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_236;

architecture SYN_behavioral of pg_net_236 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_235 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_235;

architecture SYN_behavioral of pg_net_235 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_234 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_234;

architecture SYN_behavioral of pg_net_234 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_233 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_233;

architecture SYN_behavioral of pg_net_233 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_232 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_232;

architecture SYN_behavioral of pg_net_232 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_231 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_231;

architecture SYN_behavioral of pg_net_231 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_230 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_230;

architecture SYN_behavioral of pg_net_230 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_229 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_229;

architecture SYN_behavioral of pg_net_229 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_228 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_228;

architecture SYN_behavioral of pg_net_228 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_227 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_227;

architecture SYN_behavioral of pg_net_227 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_226 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_226;

architecture SYN_behavioral of pg_net_226 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_225 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_225;

architecture SYN_behavioral of pg_net_225 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_224 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_224;

architecture SYN_behavioral of pg_net_224 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_223 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_223;

architecture SYN_behavioral of pg_net_223 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_222 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_222;

architecture SYN_behavioral of pg_net_222 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_221 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_221;

architecture SYN_behavioral of pg_net_221 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_220 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_220;

architecture SYN_behavioral of pg_net_220 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_219 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_219;

architecture SYN_behavioral of pg_net_219 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_218 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_218;

architecture SYN_behavioral of pg_net_218 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_217 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_217;

architecture SYN_behavioral of pg_net_217 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_216 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_216;

architecture SYN_behavioral of pg_net_216 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_215 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_215;

architecture SYN_behavioral of pg_net_215 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_214 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_214;

architecture SYN_behavioral of pg_net_214 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_213 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_213;

architecture SYN_behavioral of pg_net_213 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_212 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_212;

architecture SYN_behavioral of pg_net_212 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_211 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_211;

architecture SYN_behavioral of pg_net_211 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_210 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_210;

architecture SYN_behavioral of pg_net_210 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_209 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_209;

architecture SYN_behavioral of pg_net_209 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_208 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_208;

architecture SYN_behavioral of pg_net_208 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_207 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_207;

architecture SYN_behavioral of pg_net_207 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_206 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_206;

architecture SYN_behavioral of pg_net_206 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_205 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_205;

architecture SYN_behavioral of pg_net_205 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_204 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_204;

architecture SYN_behavioral of pg_net_204 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_203 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_203;

architecture SYN_behavioral of pg_net_203 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_202 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_202;

architecture SYN_behavioral of pg_net_202 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_201 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_201;

architecture SYN_behavioral of pg_net_201 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_200 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_200;

architecture SYN_behavioral of pg_net_200 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_199 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_199;

architecture SYN_behavioral of pg_net_199 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_198 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_198;

architecture SYN_behavioral of pg_net_198 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_197 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_197;

architecture SYN_behavioral of pg_net_197 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_196 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_196;

architecture SYN_behavioral of pg_net_196 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_195 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_195;

architecture SYN_behavioral of pg_net_195 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_194 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_194;

architecture SYN_behavioral of pg_net_194 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_193 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_193;

architecture SYN_behavioral of pg_net_193 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_192 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_192;

architecture SYN_behavioral of pg_net_192 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_191 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_191;

architecture SYN_behavioral of pg_net_191 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_190 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_190;

architecture SYN_behavioral of pg_net_190 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_189 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_189;

architecture SYN_behavioral of pg_net_189 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_188 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_188;

architecture SYN_behavioral of pg_net_188 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_187 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_187;

architecture SYN_behavioral of pg_net_187 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_186 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_186;

architecture SYN_behavioral of pg_net_186 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_185 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_185;

architecture SYN_behavioral of pg_net_185 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_184 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_184;

architecture SYN_behavioral of pg_net_184 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_183 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_183;

architecture SYN_behavioral of pg_net_183 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_182 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_182;

architecture SYN_behavioral of pg_net_182 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_181 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_181;

architecture SYN_behavioral of pg_net_181 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_180 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_180;

architecture SYN_behavioral of pg_net_180 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_179 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_179;

architecture SYN_behavioral of pg_net_179 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_178 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_178;

architecture SYN_behavioral of pg_net_178 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_177 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_177;

architecture SYN_behavioral of pg_net_177 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_176 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_176;

architecture SYN_behavioral of pg_net_176 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_175 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_175;

architecture SYN_behavioral of pg_net_175 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_174 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_174;

architecture SYN_behavioral of pg_net_174 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_173 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_173;

architecture SYN_behavioral of pg_net_173 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_172 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_172;

architecture SYN_behavioral of pg_net_172 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_171 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_171;

architecture SYN_behavioral of pg_net_171 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_170 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_170;

architecture SYN_behavioral of pg_net_170 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_169 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_169;

architecture SYN_behavioral of pg_net_169 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_168 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_168;

architecture SYN_behavioral of pg_net_168 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_167 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_167;

architecture SYN_behavioral of pg_net_167 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_166 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_166;

architecture SYN_behavioral of pg_net_166 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_165 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_165;

architecture SYN_behavioral of pg_net_165 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_164 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_164;

architecture SYN_behavioral of pg_net_164 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_163 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_163;

architecture SYN_behavioral of pg_net_163 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_162 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_162;

architecture SYN_behavioral of pg_net_162 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_161 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_161;

architecture SYN_behavioral of pg_net_161 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_160 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_160;

architecture SYN_behavioral of pg_net_160 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_159 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_159;

architecture SYN_behavioral of pg_net_159 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_158 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_158;

architecture SYN_behavioral of pg_net_158 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_157 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_157;

architecture SYN_behavioral of pg_net_157 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_156 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_156;

architecture SYN_behavioral of pg_net_156 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_155 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_155;

architecture SYN_behavioral of pg_net_155 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_154 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_154;

architecture SYN_behavioral of pg_net_154 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_153 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_153;

architecture SYN_behavioral of pg_net_153 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_152 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_152;

architecture SYN_behavioral of pg_net_152 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_151 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_151;

architecture SYN_behavioral of pg_net_151 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_150 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_150;

architecture SYN_behavioral of pg_net_150 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_149 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_149;

architecture SYN_behavioral of pg_net_149 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_148 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_148;

architecture SYN_behavioral of pg_net_148 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_147 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_147;

architecture SYN_behavioral of pg_net_147 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_146 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_146;

architecture SYN_behavioral of pg_net_146 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_145 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_145;

architecture SYN_behavioral of pg_net_145 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_144 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_144;

architecture SYN_behavioral of pg_net_144 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_143 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_143;

architecture SYN_behavioral of pg_net_143 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_142 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_142;

architecture SYN_behavioral of pg_net_142 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_141 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_141;

architecture SYN_behavioral of pg_net_141 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_140 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_140;

architecture SYN_behavioral of pg_net_140 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_139 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_139;

architecture SYN_behavioral of pg_net_139 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_138 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_138;

architecture SYN_behavioral of pg_net_138 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_137 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_137;

architecture SYN_behavioral of pg_net_137 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_136 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_136;

architecture SYN_behavioral of pg_net_136 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_135 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_135;

architecture SYN_behavioral of pg_net_135 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_134 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_134;

architecture SYN_behavioral of pg_net_134 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_133 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_133;

architecture SYN_behavioral of pg_net_133 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_132 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_132;

architecture SYN_behavioral of pg_net_132 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_131 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_131;

architecture SYN_behavioral of pg_net_131 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_130 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_130;

architecture SYN_behavioral of pg_net_130 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_129 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_129;

architecture SYN_behavioral of pg_net_129 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_128 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_128;

architecture SYN_behavioral of pg_net_128 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_127 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_127;

architecture SYN_behavioral of pg_net_127 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_126 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_126;

architecture SYN_behavioral_architecture80 of pg_net_126 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture80;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_125 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_125;

architecture SYN_behavioral_architecture81 of pg_net_125 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture81;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_124 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_124;

architecture SYN_behavioral_architecture82 of pg_net_124 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture82;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_123 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_123;

architecture SYN_behavioral_architecture83 of pg_net_123 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture83;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_122 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_122;

architecture SYN_behavioral_architecture84 of pg_net_122 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture84;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_121 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_121;

architecture SYN_behavioral_architecture85 of pg_net_121 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture85;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_120 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_120;

architecture SYN_behavioral_architecture86 of pg_net_120 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture86;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_119 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_119;

architecture SYN_behavioral_architecture87 of pg_net_119 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture87;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_118 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_118;

architecture SYN_behavioral_architecture88 of pg_net_118 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture88;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_117 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_117;

architecture SYN_behavioral_architecture89 of pg_net_117 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture89;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_116 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_116;

architecture SYN_behavioral_architecture90 of pg_net_116 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture90;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_115 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_115;

architecture SYN_behavioral_architecture91 of pg_net_115 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture91;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_114 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_114;

architecture SYN_behavioral_architecture92 of pg_net_114 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture92;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_113 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_113;

architecture SYN_behavioral_architecture93 of pg_net_113 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture93;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_112 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_112;

architecture SYN_behavioral_architecture94 of pg_net_112 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture94;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_111 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_111;

architecture SYN_behavioral_architecture95 of pg_net_111 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture95;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_110 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_110;

architecture SYN_behavioral_architecture96 of pg_net_110 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture96;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_109 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_109;

architecture SYN_behavioral_architecture97 of pg_net_109 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture97;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_108 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_108;

architecture SYN_behavioral_architecture98 of pg_net_108 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture98;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_107 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_107;

architecture SYN_behavioral_architecture99 of pg_net_107 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture99;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_106 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_106;

architecture SYN_behavioral_architecture100 of pg_net_106 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture100;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_105 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_105;

architecture SYN_behavioral_architecture101 of pg_net_105 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture101;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_104 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_104;

architecture SYN_behavioral_architecture102 of pg_net_104 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture102;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_103 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_103;

architecture SYN_behavioral_architecture103 of pg_net_103 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture103;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_102 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_102;

architecture SYN_behavioral_architecture104 of pg_net_102 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture104;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_101 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_101;

architecture SYN_behavioral_architecture105 of pg_net_101 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture105;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_100 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_100;

architecture SYN_behavioral_architecture106 of pg_net_100 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture106;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_99 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_99;

architecture SYN_behavioral_architecture107 of pg_net_99 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture107;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_98 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_98;

architecture SYN_behavioral_architecture108 of pg_net_98 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture108;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_97 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_97;

architecture SYN_behavioral_architecture109 of pg_net_97 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture109;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_96 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_96;

architecture SYN_behavioral_architecture110 of pg_net_96 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture110;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_95 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_95;

architecture SYN_behavioral_architecture111 of pg_net_95 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture111;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_94 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_94;

architecture SYN_behavioral_architecture112 of pg_net_94 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture112;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_93 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_93;

architecture SYN_behavioral_architecture113 of pg_net_93 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture113;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_92 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_92;

architecture SYN_behavioral_architecture114 of pg_net_92 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture114;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_91 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_91;

architecture SYN_behavioral_architecture115 of pg_net_91 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture115;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_90 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_90;

architecture SYN_behavioral_architecture116 of pg_net_90 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture116;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_89 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_89;

architecture SYN_behavioral_architecture117 of pg_net_89 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture117;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_88 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_88;

architecture SYN_behavioral_architecture118 of pg_net_88 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture118;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_87 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_87;

architecture SYN_behavioral_architecture119 of pg_net_87 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture119;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_86 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_86;

architecture SYN_behavioral_architecture120 of pg_net_86 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture120;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_85 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_85;

architecture SYN_behavioral_architecture121 of pg_net_85 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture121;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_84 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_84;

architecture SYN_behavioral_architecture122 of pg_net_84 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture122;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_83 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_83;

architecture SYN_behavioral_architecture123 of pg_net_83 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture123;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_82 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_82;

architecture SYN_behavioral_architecture124 of pg_net_82 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture124;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_81 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_81;

architecture SYN_behavioral_architecture125 of pg_net_81 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture125;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_80 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_80;

architecture SYN_behavioral_architecture126 of pg_net_80 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture126;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_79 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_79;

architecture SYN_behavioral_architecture127 of pg_net_79 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture127;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_78 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_78;

architecture SYN_behavioral_architecture128 of pg_net_78 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture128;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_77 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_77;

architecture SYN_behavioral_architecture129 of pg_net_77 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture129;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_76 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_76;

architecture SYN_behavioral_architecture130 of pg_net_76 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture130;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_75 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_75;

architecture SYN_behavioral_architecture131 of pg_net_75 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture131;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_74 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_74;

architecture SYN_behavioral_architecture132 of pg_net_74 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture132;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_73 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_73;

architecture SYN_behavioral_architecture133 of pg_net_73 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture133;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_72 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_72;

architecture SYN_behavioral_architecture134 of pg_net_72 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture134;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_71 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_71;

architecture SYN_behavioral_architecture135 of pg_net_71 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture135;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_70 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_70;

architecture SYN_behavioral_architecture136 of pg_net_70 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture136;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_69 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_69;

architecture SYN_behavioral_architecture137 of pg_net_69 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture137;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_68 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_68;

architecture SYN_behavioral_architecture138 of pg_net_68 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture138;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_67 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_67;

architecture SYN_behavioral_architecture139 of pg_net_67 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture139;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_66 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_66;

architecture SYN_behavioral_architecture140 of pg_net_66 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture140;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_65 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_65;

architecture SYN_behavioral_architecture141 of pg_net_65 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture141;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_64 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_64;

architecture SYN_behavioral_architecture142 of pg_net_64 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture142;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_63 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_63;

architecture SYN_behavioral_architecture80 of pg_net_63 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture80;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_62 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_62;

architecture SYN_behavioral_architecture81 of pg_net_62 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture81;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_61 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_61;

architecture SYN_behavioral_architecture82 of pg_net_61 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture82;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_60 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_60;

architecture SYN_behavioral_architecture83 of pg_net_60 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture83;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_59 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_59;

architecture SYN_behavioral_architecture84 of pg_net_59 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture84;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_58 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_58;

architecture SYN_behavioral_architecture85 of pg_net_58 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture85;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_57 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_57;

architecture SYN_behavioral_architecture86 of pg_net_57 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture86;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_56 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_56;

architecture SYN_behavioral_architecture87 of pg_net_56 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture87;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_55 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_55;

architecture SYN_behavioral_architecture88 of pg_net_55 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture88;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_54 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_54;

architecture SYN_behavioral_architecture89 of pg_net_54 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture89;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_53 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_53;

architecture SYN_behavioral_architecture90 of pg_net_53 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture90;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_52 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_52;

architecture SYN_behavioral_architecture91 of pg_net_52 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture91;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_51 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_51;

architecture SYN_behavioral_architecture92 of pg_net_51 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture92;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_50 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_50;

architecture SYN_behavioral_architecture93 of pg_net_50 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture93;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_49 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_49;

architecture SYN_behavioral_architecture94 of pg_net_49 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture94;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_48 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_48;

architecture SYN_behavioral_architecture95 of pg_net_48 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture95;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_47 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_47;

architecture SYN_behavioral_architecture96 of pg_net_47 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture96;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_46 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_46;

architecture SYN_behavioral_architecture97 of pg_net_46 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture97;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_45 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_45;

architecture SYN_behavioral_architecture98 of pg_net_45 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture98;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_44 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_44;

architecture SYN_behavioral_architecture99 of pg_net_44 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture99;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_43 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_43;

architecture SYN_behavioral_architecture100 of pg_net_43 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture100;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_42 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_42;

architecture SYN_behavioral_architecture101 of pg_net_42 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture101;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_41 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_41;

architecture SYN_behavioral_architecture102 of pg_net_41 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture102;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_40 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_40;

architecture SYN_behavioral_architecture103 of pg_net_40 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture103;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_39 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_39;

architecture SYN_behavioral_architecture104 of pg_net_39 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture104;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_38 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_38;

architecture SYN_behavioral_architecture105 of pg_net_38 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture105;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_37 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_37;

architecture SYN_behavioral_architecture106 of pg_net_37 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture106;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_36 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_36;

architecture SYN_behavioral_architecture107 of pg_net_36 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture107;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_35 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_35;

architecture SYN_behavioral_architecture108 of pg_net_35 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture108;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_34 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_34;

architecture SYN_behavioral_architecture109 of pg_net_34 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture109;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_33 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_33;

architecture SYN_behavioral_architecture110 of pg_net_33 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture110;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_32 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_32;

architecture SYN_behavioral_architecture111 of pg_net_32 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture111;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_31 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_31;

architecture SYN_behavioral_architecture112 of pg_net_31 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture112;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_30 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_30;

architecture SYN_behavioral_architecture113 of pg_net_30 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture113;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_29 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_29;

architecture SYN_behavioral_architecture114 of pg_net_29 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture114;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_28 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_28;

architecture SYN_behavioral_architecture115 of pg_net_28 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture115;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_27 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_27;

architecture SYN_behavioral_architecture116 of pg_net_27 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture116;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_26 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_26;

architecture SYN_behavioral_architecture117 of pg_net_26 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture117;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_25 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_25;

architecture SYN_behavioral_architecture118 of pg_net_25 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture118;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_24 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_24;

architecture SYN_behavioral_architecture119 of pg_net_24 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture119;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_23 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_23;

architecture SYN_behavioral_architecture120 of pg_net_23 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture120;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_22 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_22;

architecture SYN_behavioral_architecture121 of pg_net_22 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture121;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_21 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_21;

architecture SYN_behavioral_architecture122 of pg_net_21 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture122;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_20 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_20;

architecture SYN_behavioral_architecture123 of pg_net_20 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture123;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_19 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_19;

architecture SYN_behavioral_architecture124 of pg_net_19 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture124;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_18 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_18;

architecture SYN_behavioral_architecture125 of pg_net_18 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture125;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_17 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_17;

architecture SYN_behavioral_architecture126 of pg_net_17 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture126;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_16 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_16;

architecture SYN_behavioral_architecture127 of pg_net_16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture127;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_15 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_15;

architecture SYN_behavioral_architecture128 of pg_net_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture128;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_14 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_14;

architecture SYN_behavioral_architecture129 of pg_net_14 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture129;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_13 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_13;

architecture SYN_behavioral_architecture130 of pg_net_13 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture130;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_12 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_12;

architecture SYN_behavioral_architecture131 of pg_net_12 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture131;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_11 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_11;

architecture SYN_behavioral_architecture132 of pg_net_11 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture132;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_10 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_10;

architecture SYN_behavioral_architecture133 of pg_net_10 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture133;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_9 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_9;

architecture SYN_behavioral_architecture134 of pg_net_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture134;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_8 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_8;

architecture SYN_behavioral_architecture135 of pg_net_8 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture135;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_7 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_7;

architecture SYN_behavioral_architecture136 of pg_net_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture136;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_6 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_6;

architecture SYN_behavioral_architecture137 of pg_net_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture137;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_5 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_5;

architecture SYN_behavioral_architecture138 of pg_net_5 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture138;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_4 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_4;

architecture SYN_behavioral_architecture139 of pg_net_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture139;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_3 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_3;

architecture SYN_behavioral_architecture140 of pg_net_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture140;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_2 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_2;

architecture SYN_behavioral_architecture141 of pg_net_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture141;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_1 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_1;

architecture SYN_behavioral_architecture142 of pg_net_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral_architecture142;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX51_31 is

   port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0);  
         Y : out std_logic);

end MUX51_31;

architecture SYN_BEHAVIORAL of MUX51_31 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n9, n10, n11, n12 : std_logic;

begin
   
   U1 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S(0), B2 => B, ZN => n9);
   U2 : AOI22_X1 port map( A1 => C, A2 => n1, B1 => D, B2 => S(0), ZN => n10);
   U3 : INV_X1 port map( A => n12, ZN => Y);
   U4 : AOI22_X1 port map( A1 => n11, A2 => n3, B1 => S(2), B2 => E, ZN => n12)
                           ;
   U5 : OAI22_X1 port map( A1 => n10, A2 => n2, B1 => S(1), B2 => n9, ZN => n11
                           );
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);
   U8 : INV_X1 port map( A => S(2), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX51_30 is

   port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0);  
         Y : out std_logic);

end MUX51_30;

architecture SYN_BEHAVIORAL of MUX51_30 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n9, n10, n11, n12 : std_logic;

begin
   
   U1 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S(0), B2 => B, ZN => n9);
   U2 : AOI22_X1 port map( A1 => C, A2 => n1, B1 => D, B2 => S(0), ZN => n10);
   U3 : INV_X1 port map( A => n12, ZN => Y);
   U4 : AOI22_X1 port map( A1 => n11, A2 => n3, B1 => S(2), B2 => E, ZN => n12)
                           ;
   U5 : OAI22_X1 port map( A1 => n10, A2 => n2, B1 => S(1), B2 => n9, ZN => n11
                           );
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);
   U8 : INV_X1 port map( A => S(2), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX51_29 is

   port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0);  
         Y : out std_logic);

end MUX51_29;

architecture SYN_BEHAVIORAL of MUX51_29 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n9, n10, n11, n12 : std_logic;

begin
   
   U1 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S(0), B2 => B, ZN => n9);
   U2 : AOI22_X1 port map( A1 => C, A2 => n1, B1 => D, B2 => S(0), ZN => n10);
   U3 : INV_X1 port map( A => n12, ZN => Y);
   U4 : AOI22_X1 port map( A1 => n11, A2 => n3, B1 => S(2), B2 => E, ZN => n12)
                           ;
   U5 : OAI22_X1 port map( A1 => n10, A2 => n2, B1 => S(1), B2 => n9, ZN => n11
                           );
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);
   U8 : INV_X1 port map( A => S(2), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX51_28 is

   port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0);  
         Y : out std_logic);

end MUX51_28;

architecture SYN_BEHAVIORAL of MUX51_28 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n9, n10, n11, n12 : std_logic;

begin
   
   U1 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S(0), B2 => B, ZN => n9);
   U2 : AOI22_X1 port map( A1 => C, A2 => n1, B1 => D, B2 => S(0), ZN => n10);
   U3 : INV_X1 port map( A => n12, ZN => Y);
   U4 : AOI22_X1 port map( A1 => n11, A2 => n3, B1 => S(2), B2 => E, ZN => n12)
                           ;
   U5 : OAI22_X1 port map( A1 => n10, A2 => n2, B1 => S(1), B2 => n9, ZN => n11
                           );
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);
   U8 : INV_X1 port map( A => S(2), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX51_27 is

   port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0);  
         Y : out std_logic);

end MUX51_27;

architecture SYN_BEHAVIORAL of MUX51_27 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n9, n10, n11, n12 : std_logic;

begin
   
   U1 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S(0), B2 => B, ZN => n9);
   U2 : AOI22_X1 port map( A1 => C, A2 => n1, B1 => D, B2 => S(0), ZN => n10);
   U3 : INV_X1 port map( A => n12, ZN => Y);
   U4 : AOI22_X1 port map( A1 => n11, A2 => n3, B1 => S(2), B2 => E, ZN => n12)
                           ;
   U5 : OAI22_X1 port map( A1 => n10, A2 => n2, B1 => S(1), B2 => n9, ZN => n11
                           );
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);
   U8 : INV_X1 port map( A => S(2), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX51_26 is

   port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0);  
         Y : out std_logic);

end MUX51_26;

architecture SYN_BEHAVIORAL of MUX51_26 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n9, n10, n11, n12 : std_logic;

begin
   
   U1 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S(0), B2 => B, ZN => n9);
   U2 : AOI22_X1 port map( A1 => C, A2 => n1, B1 => D, B2 => S(0), ZN => n10);
   U3 : INV_X1 port map( A => n12, ZN => Y);
   U4 : AOI22_X1 port map( A1 => n11, A2 => n3, B1 => S(2), B2 => E, ZN => n12)
                           ;
   U5 : OAI22_X1 port map( A1 => n10, A2 => n2, B1 => S(1), B2 => n9, ZN => n11
                           );
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);
   U8 : INV_X1 port map( A => S(2), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX51_25 is

   port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0);  
         Y : out std_logic);

end MUX51_25;

architecture SYN_BEHAVIORAL of MUX51_25 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n9, n10, n11, n12 : std_logic;

begin
   
   U1 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S(0), B2 => B, ZN => n9);
   U2 : AOI22_X1 port map( A1 => C, A2 => n1, B1 => D, B2 => S(0), ZN => n10);
   U3 : INV_X1 port map( A => n12, ZN => Y);
   U4 : AOI22_X1 port map( A1 => n11, A2 => n3, B1 => S(2), B2 => E, ZN => n12)
                           ;
   U5 : OAI22_X1 port map( A1 => n10, A2 => n2, B1 => S(1), B2 => n9, ZN => n11
                           );
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);
   U8 : INV_X1 port map( A => S(2), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX51_24 is

   port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0);  
         Y : out std_logic);

end MUX51_24;

architecture SYN_BEHAVIORAL of MUX51_24 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n9, n10, n11, n12 : std_logic;

begin
   
   U1 : AOI22_X1 port map( A1 => C, A2 => n1, B1 => D, B2 => S(0), ZN => n10);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S(0), B2 => B, ZN => n9);
   U3 : INV_X1 port map( A => n12, ZN => Y);
   U4 : AOI22_X1 port map( A1 => n11, A2 => n3, B1 => S(2), B2 => E, ZN => n12)
                           ;
   U5 : OAI22_X1 port map( A1 => n10, A2 => n2, B1 => S(1), B2 => n9, ZN => n11
                           );
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);
   U8 : INV_X1 port map( A => S(2), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX51_23 is

   port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0);  
         Y : out std_logic);

end MUX51_23;

architecture SYN_BEHAVIORAL of MUX51_23 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n9, n10, n11, n12 : std_logic;

begin
   
   U1 : AOI22_X1 port map( A1 => C, A2 => n1, B1 => D, B2 => S(0), ZN => n10);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S(0), B2 => B, ZN => n9);
   U3 : INV_X1 port map( A => n12, ZN => Y);
   U4 : AOI22_X1 port map( A1 => n11, A2 => n3, B1 => S(2), B2 => E, ZN => n12)
                           ;
   U5 : OAI22_X1 port map( A1 => n10, A2 => n2, B1 => S(1), B2 => n9, ZN => n11
                           );
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);
   U8 : INV_X1 port map( A => S(2), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX51_22 is

   port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0);  
         Y : out std_logic);

end MUX51_22;

architecture SYN_BEHAVIORAL of MUX51_22 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n9, n10, n11, n12 : std_logic;

begin
   
   U1 : AOI22_X1 port map( A1 => C, A2 => n1, B1 => D, B2 => S(0), ZN => n10);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S(0), B2 => B, ZN => n9);
   U3 : INV_X1 port map( A => n12, ZN => Y);
   U4 : AOI22_X1 port map( A1 => n11, A2 => n3, B1 => S(2), B2 => E, ZN => n12)
                           ;
   U5 : OAI22_X1 port map( A1 => n10, A2 => n2, B1 => S(1), B2 => n9, ZN => n11
                           );
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);
   U8 : INV_X1 port map( A => S(2), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX51_21 is

   port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0);  
         Y : out std_logic);

end MUX51_21;

architecture SYN_BEHAVIORAL of MUX51_21 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n9, n10, n11, n12 : std_logic;

begin
   
   U1 : AOI22_X1 port map( A1 => C, A2 => n1, B1 => D, B2 => S(0), ZN => n10);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S(0), B2 => B, ZN => n9);
   U3 : INV_X1 port map( A => n12, ZN => Y);
   U4 : AOI22_X1 port map( A1 => n11, A2 => n3, B1 => S(2), B2 => E, ZN => n12)
                           ;
   U5 : OAI22_X1 port map( A1 => n10, A2 => n2, B1 => S(1), B2 => n9, ZN => n11
                           );
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);
   U8 : INV_X1 port map( A => S(2), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX51_20 is

   port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0);  
         Y : out std_logic);

end MUX51_20;

architecture SYN_BEHAVIORAL of MUX51_20 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n9, n10, n11, n12 : std_logic;

begin
   
   U1 : AOI22_X1 port map( A1 => C, A2 => n1, B1 => D, B2 => S(0), ZN => n10);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S(0), B2 => B, ZN => n9);
   U3 : INV_X1 port map( A => n12, ZN => Y);
   U4 : AOI22_X1 port map( A1 => n11, A2 => n3, B1 => S(2), B2 => E, ZN => n12)
                           ;
   U5 : OAI22_X1 port map( A1 => n10, A2 => n2, B1 => S(1), B2 => n9, ZN => n11
                           );
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);
   U8 : INV_X1 port map( A => S(2), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX51_19 is

   port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0);  
         Y : out std_logic);

end MUX51_19;

architecture SYN_BEHAVIORAL of MUX51_19 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n9, n10, n11, n12 : std_logic;

begin
   
   U1 : AOI22_X1 port map( A1 => C, A2 => n1, B1 => D, B2 => S(0), ZN => n10);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S(0), B2 => B, ZN => n9);
   U3 : INV_X1 port map( A => n12, ZN => Y);
   U4 : AOI22_X1 port map( A1 => n11, A2 => n3, B1 => S(2), B2 => E, ZN => n12)
                           ;
   U5 : OAI22_X1 port map( A1 => n10, A2 => n2, B1 => S(1), B2 => n9, ZN => n11
                           );
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);
   U8 : INV_X1 port map( A => S(2), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX51_18 is

   port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0);  
         Y : out std_logic);

end MUX51_18;

architecture SYN_BEHAVIORAL of MUX51_18 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n9, n10, n11, n12 : std_logic;

begin
   
   U1 : AOI22_X1 port map( A1 => C, A2 => n1, B1 => D, B2 => S(0), ZN => n10);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S(0), B2 => B, ZN => n9);
   U3 : INV_X1 port map( A => n12, ZN => Y);
   U4 : AOI22_X1 port map( A1 => n11, A2 => n3, B1 => S(2), B2 => E, ZN => n12)
                           ;
   U5 : OAI22_X1 port map( A1 => n10, A2 => n2, B1 => S(1), B2 => n9, ZN => n11
                           );
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);
   U8 : INV_X1 port map( A => S(2), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX51_17 is

   port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0);  
         Y : out std_logic);

end MUX51_17;

architecture SYN_BEHAVIORAL of MUX51_17 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n9, n10, n11, n12 : std_logic;

begin
   
   U1 : AOI22_X1 port map( A1 => C, A2 => n1, B1 => D, B2 => S(0), ZN => n10);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S(0), B2 => B, ZN => n9);
   U3 : INV_X1 port map( A => n12, ZN => Y);
   U4 : AOI22_X1 port map( A1 => n11, A2 => n3, B1 => S(2), B2 => E, ZN => n12)
                           ;
   U5 : OAI22_X1 port map( A1 => n10, A2 => n2, B1 => S(1), B2 => n9, ZN => n11
                           );
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);
   U8 : INV_X1 port map( A => S(2), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX51_16 is

   port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0);  
         Y : out std_logic);

end MUX51_16;

architecture SYN_BEHAVIORAL of MUX51_16 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n9, n10, n11, n12 : std_logic;

begin
   
   U1 : AOI22_X1 port map( A1 => C, A2 => n1, B1 => D, B2 => S(0), ZN => n10);
   U2 : INV_X1 port map( A => n12, ZN => Y);
   U3 : AOI22_X1 port map( A1 => n11, A2 => n3, B1 => S(2), B2 => E, ZN => n12)
                           ;
   U4 : OAI22_X1 port map( A1 => n10, A2 => n2, B1 => S(1), B2 => n9, ZN => n11
                           );
   U5 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S(0), B2 => B, ZN => n9);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);
   U8 : INV_X1 port map( A => S(2), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX51_15 is

   port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0);  
         Y : out std_logic);

end MUX51_15;

architecture SYN_BEHAVIORAL of MUX51_15 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n9, n10, n11, n12 : std_logic;

begin
   
   U1 : AOI22_X1 port map( A1 => C, A2 => n1, B1 => D, B2 => S(0), ZN => n10);
   U2 : INV_X1 port map( A => n12, ZN => Y);
   U3 : AOI22_X1 port map( A1 => n11, A2 => n3, B1 => S(2), B2 => E, ZN => n12)
                           ;
   U4 : OAI22_X1 port map( A1 => n10, A2 => n2, B1 => S(1), B2 => n9, ZN => n11
                           );
   U5 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S(0), B2 => B, ZN => n9);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);
   U8 : INV_X1 port map( A => S(2), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX51_14 is

   port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0);  
         Y : out std_logic);

end MUX51_14;

architecture SYN_BEHAVIORAL of MUX51_14 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n9, n10, n11, n12 : std_logic;

begin
   
   U1 : AOI22_X1 port map( A1 => C, A2 => n1, B1 => D, B2 => S(0), ZN => n10);
   U2 : INV_X1 port map( A => n12, ZN => Y);
   U3 : AOI22_X1 port map( A1 => n11, A2 => n3, B1 => S(2), B2 => E, ZN => n12)
                           ;
   U4 : OAI22_X1 port map( A1 => n10, A2 => n2, B1 => S(1), B2 => n9, ZN => n11
                           );
   U5 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S(0), B2 => B, ZN => n9);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);
   U8 : INV_X1 port map( A => S(2), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX51_13 is

   port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0);  
         Y : out std_logic);

end MUX51_13;

architecture SYN_BEHAVIORAL of MUX51_13 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n9, n10, n11, n12 : std_logic;

begin
   
   U1 : AOI22_X1 port map( A1 => C, A2 => n1, B1 => D, B2 => S(0), ZN => n10);
   U2 : INV_X1 port map( A => n12, ZN => Y);
   U3 : AOI22_X1 port map( A1 => n11, A2 => n3, B1 => S(2), B2 => E, ZN => n12)
                           ;
   U4 : OAI22_X1 port map( A1 => n10, A2 => n2, B1 => S(1), B2 => n9, ZN => n11
                           );
   U5 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S(0), B2 => B, ZN => n9);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);
   U8 : INV_X1 port map( A => S(2), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX51_12 is

   port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0);  
         Y : out std_logic);

end MUX51_12;

architecture SYN_BEHAVIORAL of MUX51_12 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n9, n10, n11, n12 : std_logic;

begin
   
   U1 : AOI22_X1 port map( A1 => C, A2 => n1, B1 => D, B2 => S(0), ZN => n10);
   U2 : INV_X1 port map( A => n12, ZN => Y);
   U3 : AOI22_X1 port map( A1 => n11, A2 => n3, B1 => S(2), B2 => E, ZN => n12)
                           ;
   U4 : OAI22_X1 port map( A1 => n10, A2 => n2, B1 => S(1), B2 => n9, ZN => n11
                           );
   U5 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S(0), B2 => B, ZN => n9);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);
   U8 : INV_X1 port map( A => S(2), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX51_11 is

   port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0);  
         Y : out std_logic);

end MUX51_11;

architecture SYN_BEHAVIORAL of MUX51_11 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n9, n10, n11, n12 : std_logic;

begin
   
   U1 : AOI22_X1 port map( A1 => C, A2 => n1, B1 => D, B2 => S(0), ZN => n10);
   U2 : INV_X1 port map( A => n12, ZN => Y);
   U3 : AOI22_X1 port map( A1 => n11, A2 => n3, B1 => S(2), B2 => E, ZN => n12)
                           ;
   U4 : OAI22_X1 port map( A1 => n10, A2 => n2, B1 => S(1), B2 => n9, ZN => n11
                           );
   U5 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S(0), B2 => B, ZN => n9);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);
   U8 : INV_X1 port map( A => S(2), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX51_10 is

   port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0);  
         Y : out std_logic);

end MUX51_10;

architecture SYN_BEHAVIORAL of MUX51_10 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n9, n10, n11, n12 : std_logic;

begin
   
   U1 : AOI22_X1 port map( A1 => C, A2 => n1, B1 => D, B2 => S(0), ZN => n10);
   U2 : INV_X1 port map( A => n12, ZN => Y);
   U3 : AOI22_X1 port map( A1 => n11, A2 => n3, B1 => S(2), B2 => E, ZN => n12)
                           ;
   U4 : OAI22_X1 port map( A1 => n10, A2 => n2, B1 => S(1), B2 => n9, ZN => n11
                           );
   U5 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S(0), B2 => B, ZN => n9);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);
   U8 : INV_X1 port map( A => S(2), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX51_9 is

   port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0);  
         Y : out std_logic);

end MUX51_9;

architecture SYN_BEHAVIORAL of MUX51_9 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n9, n10, n11, n12 : std_logic;

begin
   
   U1 : AOI22_X1 port map( A1 => C, A2 => n1, B1 => D, B2 => S(0), ZN => n10);
   U2 : INV_X1 port map( A => n12, ZN => Y);
   U3 : AOI22_X1 port map( A1 => n11, A2 => n3, B1 => S(2), B2 => E, ZN => n12)
                           ;
   U4 : OAI22_X1 port map( A1 => n10, A2 => n2, B1 => S(1), B2 => n9, ZN => n11
                           );
   U5 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S(0), B2 => B, ZN => n9);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);
   U8 : INV_X1 port map( A => S(2), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX51_8 is

   port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0);  
         Y : out std_logic);

end MUX51_8;

architecture SYN_BEHAVIORAL of MUX51_8 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n9, n10, n11, n12 : std_logic;

begin
   
   U1 : AOI22_X1 port map( A1 => C, A2 => n1, B1 => D, B2 => S(0), ZN => n10);
   U2 : INV_X1 port map( A => n12, ZN => Y);
   U3 : AOI22_X1 port map( A1 => n11, A2 => n3, B1 => S(2), B2 => E, ZN => n12)
                           ;
   U4 : OAI22_X1 port map( A1 => n10, A2 => n2, B1 => S(1), B2 => n9, ZN => n11
                           );
   U5 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S(0), B2 => B, ZN => n9);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);
   U8 : INV_X1 port map( A => S(2), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX51_7 is

   port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0);  
         Y : out std_logic);

end MUX51_7;

architecture SYN_BEHAVIORAL of MUX51_7 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n9, n10, n11, n12 : std_logic;

begin
   
   U1 : AOI22_X1 port map( A1 => C, A2 => n1, B1 => D, B2 => S(0), ZN => n10);
   U2 : INV_X1 port map( A => n12, ZN => Y);
   U3 : AOI22_X1 port map( A1 => n11, A2 => n3, B1 => S(2), B2 => E, ZN => n12)
                           ;
   U4 : OAI22_X1 port map( A1 => n10, A2 => n2, B1 => S(1), B2 => n9, ZN => n11
                           );
   U5 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S(0), B2 => B, ZN => n9);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);
   U8 : INV_X1 port map( A => S(2), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX51_6 is

   port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0);  
         Y : out std_logic);

end MUX51_6;

architecture SYN_BEHAVIORAL of MUX51_6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n9, n10, n11, n12 : std_logic;

begin
   
   U1 : AOI22_X1 port map( A1 => C, A2 => n1, B1 => D, B2 => S(0), ZN => n10);
   U2 : INV_X1 port map( A => n12, ZN => Y);
   U3 : AOI22_X1 port map( A1 => n11, A2 => n3, B1 => S(2), B2 => E, ZN => n12)
                           ;
   U4 : OAI22_X1 port map( A1 => n10, A2 => n2, B1 => S(1), B2 => n9, ZN => n11
                           );
   U5 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S(0), B2 => B, ZN => n9);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);
   U8 : INV_X1 port map( A => S(2), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX51_5 is

   port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0);  
         Y : out std_logic);

end MUX51_5;

architecture SYN_BEHAVIORAL of MUX51_5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n9, n10, n11, n12 : std_logic;

begin
   
   U1 : AOI22_X1 port map( A1 => C, A2 => n1, B1 => D, B2 => S(0), ZN => n10);
   U2 : INV_X1 port map( A => n12, ZN => Y);
   U3 : AOI22_X1 port map( A1 => n11, A2 => n3, B1 => S(2), B2 => E, ZN => n12)
                           ;
   U4 : OAI22_X1 port map( A1 => n10, A2 => n2, B1 => S(1), B2 => n9, ZN => n11
                           );
   U5 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S(0), B2 => B, ZN => n9);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);
   U8 : INV_X1 port map( A => S(2), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX51_4 is

   port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0);  
         Y : out std_logic);

end MUX51_4;

architecture SYN_BEHAVIORAL of MUX51_4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n9, n10, n11, n12 : std_logic;

begin
   
   U1 : AOI22_X1 port map( A1 => C, A2 => n1, B1 => D, B2 => S(0), ZN => n10);
   U2 : INV_X1 port map( A => n12, ZN => Y);
   U3 : AOI22_X1 port map( A1 => n11, A2 => n3, B1 => S(2), B2 => E, ZN => n12)
                           ;
   U4 : OAI22_X1 port map( A1 => n10, A2 => n2, B1 => S(1), B2 => n9, ZN => n11
                           );
   U5 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S(0), B2 => B, ZN => n9);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);
   U8 : INV_X1 port map( A => S(2), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX51_3 is

   port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0);  
         Y : out std_logic);

end MUX51_3;

architecture SYN_BEHAVIORAL of MUX51_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n9, n10, n11, n12 : std_logic;

begin
   
   U1 : AOI22_X1 port map( A1 => C, A2 => n1, B1 => D, B2 => S(0), ZN => n10);
   U2 : INV_X1 port map( A => n12, ZN => Y);
   U3 : AOI22_X1 port map( A1 => n11, A2 => n3, B1 => S(2), B2 => E, ZN => n12)
                           ;
   U4 : OAI22_X1 port map( A1 => n10, A2 => n2, B1 => S(1), B2 => n9, ZN => n11
                           );
   U5 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S(0), B2 => B, ZN => n9);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);
   U8 : INV_X1 port map( A => S(2), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX51_2 is

   port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0);  
         Y : out std_logic);

end MUX51_2;

architecture SYN_BEHAVIORAL of MUX51_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n9, n10, n11, n12 : std_logic;

begin
   
   U1 : AOI22_X1 port map( A1 => C, A2 => n1, B1 => D, B2 => S(0), ZN => n10);
   U2 : INV_X1 port map( A => n12, ZN => Y);
   U3 : AOI22_X1 port map( A1 => n11, A2 => n3, B1 => S(2), B2 => E, ZN => n12)
                           ;
   U4 : OAI22_X1 port map( A1 => n10, A2 => n2, B1 => S(1), B2 => n9, ZN => n11
                           );
   U5 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S(0), B2 => B, ZN => n9);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);
   U8 : INV_X1 port map( A => S(2), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX51_1 is

   port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0);  
         Y : out std_logic);

end MUX51_1;

architecture SYN_BEHAVIORAL of MUX51_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n9, n10, n11, n12 : std_logic;

begin
   
   U1 : AOI22_X1 port map( A1 => C, A2 => n1, B1 => D, B2 => S(0), ZN => n10);
   U2 : INV_X1 port map( A => n12, ZN => Y);
   U3 : AOI22_X1 port map( A1 => n11, A2 => n3, B1 => S(2), B2 => E, ZN => n12)
                           ;
   U4 : OAI22_X1 port map( A1 => n10, A2 => n2, B1 => S(1), B2 => n9, ZN => n11
                           );
   U5 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S(0), B2 => B, ZN => n9);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);
   U8 : INV_X1 port map( A => S(2), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_167 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_167;

architecture SYN_BEHAVIORAL_1 of MUX41_167 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X4
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : OAI211_X4 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U2 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U3 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U4 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U5 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_166 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_166;

architecture SYN_BEHAVIORAL_1 of MUX41_166 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X4
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : OAI211_X4 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U2 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U3 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U4 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U5 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_165 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_165;

architecture SYN_BEHAVIORAL_1 of MUX41_165 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X4
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : OAI211_X4 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U2 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U3 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U4 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U5 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_164 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_164;

architecture SYN_BEHAVIORAL_1 of MUX41_164 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X4
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : OAI211_X4 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U2 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U3 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U4 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U5 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_163 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_163;

architecture SYN_BEHAVIORAL_1 of MUX41_163 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X4
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : OAI211_X4 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U2 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U3 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U4 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U5 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_162 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_162;

architecture SYN_BEHAVIORAL_1 of MUX41_162 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X4
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : OAI211_X4 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U2 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U3 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_161 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_161;

architecture SYN_BEHAVIORAL_1 of MUX41_161 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X4
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : OAI211_X4 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U2 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U3 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_160 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_160;

architecture SYN_BEHAVIORAL_1 of MUX41_160 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X2
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U1 : OAI211_X2 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U2 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U3 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_159 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_159;

architecture SYN_BEHAVIORAL_1 of MUX41_159 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X2
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U1 : OAI211_X2 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U2 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U3 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_158 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_158;

architecture SYN_BEHAVIORAL_1 of MUX41_158 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X2
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U1 : OAI211_X2 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U2 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U3 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_157 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_157;

architecture SYN_BEHAVIORAL_1 of MUX41_157 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X2
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U1 : OAI211_X2 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U2 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U3 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_156 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_156;

architecture SYN_BEHAVIORAL_1 of MUX41_156 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X2
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : OAI211_X2 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U2 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U3 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U4 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U5 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_155 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_155;

architecture SYN_BEHAVIORAL_1 of MUX41_155 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X2
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : OAI211_X2 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U2 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U3 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U4 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U5 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_154 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_154;

architecture SYN_BEHAVIORAL_1 of MUX41_154 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X2
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : OAI211_X2 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U2 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U3 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U4 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U5 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_153 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_153;

architecture SYN_BEHAVIORAL_1 of MUX41_153 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X2
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : OAI211_X2 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U2 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U3 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U4 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U5 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_152 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_152;

architecture SYN_BEHAVIORAL_1 of MUX41_152 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X2
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : OAI211_X2 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U2 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U3 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U4 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U5 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_151 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_151;

architecture SYN_BEHAVIORAL_1 of MUX41_151 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X2
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U1 : OAI211_X2 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U2 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U3 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_150 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_150;

architecture SYN_BEHAVIORAL_1 of MUX41_150 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X2
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U1 : OAI211_X2 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U2 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U3 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_149 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_149;

architecture SYN_BEHAVIORAL_1 of MUX41_149 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X2
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U1 : OAI211_X2 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U2 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U3 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_148 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_148;

architecture SYN_BEHAVIORAL_1 of MUX41_148 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X2
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U1 : OAI211_X2 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U2 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U3 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_147 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_147;

architecture SYN_BEHAVIORAL_1 of MUX41_147 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X2
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U1 : OAI211_X2 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U2 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U3 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_146 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_146;

architecture SYN_BEHAVIORAL_1 of MUX41_146 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X2
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U1 : OAI211_X2 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U2 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U3 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_145 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_145;

architecture SYN_BEHAVIORAL_1 of MUX41_145 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X2
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : OAI211_X2 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U2 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U3 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U4 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U5 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_144 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_144;

architecture SYN_BEHAVIORAL_1 of MUX41_144 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X4
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : OAI211_X4 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U2 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U3 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U4 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U5 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_143 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_143;

architecture SYN_BEHAVIORAL_1 of MUX41_143 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X4
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : OAI211_X4 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U2 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U3 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U4 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U5 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_142 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_142;

architecture SYN_BEHAVIORAL_1 of MUX41_142 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X4
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : OAI211_X4 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U2 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U3 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_141 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_141;

architecture SYN_BEHAVIORAL_1 of MUX41_141 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X4
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : OAI211_X4 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U2 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U3 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_140 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_140;

architecture SYN_BEHAVIORAL_1 of MUX41_140 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X4
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : OAI211_X4 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U2 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U3 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_139 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_139;

architecture SYN_BEHAVIORAL_1 of MUX41_139 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X2
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U1 : OAI211_X2 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U2 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U3 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_138 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_138;

architecture SYN_BEHAVIORAL_1 of MUX41_138 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X2
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U1 : OAI211_X2 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U2 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U3 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_137 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_137;

architecture SYN_BEHAVIORAL_1 of MUX41_137 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U2 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U3 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_136 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_136;

architecture SYN_BEHAVIORAL_1 of MUX41_136 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U2 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U3 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U5 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_135 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_135;

architecture SYN_BEHAVIORAL_1 of MUX41_135 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X2
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U1 : OAI211_X2 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U2 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U3 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U4 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U5 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_134 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_134;

architecture SYN_BEHAVIORAL_1 of MUX41_134 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U2 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U3 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U5 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_133 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_133;

architecture SYN_BEHAVIORAL_1 of MUX41_133 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U2 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U3 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U4 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U5 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_132 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_132;

architecture SYN_BEHAVIORAL_1 of MUX41_132 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U2 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U3 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U5 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_131 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_131;

architecture SYN_BEHAVIORAL_1 of MUX41_131 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U2 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U3 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_130 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_130;

architecture SYN_BEHAVIORAL_1 of MUX41_130 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U2 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U3 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_129 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_129;

architecture SYN_BEHAVIORAL_1 of MUX41_129 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U2 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U3 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_128 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_128;

architecture SYN_BEHAVIORAL_1 of MUX41_128 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U2 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U3 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_127 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_127;

architecture SYN_BEHAVIORAL_1 of MUX41_127 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U2 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U3 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_126 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_126;

architecture SYN_BEHAVIORAL_1 of MUX41_126 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U2 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U3 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_125 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_125;

architecture SYN_BEHAVIORAL_1 of MUX41_125 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U2 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U3 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U5 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_124 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_124;

architecture SYN_BEHAVIORAL_1 of MUX41_124 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U2 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U3 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U5 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_123 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_123;

architecture SYN_BEHAVIORAL_1 of MUX41_123 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U2 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U3 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U5 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_122 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_122;

architecture SYN_BEHAVIORAL_1 of MUX41_122 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U2 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U3 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U5 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_121 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_121;

architecture SYN_BEHAVIORAL_1 of MUX41_121 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U2 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U3 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U5 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_120 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_120;

architecture SYN_BEHAVIORAL_1 of MUX41_120 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U2 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U3 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_119 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_119;

architecture SYN_BEHAVIORAL_1 of MUX41_119 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U2 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U3 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_118 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_118;

architecture SYN_BEHAVIORAL_1 of MUX41_118 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U2 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U3 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_117 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_117;

architecture SYN_BEHAVIORAL_1 of MUX41_117 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U2 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U3 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_116 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_116;

architecture SYN_BEHAVIORAL_1 of MUX41_116 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U2 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U3 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_115 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_115;

architecture SYN_BEHAVIORAL_1 of MUX41_115 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U2 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U3 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_114 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_114;

architecture SYN_BEHAVIORAL_1 of MUX41_114 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U2 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U3 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U5 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_113 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_113;

architecture SYN_BEHAVIORAL_1 of MUX41_113 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U2 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U3 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U5 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_112 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_112;

architecture SYN_BEHAVIORAL_1 of MUX41_112 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U2 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U3 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U5 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_111 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_111;

architecture SYN_BEHAVIORAL_1 of MUX41_111 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U2 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U3 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_110 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_110;

architecture SYN_BEHAVIORAL_1 of MUX41_110 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U2 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U3 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_109 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_109;

architecture SYN_BEHAVIORAL_1 of MUX41_109 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U2 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U3 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_108 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_108;

architecture SYN_BEHAVIORAL_1 of MUX41_108 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U2 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U3 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_107 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_107;

architecture SYN_BEHAVIORAL_1 of MUX41_107 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U2 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U3 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_106 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_106;

architecture SYN_BEHAVIORAL_1 of MUX41_106 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U2 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U3 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_105 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_105;

architecture SYN_BEHAVIORAL_1 of MUX41_105 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U2 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U3 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_104 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_104;

architecture SYN_BEHAVIORAL_1 of MUX41_104 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U2 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U3 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U5 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_103 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_103;

architecture SYN_BEHAVIORAL_1 of MUX41_103 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U2 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U3 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U5 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_102 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_102;

architecture SYN_BEHAVIORAL_1 of MUX41_102 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U2 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U3 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U5 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_101 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_101;

architecture SYN_BEHAVIORAL_1 of MUX41_101 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U2 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U3 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U5 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_100 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_100;

architecture SYN_BEHAVIORAL_1 of MUX41_100 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U2 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U3 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U5 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_99 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_99;

architecture SYN_BEHAVIORAL_1 of MUX41_99 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U2 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U3 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_98 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_98;

architecture SYN_BEHAVIORAL_1 of MUX41_98 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U2 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U3 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_97 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_97;

architecture SYN_BEHAVIORAL_1 of MUX41_97 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U2 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U3 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_96 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_96;

architecture SYN_BEHAVIORAL_1 of MUX41_96 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U2 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U3 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_95 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_95;

architecture SYN_BEHAVIORAL_1 of MUX41_95 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U2 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U3 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_94 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_94;

architecture SYN_BEHAVIORAL_1 of MUX41_94 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U2 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U3 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_93 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_93;

architecture SYN_BEHAVIORAL_1 of MUX41_93 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U2 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U3 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U5 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_92 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_92;

architecture SYN_BEHAVIORAL_1 of MUX41_92 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U2 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U3 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U5 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_91 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_91;

architecture SYN_BEHAVIORAL_1 of MUX41_91 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U2 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U3 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U5 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_90 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_90;

architecture SYN_BEHAVIORAL_1 of MUX41_90 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U2 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U3 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U5 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_89 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_89;

architecture SYN_BEHAVIORAL_1 of MUX41_89 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U2 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U3 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U5 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_88 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_88;

architecture SYN_BEHAVIORAL_1 of MUX41_88 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U2 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U3 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_87 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_87;

architecture SYN_BEHAVIORAL_1 of MUX41_87 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U2 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U3 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_86 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_86;

architecture SYN_BEHAVIORAL_1 of MUX41_86 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U2 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U3 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_85 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_85;

architecture SYN_BEHAVIORAL_1 of MUX41_85 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U2 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U3 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_84 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_84;

architecture SYN_BEHAVIORAL_1 of MUX41_84 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U2 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U3 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_83 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_83;

architecture SYN_BEHAVIORAL_1 of MUX41_83 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U2 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U3 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_82 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_82;

architecture SYN_BEHAVIORAL_1 of MUX41_82 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U2 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U3 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U5 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_81 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_81;

architecture SYN_BEHAVIORAL_1 of MUX41_81 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U2 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U3 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U5 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_80 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_80;

architecture SYN_BEHAVIORAL_1 of MUX41_80 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U2 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U3 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U5 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_79 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_79;

architecture SYN_BEHAVIORAL_1 of MUX41_79 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U2 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U3 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_78 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_78;

architecture SYN_BEHAVIORAL_1 of MUX41_78 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U2 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U3 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_77 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_77;

architecture SYN_BEHAVIORAL_1 of MUX41_77 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U2 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U3 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_76 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_76;

architecture SYN_BEHAVIORAL_1 of MUX41_76 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U2 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U3 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_75 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_75;

architecture SYN_BEHAVIORAL_1 of MUX41_75 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U2 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U3 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_74 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_74;

architecture SYN_BEHAVIORAL_1 of MUX41_74 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U2 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U3 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_73 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_73;

architecture SYN_BEHAVIORAL_1 of MUX41_73 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U2 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U3 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_72 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_72;

architecture SYN_BEHAVIORAL_1 of MUX41_72 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U2 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U3 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U4 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U5 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_71 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_71;

architecture SYN_BEHAVIORAL_1 of MUX41_71 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U2 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U3 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U4 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U5 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_70 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_70;

architecture SYN_BEHAVIORAL_1 of MUX41_70 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U2 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U3 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U5 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_69 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_69;

architecture SYN_BEHAVIORAL_1 of MUX41_69 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U2 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U3 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U5 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_68 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_68;

architecture SYN_BEHAVIORAL_1 of MUX41_68 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U2 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U3 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U5 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_67 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_67;

architecture SYN_BEHAVIORAL_1 of MUX41_67 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U2 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U3 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_66 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_66;

architecture SYN_BEHAVIORAL_1 of MUX41_66 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U2 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U3 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_65 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_65;

architecture SYN_BEHAVIORAL_1 of MUX41_65 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U2 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U3 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_64 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_64;

architecture SYN_BEHAVIORAL_1 of MUX41_64 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U2 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U3 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_63 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_63;

architecture SYN_BEHAVIORAL_1 of MUX41_63 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U2 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U3 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_62 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_62;

architecture SYN_BEHAVIORAL_1 of MUX41_62 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U2 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U3 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_61 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_61;

architecture SYN_BEHAVIORAL_1 of MUX41_61 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U2 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U3 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U5 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_60 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_60;

architecture SYN_BEHAVIORAL_1 of MUX41_60 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U2 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U3 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U5 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_59 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_59;

architecture SYN_BEHAVIORAL_1 of MUX41_59 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U2 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U3 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U5 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_58 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_58;

architecture SYN_BEHAVIORAL_1 of MUX41_58 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U2 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U3 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U5 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_57 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_57;

architecture SYN_BEHAVIORAL_1 of MUX41_57 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U2 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U3 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U5 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_56 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_56;

architecture SYN_BEHAVIORAL_1 of MUX41_56 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U2 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U3 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_55 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_55;

architecture SYN_BEHAVIORAL_1 of MUX41_55 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U2 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U3 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_54 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_54;

architecture SYN_BEHAVIORAL_1 of MUX41_54 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U2 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U3 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_53 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_53;

architecture SYN_BEHAVIORAL_1 of MUX41_53 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U2 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U3 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_52 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_52;

architecture SYN_BEHAVIORAL_1 of MUX41_52 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U2 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U3 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_51 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_51;

architecture SYN_BEHAVIORAL_1 of MUX41_51 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U2 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U3 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_50 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_50;

architecture SYN_BEHAVIORAL_1 of MUX41_50 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U2 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U3 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U5 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_49 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_49;

architecture SYN_BEHAVIORAL_1 of MUX41_49 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U2 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U3 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U5 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_48 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_48;

architecture SYN_BEHAVIORAL_1 of MUX41_48 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U2 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U3 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U5 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_47 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_47;

architecture SYN_BEHAVIORAL_1 of MUX41_47 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U2 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U3 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U5 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_46 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_46;

architecture SYN_BEHAVIORAL_1 of MUX41_46 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U2 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U3 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U5 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_45 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_45;

architecture SYN_BEHAVIORAL_1 of MUX41_45 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U2 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U3 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_44 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_44;

architecture SYN_BEHAVIORAL_1 of MUX41_44 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U2 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U3 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_43 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_43;

architecture SYN_BEHAVIORAL_1 of MUX41_43 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U2 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U3 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_42 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_42;

architecture SYN_BEHAVIORAL_1 of MUX41_42 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U2 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U3 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_41 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_41;

architecture SYN_BEHAVIORAL_1 of MUX41_41 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U2 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U3 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_40 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_40;

architecture SYN_BEHAVIORAL_1 of MUX41_40 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U2 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U3 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_39 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_39;

architecture SYN_BEHAVIORAL_1 of MUX41_39 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U2 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U3 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_38 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_38;

architecture SYN_BEHAVIORAL_1 of MUX41_38 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U2 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U3 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_37 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_37;

architecture SYN_BEHAVIORAL_1 of MUX41_37 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U2 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U3 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_36 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_36;

architecture SYN_BEHAVIORAL_1 of MUX41_36 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U2 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U3 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_35 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_35;

architecture SYN_BEHAVIORAL_1 of MUX41_35 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U2 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U3 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_34 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_34;

architecture SYN_BEHAVIORAL_1 of MUX41_34 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U2 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U3 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U4 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U5 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_33 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_33;

architecture SYN_BEHAVIORAL_1 of MUX41_33 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U2 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U3 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U4 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U5 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_32 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_32;

architecture SYN_BEHAVIORAL_1 of MUX41_32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U2 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U3 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U4 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U5 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_31 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_31;

architecture SYN_BEHAVIORAL_1 of MUX41_31 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U2 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U3 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U4 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U5 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_30 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_30;

architecture SYN_BEHAVIORAL_1 of MUX41_30 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U2 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U3 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U4 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U5 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_29 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_29;

architecture SYN_BEHAVIORAL_1 of MUX41_29 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U2 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U3 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U4 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U5 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_28 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_28;

architecture SYN_BEHAVIORAL_1 of MUX41_28 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U2 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U3 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U4 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U5 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_27 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_27;

architecture SYN_BEHAVIORAL_1 of MUX41_27 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U2 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U3 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U4 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U5 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_26 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_26;

architecture SYN_BEHAVIORAL_1 of MUX41_26 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U2 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U3 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U4 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U5 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_25 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_25;

architecture SYN_BEHAVIORAL_1 of MUX41_25 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U2 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U3 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U4 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U5 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_24 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_24;

architecture SYN_BEHAVIORAL_1 of MUX41_24 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U2 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U3 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U4 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U5 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_23 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_23;

architecture SYN_BEHAVIORAL_1_architecture of MUX41_23 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U2 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U3 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U4 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U5 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_22 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_22;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX41_22 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U2 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U3 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U4 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U5 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_21 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_21;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX41_21 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U2 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U3 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U4 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U5 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_20 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_20;

architecture SYN_BEHAVIORAL_1_architecture4 of MUX41_20 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U2 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U3 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U4 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U5 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_19 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_19;

architecture SYN_BEHAVIORAL_1_architecture5 of MUX41_19 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U2 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U3 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U4 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U5 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1_architecture5;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_18 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_18;

architecture SYN_BEHAVIORAL_1_architecture6 of MUX41_18 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U2 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U3 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U4 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U5 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1_architecture6;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_17 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_17;

architecture SYN_BEHAVIORAL_1_architecture7 of MUX41_17 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U2 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U3 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U4 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U5 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1_architecture7;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_16 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_16;

architecture SYN_BEHAVIORAL_1 of MUX41_16 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U2 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U3 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U4 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U5 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_15 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_15;

architecture SYN_BEHAVIORAL_1_architecture of MUX41_15 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U2 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U3 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U4 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U5 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_14 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_14;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX41_14 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U2 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U3 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U4 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U5 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_13 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_13;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX41_13 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U2 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U3 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U4 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U5 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_12 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_12;

architecture SYN_BEHAVIORAL_1_architecture4 of MUX41_12 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U2 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U3 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U4 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U5 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_11 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_11;

architecture SYN_BEHAVIORAL_1_architecture5 of MUX41_11 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U2 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U3 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U4 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U5 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1_architecture5;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_10 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_10;

architecture SYN_BEHAVIORAL_1_architecture6 of MUX41_10 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U2 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U3 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U4 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U5 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1_architecture6;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_9 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_9;

architecture SYN_BEHAVIORAL_1_architecture7 of MUX41_9 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U2 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U3 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U4 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U5 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1_architecture7;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_8 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_8;

architecture SYN_BEHAVIORAL_1 of MUX41_8 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12, n13 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n2, A2 => n8, A3 => A, ZN => n10);
   U1 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => n9);
   U2 : OAI211_X1 port map( C1 => n13, C2 => n12, A => n11, B => n10, ZN => Y);
   U3 : NAND2_X1 port map( A1 => B, A2 => n13, ZN => n11);
   U4 : AOI22_X1 port map( A1 => D, A2 => n1, B1 => n9, B2 => C, ZN => n12);
   U5 : NOR2_X1 port map( A1 => n2, A2 => S(1), ZN => n13);
   U6 : INV_X1 port map( A => n2, ZN => n1);
   U7 : INV_X1 port map( A => S(0), ZN => n2);
   U9 : INV_X1 port map( A => S(1), ZN => n8);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_7 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_7;

architecture SYN_BEHAVIORAL_1_architecture of MUX41_7 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U2 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U3 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U4 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U5 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_6 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_6;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX41_6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U2 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U3 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U4 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U5 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_5 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_5;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX41_5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U2 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U3 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U4 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U5 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_4 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_4;

architecture SYN_BEHAVIORAL_1_architecture4 of MUX41_4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U2 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U3 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U4 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U5 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_3 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_3;

architecture SYN_BEHAVIORAL_1_architecture5 of MUX41_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U2 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U3 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U4 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U5 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1_architecture5;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_2 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_2;

architecture SYN_BEHAVIORAL_1_architecture6 of MUX41_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U2 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U3 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1_architecture6;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_1 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_1;

architecture SYN_BEHAVIORAL_1_architecture7 of MUX41_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n9);
   U1 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n8, B2 => C, ZN => n11);
   U2 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n8);
   U3 : OAI211_X1 port map( C1 => n12, C2 => n11, A => n10, B => n9, ZN => Y);
   U4 : NAND2_X1 port map( A1 => B, A2 => n12, ZN => n10);
   U5 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n12);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1_architecture7;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity sum_generator_n_bit32_n_CSB8_1 is

   port( A, B : in std_logic_vector (31 downto 0);  C_in : in std_logic_vector 
         (7 downto 0);  S : out std_logic_vector (31 downto 0));

end sum_generator_n_bit32_n_CSB8_1;

architecture SYN_STRUCTURAL of sum_generator_n_bit32_n_CSB8_1 is

   component carry_select_block_n4_49
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_n4_50
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_n4_51
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_n4_52
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_n4_53
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_n4_54
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_n4_55
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_n4_56
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;

begin
   
   csb_0 : carry_select_block_n4_56 port map( A(3) => A(3), A(2) => A(2), A(1) 
                           => A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), 
                           B(1) => B(1), B(0) => B(0), C_sel => C_in(0), S(3) 
                           => S(3), S(2) => S(2), S(1) => S(1), S(0) => S(0));
   csb_1 : carry_select_block_n4_55 port map( A(3) => A(7), A(2) => A(6), A(1) 
                           => A(5), A(0) => A(4), B(3) => B(7), B(2) => B(6), 
                           B(1) => B(5), B(0) => B(4), C_sel => C_in(1), S(3) 
                           => S(7), S(2) => S(6), S(1) => S(5), S(0) => S(4));
   csb_2 : carry_select_block_n4_54 port map( A(3) => A(11), A(2) => A(10), 
                           A(1) => A(9), A(0) => A(8), B(3) => B(11), B(2) => 
                           B(10), B(1) => B(9), B(0) => B(8), C_sel => C_in(2),
                           S(3) => S(11), S(2) => S(10), S(1) => S(9), S(0) => 
                           S(8));
   csb_3 : carry_select_block_n4_53 port map( A(3) => A(15), A(2) => A(14), 
                           A(1) => A(13), A(0) => A(12), B(3) => B(15), B(2) =>
                           B(14), B(1) => B(13), B(0) => B(12), C_sel => 
                           C_in(3), S(3) => S(15), S(2) => S(14), S(1) => S(13)
                           , S(0) => S(12));
   csb_4 : carry_select_block_n4_52 port map( A(3) => A(19), A(2) => A(18), 
                           A(1) => A(17), A(0) => A(16), B(3) => B(19), B(2) =>
                           B(18), B(1) => B(17), B(0) => B(16), C_sel => 
                           C_in(4), S(3) => S(19), S(2) => S(18), S(1) => S(17)
                           , S(0) => S(16));
   csb_5 : carry_select_block_n4_51 port map( A(3) => A(23), A(2) => A(22), 
                           A(1) => A(21), A(0) => A(20), B(3) => B(23), B(2) =>
                           B(22), B(1) => B(21), B(0) => B(20), C_sel => 
                           C_in(5), S(3) => S(23), S(2) => S(22), S(1) => S(21)
                           , S(0) => S(20));
   csb_6 : carry_select_block_n4_50 port map( A(3) => A(27), A(2) => A(26), 
                           A(1) => A(25), A(0) => A(24), B(3) => B(27), B(2) =>
                           B(26), B(1) => B(25), B(0) => B(24), C_sel => 
                           C_in(6), S(3) => S(27), S(2) => S(26), S(1) => S(25)
                           , S(0) => S(24));
   csb_7 : carry_select_block_n4_49 port map( A(3) => A(31), A(2) => A(30), 
                           A(1) => A(29), A(0) => A(28), B(3) => B(31), B(2) =>
                           B(30), B(1) => B(29), B(0) => B(28), C_sel => 
                           C_in(7), S(3) => S(31), S(2) => S(30), S(1) => S(29)
                           , S(0) => S(28));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_1 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co : 
         out std_logic_vector (7 downto 0));

end CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_1;

architecture SYN_structural of CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_1 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component G_BLOCK_52
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component G_BLOCK_53
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component G_BLOCK_54
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component G_BLOCK_55
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component G_BLOCK_56
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component G_BLOCK_57
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component PG_BLOCK_190
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_191
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component G_BLOCK_58
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component PG_BLOCK_192
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_193
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_194
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component G_BLOCK_59
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component PG_BLOCK_195
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_196
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_197
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_198
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_199
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_200
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_201
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component G_BLOCK_60
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component PG_BLOCK_202
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_203
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_204
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_205
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_206
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_207
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_208
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_209
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_210
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_211
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_212
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_213
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_214
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_215
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_216
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component pg_net_190
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_191
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_192
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_193
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_194
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_195
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_196
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_197
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_198
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_199
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_200
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_201
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_202
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_203
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_204
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_205
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_206
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_207
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_208
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_209
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_210
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_211
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_212
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_213
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_214
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_215
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_216
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_217
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_218
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_219
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_220
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   signal Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, Co_2_port, 
      Co_1_port, Co_0_port, g_vector_4_31_port, g_vector_4_27_port, 
      g_vector_3_31_port, g_vector_3_23_port, g_vector_3_15_port, 
      g_vector_2_31_port, g_vector_2_27_port, g_vector_2_23_port, 
      g_vector_2_19_port, g_vector_2_15_port, g_vector_2_11_port, 
      g_vector_2_7_port, g_vector_1_31_port, g_vector_1_29_port, 
      g_vector_1_27_port, g_vector_1_25_port, g_vector_1_23_port, 
      g_vector_1_21_port, g_vector_1_19_port, g_vector_1_17_port, 
      g_vector_1_15_port, g_vector_1_13_port, g_vector_1_11_port, 
      g_vector_1_9_port, g_vector_1_7_port, g_vector_1_5_port, 
      g_vector_1_3_port, g_vector_1_1_port, g_vector_0_31_port, 
      g_vector_0_30_port, g_vector_0_29_port, g_vector_0_28_port, 
      g_vector_0_27_port, g_vector_0_26_port, g_vector_0_25_port, 
      g_vector_0_24_port, g_vector_0_23_port, g_vector_0_22_port, 
      g_vector_0_21_port, g_vector_0_20_port, g_vector_0_19_port, 
      g_vector_0_18_port, g_vector_0_17_port, g_vector_0_16_port, 
      g_vector_0_15_port, g_vector_0_14_port, g_vector_0_13_port, 
      g_vector_0_12_port, g_vector_0_11_port, g_vector_0_10_port, 
      g_vector_0_9_port, g_vector_0_8_port, g_vector_0_7_port, 
      g_vector_0_6_port, g_vector_0_5_port, g_vector_0_4_port, 
      g_vector_0_3_port, g_vector_0_2_port, g_vector_0_1_port, 
      g_vector_0_0_port, p_vector_4_31_port, p_vector_4_27_port, 
      p_vector_3_31_port, p_vector_3_23_port, p_vector_3_15_port, 
      p_vector_2_31_port, p_vector_2_27_port, p_vector_2_23_port, 
      p_vector_2_19_port, p_vector_2_15_port, p_vector_2_11_port, 
      p_vector_2_7_port, p_vector_1_31_port, p_vector_1_29_port, 
      p_vector_1_27_port, p_vector_1_25_port, p_vector_1_23_port, 
      p_vector_1_21_port, p_vector_1_19_port, p_vector_1_17_port, 
      p_vector_1_15_port, p_vector_1_13_port, p_vector_1_11_port, 
      p_vector_1_9_port, p_vector_1_7_port, p_vector_1_5_port, 
      p_vector_1_3_port, p_vector_0_31_port, p_vector_0_30_port, 
      p_vector_0_29_port, p_vector_0_28_port, p_vector_0_27_port, 
      p_vector_0_26_port, p_vector_0_25_port, p_vector_0_24_port, 
      p_vector_0_23_port, p_vector_0_22_port, p_vector_0_21_port, 
      p_vector_0_20_port, p_vector_0_19_port, p_vector_0_18_port, 
      p_vector_0_17_port, p_vector_0_16_port, p_vector_0_15_port, 
      p_vector_0_14_port, p_vector_0_13_port, p_vector_0_12_port, 
      p_vector_0_11_port, p_vector_0_10_port, p_vector_0_9_port, 
      p_vector_0_8_port, p_vector_0_7_port, p_vector_0_6_port, 
      p_vector_0_5_port, p_vector_0_4_port, p_vector_0_3_port, 
      p_vector_0_2_port, p_vector_0_1_port, n1, n2, n4 : std_logic;

begin
   Co <= ( Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, Co_2_port, 
      Co_1_port, Co_0_port );
   
   pg_network_31 : pg_net_220 port map( a => A(31), b => B(31), p => 
                           p_vector_0_31_port, g => g_vector_0_31_port);
   pg_network_30 : pg_net_219 port map( a => A(30), b => B(30), p => 
                           p_vector_0_30_port, g => g_vector_0_30_port);
   pg_network_29 : pg_net_218 port map( a => A(29), b => B(29), p => 
                           p_vector_0_29_port, g => g_vector_0_29_port);
   pg_network_28 : pg_net_217 port map( a => A(28), b => B(28), p => 
                           p_vector_0_28_port, g => g_vector_0_28_port);
   pg_network_27 : pg_net_216 port map( a => A(27), b => B(27), p => 
                           p_vector_0_27_port, g => g_vector_0_27_port);
   pg_network_26 : pg_net_215 port map( a => A(26), b => B(26), p => 
                           p_vector_0_26_port, g => g_vector_0_26_port);
   pg_network_25 : pg_net_214 port map( a => A(25), b => B(25), p => 
                           p_vector_0_25_port, g => g_vector_0_25_port);
   pg_network_24 : pg_net_213 port map( a => A(24), b => B(24), p => 
                           p_vector_0_24_port, g => g_vector_0_24_port);
   pg_network_23 : pg_net_212 port map( a => A(23), b => B(23), p => 
                           p_vector_0_23_port, g => g_vector_0_23_port);
   pg_network_22 : pg_net_211 port map( a => A(22), b => B(22), p => 
                           p_vector_0_22_port, g => g_vector_0_22_port);
   pg_network_21 : pg_net_210 port map( a => A(21), b => B(21), p => 
                           p_vector_0_21_port, g => g_vector_0_21_port);
   pg_network_20 : pg_net_209 port map( a => A(20), b => B(20), p => 
                           p_vector_0_20_port, g => g_vector_0_20_port);
   pg_network_19 : pg_net_208 port map( a => A(19), b => B(19), p => 
                           p_vector_0_19_port, g => g_vector_0_19_port);
   pg_network_18 : pg_net_207 port map( a => A(18), b => B(18), p => 
                           p_vector_0_18_port, g => g_vector_0_18_port);
   pg_network_17 : pg_net_206 port map( a => A(17), b => B(17), p => 
                           p_vector_0_17_port, g => g_vector_0_17_port);
   pg_network_16 : pg_net_205 port map( a => A(16), b => B(16), p => 
                           p_vector_0_16_port, g => g_vector_0_16_port);
   pg_network_15 : pg_net_204 port map( a => A(15), b => B(15), p => 
                           p_vector_0_15_port, g => g_vector_0_15_port);
   pg_network_14 : pg_net_203 port map( a => A(14), b => B(14), p => 
                           p_vector_0_14_port, g => g_vector_0_14_port);
   pg_network_13 : pg_net_202 port map( a => A(13), b => B(13), p => 
                           p_vector_0_13_port, g => g_vector_0_13_port);
   pg_network_12 : pg_net_201 port map( a => A(12), b => B(12), p => 
                           p_vector_0_12_port, g => g_vector_0_12_port);
   pg_network_11 : pg_net_200 port map( a => A(11), b => B(11), p => 
                           p_vector_0_11_port, g => g_vector_0_11_port);
   pg_network_10 : pg_net_199 port map( a => A(10), b => B(10), p => 
                           p_vector_0_10_port, g => g_vector_0_10_port);
   pg_network_9 : pg_net_198 port map( a => A(9), b => B(9), p => 
                           p_vector_0_9_port, g => g_vector_0_9_port);
   pg_network_8 : pg_net_197 port map( a => A(8), b => B(8), p => 
                           p_vector_0_8_port, g => g_vector_0_8_port);
   pg_network_7 : pg_net_196 port map( a => A(7), b => B(7), p => 
                           p_vector_0_7_port, g => g_vector_0_7_port);
   pg_network_6 : pg_net_195 port map( a => A(6), b => B(6), p => 
                           p_vector_0_6_port, g => g_vector_0_6_port);
   pg_network_5 : pg_net_194 port map( a => A(5), b => B(5), p => 
                           p_vector_0_5_port, g => g_vector_0_5_port);
   pg_network_4 : pg_net_193 port map( a => A(4), b => B(4), p => 
                           p_vector_0_4_port, g => g_vector_0_4_port);
   pg_network_3 : pg_net_192 port map( a => A(3), b => B(3), p => 
                           p_vector_0_3_port, g => g_vector_0_3_port);
   pg_network_2 : pg_net_191 port map( a => A(2), b => B(2), p => 
                           p_vector_0_2_port, g => g_vector_0_2_port);
   pg_network_1 : pg_net_190 port map( a => A(1), b => B(1), p => 
                           p_vector_0_1_port, g => g_vector_0_1_port);
   std_PG_1_31 : PG_BLOCK_216 port map( p2 => p_vector_0_31_port, g2 => 
                           g_vector_0_31_port, p1 => p_vector_0_30_port, g1 => 
                           g_vector_0_30_port, PG_P => p_vector_1_31_port, PG_G
                           => g_vector_1_31_port);
   std_PG_1_29 : PG_BLOCK_215 port map( p2 => p_vector_0_29_port, g2 => 
                           g_vector_0_29_port, p1 => p_vector_0_28_port, g1 => 
                           g_vector_0_28_port, PG_P => p_vector_1_29_port, PG_G
                           => g_vector_1_29_port);
   std_PG_1_27 : PG_BLOCK_214 port map( p2 => p_vector_0_27_port, g2 => 
                           g_vector_0_27_port, p1 => p_vector_0_26_port, g1 => 
                           g_vector_0_26_port, PG_P => p_vector_1_27_port, PG_G
                           => g_vector_1_27_port);
   std_PG_1_25 : PG_BLOCK_213 port map( p2 => p_vector_0_25_port, g2 => 
                           g_vector_0_25_port, p1 => p_vector_0_24_port, g1 => 
                           g_vector_0_24_port, PG_P => p_vector_1_25_port, PG_G
                           => g_vector_1_25_port);
   std_PG_1_23 : PG_BLOCK_212 port map( p2 => p_vector_0_23_port, g2 => 
                           g_vector_0_23_port, p1 => p_vector_0_22_port, g1 => 
                           g_vector_0_22_port, PG_P => p_vector_1_23_port, PG_G
                           => g_vector_1_23_port);
   std_PG_1_21 : PG_BLOCK_211 port map( p2 => p_vector_0_21_port, g2 => 
                           g_vector_0_21_port, p1 => p_vector_0_20_port, g1 => 
                           g_vector_0_20_port, PG_P => p_vector_1_21_port, PG_G
                           => g_vector_1_21_port);
   std_PG_1_19 : PG_BLOCK_210 port map( p2 => p_vector_0_19_port, g2 => 
                           g_vector_0_19_port, p1 => p_vector_0_18_port, g1 => 
                           g_vector_0_18_port, PG_P => p_vector_1_19_port, PG_G
                           => g_vector_1_19_port);
   std_PG_1_17 : PG_BLOCK_209 port map( p2 => p_vector_0_17_port, g2 => 
                           g_vector_0_17_port, p1 => p_vector_0_16_port, g1 => 
                           g_vector_0_16_port, PG_P => p_vector_1_17_port, PG_G
                           => g_vector_1_17_port);
   std_PG_1_15 : PG_BLOCK_208 port map( p2 => p_vector_0_15_port, g2 => 
                           g_vector_0_15_port, p1 => p_vector_0_14_port, g1 => 
                           g_vector_0_14_port, PG_P => p_vector_1_15_port, PG_G
                           => g_vector_1_15_port);
   std_PG_1_13 : PG_BLOCK_207 port map( p2 => p_vector_0_13_port, g2 => 
                           g_vector_0_13_port, p1 => p_vector_0_12_port, g1 => 
                           g_vector_0_12_port, PG_P => p_vector_1_13_port, PG_G
                           => g_vector_1_13_port);
   std_PG_1_11 : PG_BLOCK_206 port map( p2 => p_vector_0_11_port, g2 => 
                           g_vector_0_11_port, p1 => p_vector_0_10_port, g1 => 
                           g_vector_0_10_port, PG_P => p_vector_1_11_port, PG_G
                           => g_vector_1_11_port);
   std_PG_1_9 : PG_BLOCK_205 port map( p2 => p_vector_0_9_port, g2 => 
                           g_vector_0_9_port, p1 => p_vector_0_8_port, g1 => 
                           g_vector_0_8_port, PG_P => p_vector_1_9_port, PG_G 
                           => g_vector_1_9_port);
   std_PG_1_7 : PG_BLOCK_204 port map( p2 => p_vector_0_7_port, g2 => 
                           g_vector_0_7_port, p1 => p_vector_0_6_port, g1 => 
                           g_vector_0_6_port, PG_P => p_vector_1_7_port, PG_G 
                           => g_vector_1_7_port);
   std_PG_1_5 : PG_BLOCK_203 port map( p2 => p_vector_0_5_port, g2 => 
                           g_vector_0_5_port, p1 => p_vector_0_4_port, g1 => 
                           g_vector_0_4_port, PG_P => p_vector_1_5_port, PG_G 
                           => g_vector_1_5_port);
   std_PG_1_3 : PG_BLOCK_202 port map( p2 => p_vector_0_3_port, g2 => 
                           g_vector_0_3_port, p1 => p_vector_0_2_port, g1 => 
                           g_vector_0_2_port, PG_P => p_vector_1_3_port, PG_G 
                           => g_vector_1_3_port);
   std_G_1_1 : G_BLOCK_60 port map( p2 => p_vector_0_1_port, g2 => 
                           g_vector_0_1_port, g1 => g_vector_0_0_port, G => 
                           g_vector_1_1_port);
   std_PG_2_31 : PG_BLOCK_201 port map( p2 => p_vector_1_31_port, g2 => 
                           g_vector_1_31_port, p1 => p_vector_1_29_port, g1 => 
                           g_vector_1_29_port, PG_P => p_vector_2_31_port, PG_G
                           => g_vector_2_31_port);
   std_PG_2_27 : PG_BLOCK_200 port map( p2 => p_vector_1_27_port, g2 => 
                           g_vector_1_27_port, p1 => p_vector_1_25_port, g1 => 
                           g_vector_1_25_port, PG_P => p_vector_2_27_port, PG_G
                           => g_vector_2_27_port);
   std_PG_2_23 : PG_BLOCK_199 port map( p2 => p_vector_1_23_port, g2 => 
                           g_vector_1_23_port, p1 => p_vector_1_21_port, g1 => 
                           g_vector_1_21_port, PG_P => p_vector_2_23_port, PG_G
                           => g_vector_2_23_port);
   std_PG_2_19 : PG_BLOCK_198 port map( p2 => p_vector_1_19_port, g2 => 
                           g_vector_1_19_port, p1 => p_vector_1_17_port, g1 => 
                           g_vector_1_17_port, PG_P => p_vector_2_19_port, PG_G
                           => g_vector_2_19_port);
   std_PG_2_15 : PG_BLOCK_197 port map( p2 => p_vector_1_15_port, g2 => 
                           g_vector_1_15_port, p1 => p_vector_1_13_port, g1 => 
                           g_vector_1_13_port, PG_P => p_vector_2_15_port, PG_G
                           => g_vector_2_15_port);
   std_PG_2_11 : PG_BLOCK_196 port map( p2 => p_vector_1_11_port, g2 => 
                           g_vector_1_11_port, p1 => p_vector_1_9_port, g1 => 
                           g_vector_1_9_port, PG_P => p_vector_2_11_port, PG_G 
                           => g_vector_2_11_port);
   std_PG_2_7 : PG_BLOCK_195 port map( p2 => p_vector_1_7_port, g2 => 
                           g_vector_1_7_port, p1 => p_vector_1_5_port, g1 => 
                           g_vector_1_5_port, PG_P => p_vector_2_7_port, PG_G 
                           => g_vector_2_7_port);
   std_G_2_3 : G_BLOCK_59 port map( p2 => p_vector_1_3_port, g2 => 
                           g_vector_1_3_port, g1 => g_vector_1_1_port, G => 
                           Co_0_port);
   std_PG_3_31 : PG_BLOCK_194 port map( p2 => p_vector_2_31_port, g2 => 
                           g_vector_2_31_port, p1 => p_vector_2_27_port, g1 => 
                           g_vector_2_27_port, PG_P => p_vector_3_31_port, PG_G
                           => g_vector_3_31_port);
   std_PG_3_23 : PG_BLOCK_193 port map( p2 => p_vector_2_23_port, g2 => 
                           g_vector_2_23_port, p1 => p_vector_2_19_port, g1 => 
                           g_vector_2_19_port, PG_P => p_vector_3_23_port, PG_G
                           => g_vector_3_23_port);
   std_PG_3_15 : PG_BLOCK_192 port map( p2 => p_vector_2_15_port, g2 => 
                           g_vector_2_15_port, p1 => p_vector_2_11_port, g1 => 
                           g_vector_2_11_port, PG_P => p_vector_3_15_port, PG_G
                           => g_vector_3_15_port);
   std_G_3_7 : G_BLOCK_58 port map( p2 => p_vector_2_7_port, g2 => 
                           g_vector_2_7_port, g1 => Co_0_port, G => Co_1_port);
   std_PG_4_31 : PG_BLOCK_191 port map( p2 => p_vector_3_31_port, g2 => 
                           g_vector_3_31_port, p1 => p_vector_3_23_port, g1 => 
                           g_vector_3_23_port, PG_P => p_vector_4_31_port, PG_G
                           => g_vector_4_31_port);
   add_PG_4_31_1 : PG_BLOCK_190 port map( p2 => p_vector_2_27_port, g2 => 
                           g_vector_2_27_port, p1 => p_vector_3_23_port, g1 => 
                           g_vector_3_23_port, PG_P => p_vector_4_27_port, PG_G
                           => g_vector_4_27_port);
   std_G_4_15 : G_BLOCK_57 port map( p2 => p_vector_3_15_port, g2 => 
                           g_vector_3_15_port, g1 => Co_1_port, G => Co_3_port)
                           ;
   add_G_4_15_1 : G_BLOCK_56 port map( p2 => p_vector_2_11_port, g2 => 
                           g_vector_2_11_port, g1 => Co_1_port, G => Co_2_port)
                           ;
   std_G_5_31 : G_BLOCK_55 port map( p2 => p_vector_4_31_port, g2 => 
                           g_vector_4_31_port, g1 => Co_3_port, G => Co_7_port)
                           ;
   add_G_5_31_1 : G_BLOCK_54 port map( p2 => p_vector_4_27_port, g2 => 
                           g_vector_4_27_port, g1 => Co_3_port, G => Co_6_port)
                           ;
   add_G_5_31_2 : G_BLOCK_53 port map( p2 => p_vector_3_23_port, g2 => 
                           g_vector_3_23_port, g1 => Co_3_port, G => Co_5_port)
                           ;
   add_G_5_31_3 : G_BLOCK_52 port map( p2 => p_vector_2_19_port, g2 => 
                           g_vector_2_19_port, g1 => Co_3_port, G => Co_4_port)
                           ;
   U1 : OAI21_X1 port map( B1 => n2, B2 => n1, A => n4, ZN => g_vector_0_0_port
                           );
   U2 : INV_X1 port map( A => A(0), ZN => n2);
   U3 : INV_X1 port map( A => B(0), ZN => n1);
   U4 : OAI21_X1 port map( B1 => A(0), B2 => B(0), A => Cin, ZN => n4);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_255 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_255;

architecture SYN_behavioral of my_xor_255 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_254 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_254;

architecture SYN_behavioral of my_xor_254 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_253 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_253;

architecture SYN_behavioral of my_xor_253 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_252 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_252;

architecture SYN_behavioral of my_xor_252 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_251 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_251;

architecture SYN_behavioral of my_xor_251 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_250 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_250;

architecture SYN_behavioral of my_xor_250 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_249 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_249;

architecture SYN_behavioral of my_xor_249 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_248 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_248;

architecture SYN_behavioral of my_xor_248 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_247 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_247;

architecture SYN_behavioral of my_xor_247 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_246 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_246;

architecture SYN_behavioral of my_xor_246 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_245 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_245;

architecture SYN_behavioral of my_xor_245 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_244 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_244;

architecture SYN_behavioral of my_xor_244 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_243 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_243;

architecture SYN_behavioral of my_xor_243 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_242 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_242;

architecture SYN_behavioral of my_xor_242 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_241 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_241;

architecture SYN_behavioral of my_xor_241 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_240 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_240;

architecture SYN_behavioral of my_xor_240 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_239 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_239;

architecture SYN_behavioral of my_xor_239 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_238 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_238;

architecture SYN_behavioral of my_xor_238 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_237 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_237;

architecture SYN_behavioral of my_xor_237 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_236 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_236;

architecture SYN_behavioral of my_xor_236 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_235 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_235;

architecture SYN_behavioral of my_xor_235 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_234 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_234;

architecture SYN_behavioral of my_xor_234 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_233 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_233;

architecture SYN_behavioral of my_xor_233 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_232 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_232;

architecture SYN_behavioral of my_xor_232 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_231 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_231;

architecture SYN_behavioral of my_xor_231 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_230 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_230;

architecture SYN_behavioral of my_xor_230 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_229 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_229;

architecture SYN_behavioral of my_xor_229 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_228 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_228;

architecture SYN_behavioral of my_xor_228 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_227 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_227;

architecture SYN_behavioral of my_xor_227 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_226 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_226;

architecture SYN_behavioral of my_xor_226 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_225 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_225;

architecture SYN_behavioral of my_xor_225 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_224 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_224;

architecture SYN_behavioral of my_xor_224 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_223 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_223;

architecture SYN_behavioral of my_xor_223 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_222 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_222;

architecture SYN_behavioral of my_xor_222 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_221 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_221;

architecture SYN_behavioral of my_xor_221 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_220 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_220;

architecture SYN_behavioral of my_xor_220 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_219 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_219;

architecture SYN_behavioral of my_xor_219 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_218 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_218;

architecture SYN_behavioral of my_xor_218 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_217 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_217;

architecture SYN_behavioral of my_xor_217 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_216 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_216;

architecture SYN_behavioral of my_xor_216 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_215 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_215;

architecture SYN_behavioral of my_xor_215 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_214 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_214;

architecture SYN_behavioral of my_xor_214 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_213 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_213;

architecture SYN_behavioral of my_xor_213 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_212 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_212;

architecture SYN_behavioral of my_xor_212 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_211 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_211;

architecture SYN_behavioral of my_xor_211 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_210 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_210;

architecture SYN_behavioral of my_xor_210 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_209 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_209;

architecture SYN_behavioral of my_xor_209 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_208 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_208;

architecture SYN_behavioral of my_xor_208 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_207 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_207;

architecture SYN_behavioral of my_xor_207 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_206 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_206;

architecture SYN_behavioral of my_xor_206 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_205 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_205;

architecture SYN_behavioral of my_xor_205 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_204 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_204;

architecture SYN_behavioral of my_xor_204 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_203 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_203;

architecture SYN_behavioral of my_xor_203 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_202 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_202;

architecture SYN_behavioral of my_xor_202 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_201 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_201;

architecture SYN_behavioral of my_xor_201 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_200 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_200;

architecture SYN_behavioral of my_xor_200 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_199 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_199;

architecture SYN_behavioral of my_xor_199 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_198 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_198;

architecture SYN_behavioral of my_xor_198 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_197 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_197;

architecture SYN_behavioral of my_xor_197 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_196 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_196;

architecture SYN_behavioral of my_xor_196 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_195 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_195;

architecture SYN_behavioral of my_xor_195 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_194 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_194;

architecture SYN_behavioral of my_xor_194 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_193 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_193;

architecture SYN_behavioral of my_xor_193 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_192 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_192;

architecture SYN_behavioral of my_xor_192 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_191 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_191;

architecture SYN_behavioral of my_xor_191 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_190 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_190;

architecture SYN_behavioral of my_xor_190 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_189 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_189;

architecture SYN_behavioral of my_xor_189 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_188 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_188;

architecture SYN_behavioral of my_xor_188 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_187 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_187;

architecture SYN_behavioral of my_xor_187 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_186 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_186;

architecture SYN_behavioral of my_xor_186 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_185 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_185;

architecture SYN_behavioral of my_xor_185 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_184 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_184;

architecture SYN_behavioral of my_xor_184 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_183 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_183;

architecture SYN_behavioral of my_xor_183 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_182 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_182;

architecture SYN_behavioral of my_xor_182 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_181 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_181;

architecture SYN_behavioral of my_xor_181 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_180 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_180;

architecture SYN_behavioral of my_xor_180 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_179 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_179;

architecture SYN_behavioral of my_xor_179 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_178 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_178;

architecture SYN_behavioral of my_xor_178 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_177 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_177;

architecture SYN_behavioral of my_xor_177 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_176 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_176;

architecture SYN_behavioral of my_xor_176 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_175 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_175;

architecture SYN_behavioral of my_xor_175 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_174 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_174;

architecture SYN_behavioral of my_xor_174 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_173 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_173;

architecture SYN_behavioral of my_xor_173 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_172 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_172;

architecture SYN_behavioral of my_xor_172 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_171 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_171;

architecture SYN_behavioral of my_xor_171 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_170 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_170;

architecture SYN_behavioral of my_xor_170 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_169 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_169;

architecture SYN_behavioral of my_xor_169 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_168 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_168;

architecture SYN_behavioral of my_xor_168 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_167 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_167;

architecture SYN_behavioral of my_xor_167 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_166 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_166;

architecture SYN_behavioral of my_xor_166 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_165 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_165;

architecture SYN_behavioral of my_xor_165 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_164 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_164;

architecture SYN_behavioral of my_xor_164 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_163 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_163;

architecture SYN_behavioral of my_xor_163 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_162 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_162;

architecture SYN_behavioral of my_xor_162 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_161 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_161;

architecture SYN_behavioral of my_xor_161 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_160 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_160;

architecture SYN_behavioral of my_xor_160 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_159 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_159;

architecture SYN_behavioral of my_xor_159 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_158 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_158;

architecture SYN_behavioral of my_xor_158 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_157 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_157;

architecture SYN_behavioral of my_xor_157 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_156 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_156;

architecture SYN_behavioral of my_xor_156 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_155 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_155;

architecture SYN_behavioral of my_xor_155 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_154 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_154;

architecture SYN_behavioral of my_xor_154 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_153 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_153;

architecture SYN_behavioral of my_xor_153 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_152 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_152;

architecture SYN_behavioral of my_xor_152 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_151 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_151;

architecture SYN_behavioral of my_xor_151 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_150 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_150;

architecture SYN_behavioral of my_xor_150 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_149 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_149;

architecture SYN_behavioral of my_xor_149 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_148 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_148;

architecture SYN_behavioral of my_xor_148 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_147 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_147;

architecture SYN_behavioral of my_xor_147 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_146 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_146;

architecture SYN_behavioral of my_xor_146 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_145 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_145;

architecture SYN_behavioral of my_xor_145 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_144 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_144;

architecture SYN_behavioral of my_xor_144 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_143 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_143;

architecture SYN_behavioral of my_xor_143 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_142 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_142;

architecture SYN_behavioral of my_xor_142 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_141 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_141;

architecture SYN_behavioral of my_xor_141 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_140 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_140;

architecture SYN_behavioral of my_xor_140 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_139 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_139;

architecture SYN_behavioral of my_xor_139 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_138 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_138;

architecture SYN_behavioral of my_xor_138 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_137 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_137;

architecture SYN_behavioral of my_xor_137 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_136 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_136;

architecture SYN_behavioral of my_xor_136 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_135 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_135;

architecture SYN_behavioral of my_xor_135 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_134 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_134;

architecture SYN_behavioral of my_xor_134 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_133 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_133;

architecture SYN_behavioral of my_xor_133 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_132 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_132;

architecture SYN_behavioral of my_xor_132 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_131 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_131;

architecture SYN_behavioral of my_xor_131 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_130 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_130;

architecture SYN_behavioral of my_xor_130 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_129 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_129;

architecture SYN_behavioral of my_xor_129 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_128 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_128;

architecture SYN_behavioral of my_xor_128 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_127 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_127;

architecture SYN_behavioral_architecture of my_xor_127 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_126 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_126;

architecture SYN_behavioral_architecture2 of my_xor_126 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_125 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_125;

architecture SYN_behavioral_architecture3 of my_xor_125 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_124 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_124;

architecture SYN_behavioral_architecture4 of my_xor_124 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_123 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_123;

architecture SYN_behavioral_architecture5 of my_xor_123 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture5;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_122 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_122;

architecture SYN_behavioral_architecture6 of my_xor_122 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture6;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_121 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_121;

architecture SYN_behavioral_architecture7 of my_xor_121 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture7;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_120 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_120;

architecture SYN_behavioral_architecture8 of my_xor_120 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture8;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_119 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_119;

architecture SYN_behavioral_architecture9 of my_xor_119 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture9;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_118 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_118;

architecture SYN_behavioral_architecture10 of my_xor_118 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture10;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_117 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_117;

architecture SYN_behavioral_architecture11 of my_xor_117 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture11;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_116 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_116;

architecture SYN_behavioral_architecture12 of my_xor_116 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture12;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_115 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_115;

architecture SYN_behavioral_architecture13 of my_xor_115 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture13;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_114 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_114;

architecture SYN_behavioral_architecture14 of my_xor_114 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture14;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_113 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_113;

architecture SYN_behavioral_architecture15 of my_xor_113 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture15;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_112 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_112;

architecture SYN_behavioral_architecture16 of my_xor_112 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture16;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_111 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_111;

architecture SYN_behavioral_architecture17 of my_xor_111 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture17;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_110 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_110;

architecture SYN_behavioral_architecture18 of my_xor_110 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture18;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_109 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_109;

architecture SYN_behavioral_architecture19 of my_xor_109 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture19;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_108 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_108;

architecture SYN_behavioral_architecture20 of my_xor_108 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture20;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_107 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_107;

architecture SYN_behavioral_architecture21 of my_xor_107 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture21;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_106 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_106;

architecture SYN_behavioral_architecture22 of my_xor_106 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture22;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_105 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_105;

architecture SYN_behavioral_architecture23 of my_xor_105 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture23;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_104 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_104;

architecture SYN_behavioral_architecture24 of my_xor_104 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture24;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_103 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_103;

architecture SYN_behavioral_architecture25 of my_xor_103 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture25;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_102 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_102;

architecture SYN_behavioral_architecture26 of my_xor_102 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture26;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_101 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_101;

architecture SYN_behavioral_architecture27 of my_xor_101 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture27;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_100 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_100;

architecture SYN_behavioral_architecture28 of my_xor_100 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture28;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_99 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_99;

architecture SYN_behavioral_architecture29 of my_xor_99 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture29;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_98 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_98;

architecture SYN_behavioral_architecture30 of my_xor_98 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture30;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_97 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_97;

architecture SYN_behavioral_architecture31 of my_xor_97 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture31;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_96 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_96;

architecture SYN_behavioral_architecture32 of my_xor_96 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture32;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_95 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_95;

architecture SYN_behavioral_architecture33 of my_xor_95 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture33;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_94 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_94;

architecture SYN_behavioral_architecture34 of my_xor_94 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture34;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_93 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_93;

architecture SYN_behavioral_architecture35 of my_xor_93 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture35;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_92 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_92;

architecture SYN_behavioral_architecture36 of my_xor_92 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture36;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_91 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_91;

architecture SYN_behavioral_architecture37 of my_xor_91 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture37;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_90 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_90;

architecture SYN_behavioral_architecture38 of my_xor_90 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture38;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_89 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_89;

architecture SYN_behavioral_architecture39 of my_xor_89 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture39;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_88 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_88;

architecture SYN_behavioral_architecture40 of my_xor_88 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture40;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_87 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_87;

architecture SYN_behavioral_architecture41 of my_xor_87 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture41;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_86 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_86;

architecture SYN_behavioral_architecture42 of my_xor_86 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture42;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_85 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_85;

architecture SYN_behavioral_architecture43 of my_xor_85 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture43;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_84 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_84;

architecture SYN_behavioral_architecture44 of my_xor_84 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture44;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_83 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_83;

architecture SYN_behavioral_architecture45 of my_xor_83 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture45;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_82 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_82;

architecture SYN_behavioral_architecture46 of my_xor_82 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture46;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_81 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_81;

architecture SYN_behavioral_architecture47 of my_xor_81 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture47;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_80 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_80;

architecture SYN_behavioral_architecture48 of my_xor_80 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture48;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_79 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_79;

architecture SYN_behavioral_architecture49 of my_xor_79 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture49;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_78 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_78;

architecture SYN_behavioral_architecture50 of my_xor_78 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture50;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_77 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_77;

architecture SYN_behavioral_architecture51 of my_xor_77 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture51;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_76 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_76;

architecture SYN_behavioral_architecture52 of my_xor_76 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture52;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_75 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_75;

architecture SYN_behavioral_architecture53 of my_xor_75 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture53;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_74 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_74;

architecture SYN_behavioral_architecture54 of my_xor_74 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture54;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_73 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_73;

architecture SYN_behavioral_architecture55 of my_xor_73 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture55;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_72 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_72;

architecture SYN_behavioral_architecture56 of my_xor_72 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture56;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_71 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_71;

architecture SYN_behavioral_architecture57 of my_xor_71 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture57;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_70 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_70;

architecture SYN_behavioral_architecture58 of my_xor_70 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture58;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_69 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_69;

architecture SYN_behavioral_architecture59 of my_xor_69 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture59;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_68 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_68;

architecture SYN_behavioral_architecture60 of my_xor_68 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture60;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_67 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_67;

architecture SYN_behavioral_architecture61 of my_xor_67 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture61;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_66 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_66;

architecture SYN_behavioral_architecture62 of my_xor_66 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture62;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_65 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_65;

architecture SYN_behavioral_architecture63 of my_xor_65 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture63;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_64 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_64;

architecture SYN_behavioral of my_xor_64 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_63 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_63;

architecture SYN_behavioral_architecture of my_xor_63 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_62 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_62;

architecture SYN_behavioral_architecture2 of my_xor_62 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_61 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_61;

architecture SYN_behavioral_architecture3 of my_xor_61 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_60 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_60;

architecture SYN_behavioral_architecture4 of my_xor_60 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_59 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_59;

architecture SYN_behavioral_architecture5 of my_xor_59 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture5;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_58 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_58;

architecture SYN_behavioral_architecture6 of my_xor_58 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture6;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_57 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_57;

architecture SYN_behavioral_architecture7 of my_xor_57 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture7;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_56 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_56;

architecture SYN_behavioral_architecture8 of my_xor_56 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture8;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_55 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_55;

architecture SYN_behavioral_architecture9 of my_xor_55 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture9;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_54 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_54;

architecture SYN_behavioral_architecture10 of my_xor_54 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture10;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_53 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_53;

architecture SYN_behavioral_architecture11 of my_xor_53 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture11;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_52 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_52;

architecture SYN_behavioral_architecture12 of my_xor_52 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture12;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_51 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_51;

architecture SYN_behavioral_architecture13 of my_xor_51 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture13;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_50 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_50;

architecture SYN_behavioral_architecture14 of my_xor_50 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture14;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_49 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_49;

architecture SYN_behavioral_architecture15 of my_xor_49 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture15;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_48 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_48;

architecture SYN_behavioral_architecture16 of my_xor_48 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture16;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_47 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_47;

architecture SYN_behavioral_architecture17 of my_xor_47 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture17;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_46 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_46;

architecture SYN_behavioral_architecture18 of my_xor_46 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture18;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_45 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_45;

architecture SYN_behavioral_architecture19 of my_xor_45 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture19;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_44 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_44;

architecture SYN_behavioral_architecture20 of my_xor_44 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture20;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_43 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_43;

architecture SYN_behavioral_architecture21 of my_xor_43 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture21;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_42 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_42;

architecture SYN_behavioral_architecture22 of my_xor_42 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture22;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_41 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_41;

architecture SYN_behavioral_architecture23 of my_xor_41 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture23;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_40 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_40;

architecture SYN_behavioral_architecture24 of my_xor_40 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture24;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_39 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_39;

architecture SYN_behavioral_architecture25 of my_xor_39 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture25;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_38 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_38;

architecture SYN_behavioral_architecture26 of my_xor_38 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture26;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_37 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_37;

architecture SYN_behavioral_architecture27 of my_xor_37 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture27;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_36 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_36;

architecture SYN_behavioral_architecture28 of my_xor_36 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture28;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_35 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_35;

architecture SYN_behavioral_architecture29 of my_xor_35 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture29;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_34 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_34;

architecture SYN_behavioral_architecture30 of my_xor_34 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture30;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_33 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_33;

architecture SYN_behavioral_architecture31 of my_xor_33 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture31;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_32 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_32;

architecture SYN_behavioral_architecture32 of my_xor_32 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture32;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_31 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_31;

architecture SYN_behavioral_architecture33 of my_xor_31 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture33;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_30 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_30;

architecture SYN_behavioral_architecture34 of my_xor_30 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture34;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_29 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_29;

architecture SYN_behavioral_architecture35 of my_xor_29 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture35;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_28 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_28;

architecture SYN_behavioral_architecture36 of my_xor_28 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture36;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_27 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_27;

architecture SYN_behavioral_architecture37 of my_xor_27 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture37;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_26 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_26;

architecture SYN_behavioral_architecture38 of my_xor_26 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture38;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_25 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_25;

architecture SYN_behavioral_architecture39 of my_xor_25 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture39;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_24 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_24;

architecture SYN_behavioral_architecture40 of my_xor_24 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture40;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_23 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_23;

architecture SYN_behavioral_architecture41 of my_xor_23 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture41;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_22 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_22;

architecture SYN_behavioral_architecture42 of my_xor_22 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture42;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_21 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_21;

architecture SYN_behavioral_architecture43 of my_xor_21 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture43;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_20 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_20;

architecture SYN_behavioral_architecture44 of my_xor_20 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture44;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_19 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_19;

architecture SYN_behavioral_architecture45 of my_xor_19 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture45;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_18 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_18;

architecture SYN_behavioral_architecture46 of my_xor_18 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture46;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_17 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_17;

architecture SYN_behavioral_architecture47 of my_xor_17 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture47;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_16 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_16;

architecture SYN_behavioral_architecture48 of my_xor_16 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture48;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_15 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_15;

architecture SYN_behavioral_architecture49 of my_xor_15 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture49;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_14 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_14;

architecture SYN_behavioral_architecture50 of my_xor_14 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture50;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_13 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_13;

architecture SYN_behavioral_architecture51 of my_xor_13 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture51;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_12 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_12;

architecture SYN_behavioral_architecture52 of my_xor_12 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture52;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_11 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_11;

architecture SYN_behavioral_architecture53 of my_xor_11 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture53;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_10 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_10;

architecture SYN_behavioral_architecture54 of my_xor_10 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture54;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_9 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_9;

architecture SYN_behavioral_architecture55 of my_xor_9 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture55;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_8 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_8;

architecture SYN_behavioral_architecture56 of my_xor_8 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture56;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_7 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_7;

architecture SYN_behavioral_architecture57 of my_xor_7 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture57;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_6 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_6;

architecture SYN_behavioral_architecture58 of my_xor_6 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture58;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_5 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_5;

architecture SYN_behavioral_architecture59 of my_xor_5 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture59;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_4 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_4;

architecture SYN_behavioral_architecture60 of my_xor_4 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture60;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_3 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_3;

architecture SYN_behavioral_architecture61 of my_xor_3 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture61;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_2 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_2;

architecture SYN_behavioral_architecture62 of my_xor_2 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture62;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_1 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_1;

architecture SYN_behavioral_architecture63 of my_xor_1 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral_architecture63;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT5_1 is

   port( A, B : in std_logic_vector (4 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (4 downto 0));

end MUX21_GENERIC_NBIT5_1;

architecture SYN_structural of MUX21_GENERIC_NBIT5_1 is

   component MUX21_457
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_458
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_459
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_460
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_461
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_461 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_460 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_459 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_458 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));
   MUXES_4 : MUX21_457 port map( A => A(4), B => B(4), S => SEL, Y => Y(4));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_GENERIC_NBIT32_2 is

   port( A, B, C, D : in std_logic_vector (31 downto 0);  SEL : in 
         std_logic_vector (1 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end MUX41_GENERIC_NBIT32_2;

architecture SYN_structural of MUX41_GENERIC_NBIT32_2 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX41_105
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_106
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_107
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_108
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_109
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_110
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_111
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_112
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_113
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_114
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_115
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_116
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_117
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_118
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_119
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_120
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_121
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_122
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_123
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_124
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_125
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_126
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_127
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_128
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_129
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_130
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_131
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_132
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_133
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_134
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_135
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_136
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   MUXES_0 : MUX41_136 port map( A => A(0), B => B(0), C => C(0), D => D(0), 
                           S(1) => n4, S(0) => n1, Y => Y(0));
   MUXES_1 : MUX41_135 port map( A => A(1), B => B(1), C => C(1), D => D(1), 
                           S(1) => n4, S(0) => n1, Y => Y(1));
   MUXES_2 : MUX41_134 port map( A => A(2), B => B(2), C => C(2), D => D(2), 
                           S(1) => n4, S(0) => n1, Y => Y(2));
   MUXES_3 : MUX41_133 port map( A => A(3), B => B(3), C => C(3), D => D(3), 
                           S(1) => n4, S(0) => n1, Y => Y(3));
   MUXES_4 : MUX41_132 port map( A => A(4), B => B(4), C => C(4), D => D(4), 
                           S(1) => n4, S(0) => n1, Y => Y(4));
   MUXES_5 : MUX41_131 port map( A => A(5), B => B(5), C => C(5), D => D(5), 
                           S(1) => n4, S(0) => n1, Y => Y(5));
   MUXES_6 : MUX41_130 port map( A => A(6), B => B(6), C => C(6), D => D(6), 
                           S(1) => n4, S(0) => n1, Y => Y(6));
   MUXES_7 : MUX41_129 port map( A => A(7), B => B(7), C => C(7), D => D(7), 
                           S(1) => n4, S(0) => n1, Y => Y(7));
   MUXES_8 : MUX41_128 port map( A => A(8), B => B(8), C => C(8), D => D(8), 
                           S(1) => n4, S(0) => n1, Y => Y(8));
   MUXES_9 : MUX41_127 port map( A => A(9), B => B(9), C => C(9), D => D(9), 
                           S(1) => n4, S(0) => n1, Y => Y(9));
   MUXES_10 : MUX41_126 port map( A => A(10), B => B(10), C => C(10), D => 
                           D(10), S(1) => n4, S(0) => n1, Y => Y(10));
   MUXES_11 : MUX41_125 port map( A => A(11), B => B(11), C => C(11), D => 
                           D(11), S(1) => n4, S(0) => n2, Y => Y(11));
   MUXES_12 : MUX41_124 port map( A => A(12), B => B(12), C => C(12), D => 
                           D(12), S(1) => n5, S(0) => n2, Y => Y(12));
   MUXES_13 : MUX41_123 port map( A => A(13), B => B(13), C => C(13), D => 
                           D(13), S(1) => n5, S(0) => n2, Y => Y(13));
   MUXES_14 : MUX41_122 port map( A => A(14), B => B(14), C => C(14), D => 
                           D(14), S(1) => n5, S(0) => n2, Y => Y(14));
   MUXES_15 : MUX41_121 port map( A => A(15), B => B(15), C => C(15), D => 
                           D(15), S(1) => n5, S(0) => n2, Y => Y(15));
   MUXES_16 : MUX41_120 port map( A => A(16), B => B(16), C => C(16), D => 
                           D(16), S(1) => n5, S(0) => n2, Y => Y(16));
   MUXES_17 : MUX41_119 port map( A => A(17), B => B(17), C => C(17), D => 
                           D(17), S(1) => n5, S(0) => n2, Y => Y(17));
   MUXES_18 : MUX41_118 port map( A => A(18), B => B(18), C => C(18), D => 
                           D(18), S(1) => n5, S(0) => n2, Y => Y(18));
   MUXES_19 : MUX41_117 port map( A => A(19), B => B(19), C => C(19), D => 
                           D(19), S(1) => n5, S(0) => n2, Y => Y(19));
   MUXES_20 : MUX41_116 port map( A => A(20), B => B(20), C => C(20), D => 
                           D(20), S(1) => n5, S(0) => n2, Y => Y(20));
   MUXES_21 : MUX41_115 port map( A => A(21), B => B(21), C => C(21), D => 
                           D(21), S(1) => n5, S(0) => n2, Y => Y(21));
   MUXES_22 : MUX41_114 port map( A => A(22), B => B(22), C => C(22), D => 
                           D(22), S(1) => n5, S(0) => n3, Y => Y(22));
   MUXES_23 : MUX41_113 port map( A => A(23), B => B(23), C => C(23), D => 
                           D(23), S(1) => n5, S(0) => n3, Y => Y(23));
   MUXES_24 : MUX41_112 port map( A => A(24), B => B(24), C => C(24), D => 
                           D(24), S(1) => n6, S(0) => n3, Y => Y(24));
   MUXES_25 : MUX41_111 port map( A => A(25), B => B(25), C => C(25), D => 
                           D(25), S(1) => n6, S(0) => n3, Y => Y(25));
   MUXES_26 : MUX41_110 port map( A => A(26), B => B(26), C => C(26), D => 
                           D(26), S(1) => n6, S(0) => n3, Y => Y(26));
   MUXES_27 : MUX41_109 port map( A => A(27), B => B(27), C => C(27), D => 
                           D(27), S(1) => n6, S(0) => n3, Y => Y(27));
   MUXES_28 : MUX41_108 port map( A => A(28), B => B(28), C => C(28), D => 
                           D(28), S(1) => n6, S(0) => n3, Y => Y(28));
   MUXES_29 : MUX41_107 port map( A => A(29), B => B(29), C => C(29), D => 
                           D(29), S(1) => n6, S(0) => n3, Y => Y(29));
   MUXES_30 : MUX41_106 port map( A => A(30), B => B(30), C => C(30), D => 
                           D(30), S(1) => n6, S(0) => n3, Y => Y(30));
   MUXES_31 : MUX41_105 port map( A => A(31), B => B(31), C => C(31), D => 
                           D(31), S(1) => n6, S(0) => n3, Y => Y(31));
   U1 : BUF_X1 port map( A => SEL(1), Z => n5);
   U2 : BUF_X1 port map( A => SEL(1), Z => n4);
   U3 : BUF_X1 port map( A => SEL(1), Z => n6);
   U4 : BUF_X1 port map( A => SEL(0), Z => n2);
   U5 : BUF_X1 port map( A => SEL(0), Z => n1);
   U6 : BUF_X1 port map( A => SEL(0), Z => n3);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_GENERIC_NBIT32_1 is

   port( A, B, C, D : in std_logic_vector (31 downto 0);  SEL : in 
         std_logic_vector (1 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end MUX41_GENERIC_NBIT32_1;

architecture SYN_structural of MUX41_GENERIC_NBIT32_1 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX41_73
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_74
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_75
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_76
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_77
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_78
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_79
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_80
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_81
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_82
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_83
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_84
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_85
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_86
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_87
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_88
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_89
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_90
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_91
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_92
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_93
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_94
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_95
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_96
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_97
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_98
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_99
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_100
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_101
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_102
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_103
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_104
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   MUXES_0 : MUX41_104 port map( A => A(0), B => B(0), C => C(0), D => D(0), 
                           S(1) => n4, S(0) => n1, Y => Y(0));
   MUXES_1 : MUX41_103 port map( A => A(1), B => B(1), C => C(1), D => D(1), 
                           S(1) => n4, S(0) => n1, Y => Y(1));
   MUXES_2 : MUX41_102 port map( A => A(2), B => B(2), C => C(2), D => D(2), 
                           S(1) => n4, S(0) => n1, Y => Y(2));
   MUXES_3 : MUX41_101 port map( A => A(3), B => B(3), C => C(3), D => D(3), 
                           S(1) => n4, S(0) => n1, Y => Y(3));
   MUXES_4 : MUX41_100 port map( A => A(4), B => B(4), C => C(4), D => D(4), 
                           S(1) => n4, S(0) => n1, Y => Y(4));
   MUXES_5 : MUX41_99 port map( A => A(5), B => B(5), C => C(5), D => D(5), 
                           S(1) => n4, S(0) => n1, Y => Y(5));
   MUXES_6 : MUX41_98 port map( A => A(6), B => B(6), C => C(6), D => D(6), 
                           S(1) => n4, S(0) => n1, Y => Y(6));
   MUXES_7 : MUX41_97 port map( A => A(7), B => B(7), C => C(7), D => D(7), 
                           S(1) => n4, S(0) => n1, Y => Y(7));
   MUXES_8 : MUX41_96 port map( A => A(8), B => B(8), C => C(8), D => D(8), 
                           S(1) => n4, S(0) => n1, Y => Y(8));
   MUXES_9 : MUX41_95 port map( A => A(9), B => B(9), C => C(9), D => D(9), 
                           S(1) => n4, S(0) => n1, Y => Y(9));
   MUXES_10 : MUX41_94 port map( A => A(10), B => B(10), C => C(10), D => D(10)
                           , S(1) => n4, S(0) => n1, Y => Y(10));
   MUXES_11 : MUX41_93 port map( A => A(11), B => B(11), C => C(11), D => D(11)
                           , S(1) => n4, S(0) => n2, Y => Y(11));
   MUXES_12 : MUX41_92 port map( A => A(12), B => B(12), C => C(12), D => D(12)
                           , S(1) => n5, S(0) => n2, Y => Y(12));
   MUXES_13 : MUX41_91 port map( A => A(13), B => B(13), C => C(13), D => D(13)
                           , S(1) => n5, S(0) => n2, Y => Y(13));
   MUXES_14 : MUX41_90 port map( A => A(14), B => B(14), C => C(14), D => D(14)
                           , S(1) => n5, S(0) => n2, Y => Y(14));
   MUXES_15 : MUX41_89 port map( A => A(15), B => B(15), C => C(15), D => D(15)
                           , S(1) => n5, S(0) => n2, Y => Y(15));
   MUXES_16 : MUX41_88 port map( A => A(16), B => B(16), C => C(16), D => D(16)
                           , S(1) => n5, S(0) => n2, Y => Y(16));
   MUXES_17 : MUX41_87 port map( A => A(17), B => B(17), C => C(17), D => D(17)
                           , S(1) => n5, S(0) => n2, Y => Y(17));
   MUXES_18 : MUX41_86 port map( A => A(18), B => B(18), C => C(18), D => D(18)
                           , S(1) => n5, S(0) => n2, Y => Y(18));
   MUXES_19 : MUX41_85 port map( A => A(19), B => B(19), C => C(19), D => D(19)
                           , S(1) => n5, S(0) => n2, Y => Y(19));
   MUXES_20 : MUX41_84 port map( A => A(20), B => B(20), C => C(20), D => D(20)
                           , S(1) => n5, S(0) => n2, Y => Y(20));
   MUXES_21 : MUX41_83 port map( A => A(21), B => B(21), C => C(21), D => D(21)
                           , S(1) => n5, S(0) => n2, Y => Y(21));
   MUXES_22 : MUX41_82 port map( A => A(22), B => B(22), C => C(22), D => D(22)
                           , S(1) => n5, S(0) => n3, Y => Y(22));
   MUXES_23 : MUX41_81 port map( A => A(23), B => B(23), C => C(23), D => D(23)
                           , S(1) => n5, S(0) => n3, Y => Y(23));
   MUXES_24 : MUX41_80 port map( A => A(24), B => B(24), C => C(24), D => D(24)
                           , S(1) => n6, S(0) => n3, Y => Y(24));
   MUXES_25 : MUX41_79 port map( A => A(25), B => B(25), C => C(25), D => D(25)
                           , S(1) => n6, S(0) => n3, Y => Y(25));
   MUXES_26 : MUX41_78 port map( A => A(26), B => B(26), C => C(26), D => D(26)
                           , S(1) => n6, S(0) => n3, Y => Y(26));
   MUXES_27 : MUX41_77 port map( A => A(27), B => B(27), C => C(27), D => D(27)
                           , S(1) => n6, S(0) => n3, Y => Y(27));
   MUXES_28 : MUX41_76 port map( A => A(28), B => B(28), C => C(28), D => D(28)
                           , S(1) => n6, S(0) => n3, Y => Y(28));
   MUXES_29 : MUX41_75 port map( A => A(29), B => B(29), C => C(29), D => D(29)
                           , S(1) => n6, S(0) => n3, Y => Y(29));
   MUXES_30 : MUX41_74 port map( A => A(30), B => B(30), C => C(30), D => D(30)
                           , S(1) => n6, S(0) => n3, Y => Y(30));
   MUXES_31 : MUX41_73 port map( A => A(31), B => B(31), C => C(31), D => D(31)
                           , S(1) => n6, S(0) => n3, Y => Y(31));
   U1 : BUF_X1 port map( A => SEL(1), Z => n5);
   U2 : BUF_X1 port map( A => SEL(1), Z => n4);
   U3 : BUF_X1 port map( A => SEL(1), Z => n6);
   U4 : BUF_X1 port map( A => SEL(0), Z => n2);
   U5 : BUF_X1 port map( A => SEL(0), Z => n1);
   U6 : BUF_X1 port map( A => SEL(0), Z => n3);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity P4_ADDER_NBIT32_1 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  S : 
         out std_logic_vector (31 downto 0);  Cout, ovf : out std_logic);

end P4_ADDER_NBIT32_1;

architecture SYN_STRUCTURAL of P4_ADDER_NBIT32_1 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component sum_generator_n_bit32_n_CSB8_1
      port( A, B : in std_logic_vector (31 downto 0);  C_in : in 
            std_logic_vector (7 downto 0);  S : out std_logic_vector (31 downto
            0));
   end component;
   
   component CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_1
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co 
            : out std_logic_vector (7 downto 0));
   end component;
   
   component my_xor_193
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_194
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_195
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_196
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_197
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_198
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_199
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_200
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_201
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_202
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_203
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_204
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_205
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_206
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_207
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_208
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_209
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_210
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_211
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_212
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_213
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_214
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_215
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_216
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_217
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_218
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_219
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_220
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_221
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_222
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_223
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_224
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal S_31_port, S_30_port, S_29_port, S_28_port, S_27_port, S_26_port, 
      S_25_port, S_24_port, S_23_port, S_22_port, S_21_port, S_20_port, 
      S_19_port, S_18_port, S_17_port, S_16_port, S_15_port, S_14_port, 
      S_13_port, S_12_port, S_11_port, S_10_port, S_9_port, S_8_port, S_7_port,
      S_6_port, S_5_port, S_4_port, S_3_port, S_2_port, S_1_port, S_0_port, 
      xor_b_31_port, xor_b_30_port, xor_b_29_port, xor_b_28_port, xor_b_27_port
      , xor_b_26_port, xor_b_25_port, xor_b_24_port, xor_b_23_port, 
      xor_b_22_port, xor_b_21_port, xor_b_20_port, xor_b_19_port, xor_b_18_port
      , xor_b_17_port, xor_b_16_port, xor_b_15_port, xor_b_14_port, 
      xor_b_13_port, xor_b_12_port, xor_b_11_port, xor_b_10_port, xor_b_9_port,
      xor_b_8_port, xor_b_7_port, xor_b_6_port, xor_b_5_port, xor_b_4_port, 
      xor_b_3_port, xor_b_2_port, xor_b_1_port, xor_b_0_port, carry_6_port, 
      carry_5_port, carry_4_port, carry_3_port, carry_2_port, carry_1_port, 
      carry_0_port, n3, n4, n5, n6 : std_logic;

begin
   S <= ( S_31_port, S_30_port, S_29_port, S_28_port, S_27_port, S_26_port, 
      S_25_port, S_24_port, S_23_port, S_22_port, S_21_port, S_20_port, 
      S_19_port, S_18_port, S_17_port, S_16_port, S_15_port, S_14_port, 
      S_13_port, S_12_port, S_11_port, S_10_port, S_9_port, S_8_port, S_7_port,
      S_6_port, S_5_port, S_4_port, S_3_port, S_2_port, S_1_port, S_0_port );
   
   U3 : XOR2_X1 port map( A => xor_b_31_port, B => A(31), Z => n5);
   bc_xor_31 : my_xor_224 port map( A => B(31), B => n3, xor_out => 
                           xor_b_31_port);
   bc_xor_30 : my_xor_223 port map( A => B(30), B => n3, xor_out => 
                           xor_b_30_port);
   bc_xor_29 : my_xor_222 port map( A => B(29), B => n3, xor_out => 
                           xor_b_29_port);
   bc_xor_28 : my_xor_221 port map( A => B(28), B => n3, xor_out => 
                           xor_b_28_port);
   bc_xor_27 : my_xor_220 port map( A => B(27), B => n3, xor_out => 
                           xor_b_27_port);
   bc_xor_26 : my_xor_219 port map( A => B(26), B => n3, xor_out => 
                           xor_b_26_port);
   bc_xor_25 : my_xor_218 port map( A => B(25), B => n3, xor_out => 
                           xor_b_25_port);
   bc_xor_24 : my_xor_217 port map( A => B(24), B => n3, xor_out => 
                           xor_b_24_port);
   bc_xor_23 : my_xor_216 port map( A => B(23), B => n3, xor_out => 
                           xor_b_23_port);
   bc_xor_22 : my_xor_215 port map( A => B(22), B => n3, xor_out => 
                           xor_b_22_port);
   bc_xor_21 : my_xor_214 port map( A => B(21), B => n3, xor_out => 
                           xor_b_21_port);
   bc_xor_20 : my_xor_213 port map( A => B(20), B => n3, xor_out => 
                           xor_b_20_port);
   bc_xor_19 : my_xor_212 port map( A => B(19), B => n3, xor_out => 
                           xor_b_19_port);
   bc_xor_18 : my_xor_211 port map( A => B(18), B => n3, xor_out => 
                           xor_b_18_port);
   bc_xor_17 : my_xor_210 port map( A => B(17), B => n3, xor_out => 
                           xor_b_17_port);
   bc_xor_16 : my_xor_209 port map( A => B(16), B => n4, xor_out => 
                           xor_b_16_port);
   bc_xor_15 : my_xor_208 port map( A => B(15), B => n4, xor_out => 
                           xor_b_15_port);
   bc_xor_14 : my_xor_207 port map( A => B(14), B => n4, xor_out => 
                           xor_b_14_port);
   bc_xor_13 : my_xor_206 port map( A => B(13), B => n4, xor_out => 
                           xor_b_13_port);
   bc_xor_12 : my_xor_205 port map( A => B(12), B => n4, xor_out => 
                           xor_b_12_port);
   bc_xor_11 : my_xor_204 port map( A => B(11), B => n4, xor_out => 
                           xor_b_11_port);
   bc_xor_10 : my_xor_203 port map( A => B(10), B => n4, xor_out => 
                           xor_b_10_port);
   bc_xor_9 : my_xor_202 port map( A => B(9), B => n4, xor_out => xor_b_9_port)
                           ;
   bc_xor_8 : my_xor_201 port map( A => B(8), B => n4, xor_out => xor_b_8_port)
                           ;
   bc_xor_7 : my_xor_200 port map( A => B(7), B => n4, xor_out => xor_b_7_port)
                           ;
   bc_xor_6 : my_xor_199 port map( A => B(6), B => n4, xor_out => xor_b_6_port)
                           ;
   bc_xor_5 : my_xor_198 port map( A => B(5), B => n4, xor_out => xor_b_5_port)
                           ;
   bc_xor_4 : my_xor_197 port map( A => B(4), B => n4, xor_out => xor_b_4_port)
                           ;
   bc_xor_3 : my_xor_196 port map( A => B(3), B => n4, xor_out => xor_b_3_port)
                           ;
   bc_xor_2 : my_xor_195 port map( A => B(2), B => n4, xor_out => xor_b_2_port)
                           ;
   bc_xor_1 : my_xor_194 port map( A => B(1), B => n4, xor_out => xor_b_1_port)
                           ;
   bc_xor_0 : my_xor_193 port map( A => B(0), B => n4, xor_out => xor_b_0_port)
                           ;
   CG : CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_1 port map( A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(31) => 
                           xor_b_31_port, B(30) => xor_b_30_port, B(29) => 
                           xor_b_29_port, B(28) => xor_b_28_port, B(27) => 
                           xor_b_27_port, B(26) => xor_b_26_port, B(25) => 
                           xor_b_25_port, B(24) => xor_b_24_port, B(23) => 
                           xor_b_23_port, B(22) => xor_b_22_port, B(21) => 
                           xor_b_21_port, B(20) => xor_b_20_port, B(19) => 
                           xor_b_19_port, B(18) => xor_b_18_port, B(17) => 
                           xor_b_17_port, B(16) => xor_b_16_port, B(15) => 
                           xor_b_15_port, B(14) => xor_b_14_port, B(13) => 
                           xor_b_13_port, B(12) => xor_b_12_port, B(11) => 
                           xor_b_11_port, B(10) => xor_b_10_port, B(9) => 
                           xor_b_9_port, B(8) => xor_b_8_port, B(7) => 
                           xor_b_7_port, B(6) => xor_b_6_port, B(5) => 
                           xor_b_5_port, B(4) => xor_b_4_port, B(3) => 
                           xor_b_3_port, B(2) => xor_b_2_port, B(1) => 
                           xor_b_1_port, B(0) => xor_b_0_port, Cin => n3, Co(7)
                           => Cout, Co(6) => carry_6_port, Co(5) => 
                           carry_5_port, Co(4) => carry_4_port, Co(3) => 
                           carry_3_port, Co(2) => carry_2_port, Co(1) => 
                           carry_1_port, Co(0) => carry_0_port);
   SG : sum_generator_n_bit32_n_CSB8_1 port map( A(31) => A(31), A(30) => A(30)
                           , A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(31) => xor_b_31_port, B(30) =>
                           xor_b_30_port, B(29) => xor_b_29_port, B(28) => 
                           xor_b_28_port, B(27) => xor_b_27_port, B(26) => 
                           xor_b_26_port, B(25) => xor_b_25_port, B(24) => 
                           xor_b_24_port, B(23) => xor_b_23_port, B(22) => 
                           xor_b_22_port, B(21) => xor_b_21_port, B(20) => 
                           xor_b_20_port, B(19) => xor_b_19_port, B(18) => 
                           xor_b_18_port, B(17) => xor_b_17_port, B(16) => 
                           xor_b_16_port, B(15) => xor_b_15_port, B(14) => 
                           xor_b_14_port, B(13) => xor_b_13_port, B(12) => 
                           xor_b_12_port, B(11) => xor_b_11_port, B(10) => 
                           xor_b_10_port, B(9) => xor_b_9_port, B(8) => 
                           xor_b_8_port, B(7) => xor_b_7_port, B(6) => 
                           xor_b_6_port, B(5) => xor_b_5_port, B(4) => 
                           xor_b_4_port, B(3) => xor_b_3_port, B(2) => 
                           xor_b_2_port, B(1) => xor_b_1_port, B(0) => 
                           xor_b_0_port, C_in(7) => carry_6_port, C_in(6) => 
                           carry_5_port, C_in(5) => carry_4_port, C_in(4) => 
                           carry_3_port, C_in(3) => carry_2_port, C_in(2) => 
                           carry_1_port, C_in(1) => carry_0_port, C_in(0) => n3
                           , S(31) => S_31_port, S(30) => S_30_port, S(29) => 
                           S_29_port, S(28) => S_28_port, S(27) => S_27_port, 
                           S(26) => S_26_port, S(25) => S_25_port, S(24) => 
                           S_24_port, S(23) => S_23_port, S(22) => S_22_port, 
                           S(21) => S_21_port, S(20) => S_20_port, S(19) => 
                           S_19_port, S(18) => S_18_port, S(17) => S_17_port, 
                           S(16) => S_16_port, S(15) => S_15_port, S(14) => 
                           S_14_port, S(13) => S_13_port, S(12) => S_12_port, 
                           S(11) => S_11_port, S(10) => S_10_port, S(9) => 
                           S_9_port, S(8) => S_8_port, S(7) => S_7_port, S(6) 
                           => S_6_port, S(5) => S_5_port, S(4) => S_4_port, 
                           S(3) => S_3_port, S(2) => S_2_port, S(1) => S_1_port
                           , S(0) => S_0_port);
   U1 : NOR2_X1 port map( A1 => n6, A2 => n5, ZN => ovf);
   U2 : XNOR2_X1 port map( A => A(31), B => S_31_port, ZN => n6);
   U4 : BUF_X2 port map( A => Cin, Z => n3);
   U5 : BUF_X1 port map( A => Cin, Z => n4);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_593 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_593;

architecture SYN_BEHAVIORAL_1 of MUX21_593 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_592 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_592;

architecture SYN_BEHAVIORAL_1 of MUX21_592 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_591 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_591;

architecture SYN_BEHAVIORAL_1 of MUX21_591 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_590 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_590;

architecture SYN_BEHAVIORAL_1 of MUX21_590 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_589 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_589;

architecture SYN_BEHAVIORAL_1 of MUX21_589 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_588 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_588;

architecture SYN_BEHAVIORAL_1 of MUX21_588 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_587 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_587;

architecture SYN_BEHAVIORAL_1 of MUX21_587 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_586 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_586;

architecture SYN_BEHAVIORAL_1 of MUX21_586 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_585 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_585;

architecture SYN_BEHAVIORAL_1 of MUX21_585 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_584 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_584;

architecture SYN_BEHAVIORAL_1 of MUX21_584 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_583 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_583;

architecture SYN_BEHAVIORAL_1 of MUX21_583 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_582 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_582;

architecture SYN_BEHAVIORAL_1 of MUX21_582 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_581 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_581;

architecture SYN_BEHAVIORAL_1 of MUX21_581 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_580 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_580;

architecture SYN_BEHAVIORAL_1 of MUX21_580 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_579 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_579;

architecture SYN_BEHAVIORAL_1 of MUX21_579 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_578 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_578;

architecture SYN_BEHAVIORAL_1 of MUX21_578 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_577 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_577;

architecture SYN_BEHAVIORAL_1 of MUX21_577 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_576 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_576;

architecture SYN_BEHAVIORAL_1 of MUX21_576 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_575 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_575;

architecture SYN_BEHAVIORAL_1 of MUX21_575 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_574 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_574;

architecture SYN_BEHAVIORAL_1 of MUX21_574 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_573 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_573;

architecture SYN_BEHAVIORAL_1 of MUX21_573 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_572 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_572;

architecture SYN_BEHAVIORAL_1 of MUX21_572 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_571 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_571;

architecture SYN_BEHAVIORAL_1 of MUX21_571 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_570 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_570;

architecture SYN_BEHAVIORAL_1 of MUX21_570 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_569 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_569;

architecture SYN_BEHAVIORAL_1 of MUX21_569 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_568 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_568;

architecture SYN_BEHAVIORAL_1 of MUX21_568 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_567 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_567;

architecture SYN_BEHAVIORAL_1 of MUX21_567 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_566 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_566;

architecture SYN_BEHAVIORAL_1 of MUX21_566 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_565 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_565;

architecture SYN_BEHAVIORAL_1 of MUX21_565 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_564 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_564;

architecture SYN_BEHAVIORAL_1 of MUX21_564 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_563 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_563;

architecture SYN_BEHAVIORAL_1 of MUX21_563 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_562 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_562;

architecture SYN_BEHAVIORAL_1 of MUX21_562 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_561 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_561;

architecture SYN_BEHAVIORAL_1 of MUX21_561 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_560 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_560;

architecture SYN_BEHAVIORAL_1 of MUX21_560 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_559 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_559;

architecture SYN_BEHAVIORAL_1 of MUX21_559 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_558 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_558;

architecture SYN_BEHAVIORAL_1 of MUX21_558 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_557 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_557;

architecture SYN_BEHAVIORAL_1 of MUX21_557 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_556 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_556;

architecture SYN_BEHAVIORAL_1 of MUX21_556 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_555 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_555;

architecture SYN_BEHAVIORAL_1 of MUX21_555 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_554 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_554;

architecture SYN_BEHAVIORAL_1 of MUX21_554 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_553 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_553;

architecture SYN_BEHAVIORAL_1 of MUX21_553 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_552 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_552;

architecture SYN_BEHAVIORAL_1 of MUX21_552 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_551 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_551;

architecture SYN_BEHAVIORAL_1 of MUX21_551 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_550 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_550;

architecture SYN_BEHAVIORAL_1 of MUX21_550 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_549 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_549;

architecture SYN_BEHAVIORAL_1 of MUX21_549 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_548 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_548;

architecture SYN_BEHAVIORAL_1 of MUX21_548 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_547 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_547;

architecture SYN_BEHAVIORAL_1 of MUX21_547 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_546 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_546;

architecture SYN_BEHAVIORAL_1 of MUX21_546 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_545 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_545;

architecture SYN_BEHAVIORAL_1 of MUX21_545 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_544 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_544;

architecture SYN_BEHAVIORAL_1 of MUX21_544 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_543 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_543;

architecture SYN_BEHAVIORAL_1 of MUX21_543 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_542 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_542;

architecture SYN_BEHAVIORAL_1 of MUX21_542 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_541 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_541;

architecture SYN_BEHAVIORAL_1 of MUX21_541 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_540 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_540;

architecture SYN_BEHAVIORAL_1 of MUX21_540 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_539 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_539;

architecture SYN_BEHAVIORAL_1 of MUX21_539 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_538 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_538;

architecture SYN_BEHAVIORAL_1 of MUX21_538 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_537 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_537;

architecture SYN_BEHAVIORAL_1 of MUX21_537 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_536 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_536;

architecture SYN_BEHAVIORAL_1 of MUX21_536 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_535 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_535;

architecture SYN_BEHAVIORAL_1 of MUX21_535 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_534 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_534;

architecture SYN_BEHAVIORAL_1 of MUX21_534 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_533 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_533;

architecture SYN_BEHAVIORAL_1 of MUX21_533 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_532 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_532;

architecture SYN_BEHAVIORAL_1 of MUX21_532 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_531 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_531;

architecture SYN_BEHAVIORAL_1 of MUX21_531 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_530 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_530;

architecture SYN_BEHAVIORAL_1 of MUX21_530 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_529 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_529;

architecture SYN_BEHAVIORAL_1 of MUX21_529 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_528 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_528;

architecture SYN_BEHAVIORAL_1 of MUX21_528 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_527 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_527;

architecture SYN_BEHAVIORAL_1 of MUX21_527 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_526 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_526;

architecture SYN_BEHAVIORAL_1 of MUX21_526 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_525 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_525;

architecture SYN_BEHAVIORAL_1 of MUX21_525 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_524 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_524;

architecture SYN_BEHAVIORAL_1 of MUX21_524 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_523 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_523;

architecture SYN_BEHAVIORAL_1 of MUX21_523 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_522 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_522;

architecture SYN_BEHAVIORAL_1 of MUX21_522 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_521 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_521;

architecture SYN_BEHAVIORAL_1 of MUX21_521 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_520 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_520;

architecture SYN_BEHAVIORAL_1 of MUX21_520 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_519 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_519;

architecture SYN_BEHAVIORAL_1 of MUX21_519 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_518 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_518;

architecture SYN_BEHAVIORAL_1 of MUX21_518 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_517 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_517;

architecture SYN_BEHAVIORAL_1 of MUX21_517 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_516 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_516;

architecture SYN_BEHAVIORAL_1 of MUX21_516 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_515 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_515;

architecture SYN_BEHAVIORAL_1 of MUX21_515 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_514 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_514;

architecture SYN_BEHAVIORAL_1 of MUX21_514 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_513 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_513;

architecture SYN_BEHAVIORAL_1 of MUX21_513 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_512 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_512;

architecture SYN_BEHAVIORAL_1 of MUX21_512 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_511 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_511;

architecture SYN_BEHAVIORAL_1 of MUX21_511 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_510 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_510;

architecture SYN_BEHAVIORAL_1 of MUX21_510 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_509 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_509;

architecture SYN_BEHAVIORAL_1 of MUX21_509 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_508 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_508;

architecture SYN_BEHAVIORAL_1 of MUX21_508 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_507 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_507;

architecture SYN_BEHAVIORAL_1 of MUX21_507 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_506 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_506;

architecture SYN_BEHAVIORAL_1 of MUX21_506 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_505 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_505;

architecture SYN_BEHAVIORAL_1 of MUX21_505 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_504 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_504;

architecture SYN_BEHAVIORAL_1 of MUX21_504 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_503 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_503;

architecture SYN_BEHAVIORAL_1 of MUX21_503 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_502 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_502;

architecture SYN_BEHAVIORAL_1 of MUX21_502 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_501 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_501;

architecture SYN_BEHAVIORAL_1 of MUX21_501 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_500 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_500;

architecture SYN_BEHAVIORAL_1 of MUX21_500 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_499 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_499;

architecture SYN_BEHAVIORAL_1 of MUX21_499 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_498 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_498;

architecture SYN_BEHAVIORAL_1 of MUX21_498 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_497 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_497;

architecture SYN_BEHAVIORAL_1 of MUX21_497 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_496 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_496;

architecture SYN_BEHAVIORAL_1 of MUX21_496 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_495 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_495;

architecture SYN_BEHAVIORAL_1 of MUX21_495 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_494 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_494;

architecture SYN_BEHAVIORAL_1 of MUX21_494 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_493 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_493;

architecture SYN_BEHAVIORAL_1 of MUX21_493 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_492 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_492;

architecture SYN_BEHAVIORAL_1 of MUX21_492 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_491 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_491;

architecture SYN_BEHAVIORAL_1 of MUX21_491 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_490 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_490;

architecture SYN_BEHAVIORAL_1 of MUX21_490 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_489 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_489;

architecture SYN_BEHAVIORAL_1 of MUX21_489 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_488 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_488;

architecture SYN_BEHAVIORAL_1 of MUX21_488 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_487 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_487;

architecture SYN_BEHAVIORAL_1 of MUX21_487 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_486 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_486;

architecture SYN_BEHAVIORAL_1 of MUX21_486 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_485 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_485;

architecture SYN_BEHAVIORAL_1 of MUX21_485 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_484 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_484;

architecture SYN_BEHAVIORAL_1 of MUX21_484 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_483 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_483;

architecture SYN_BEHAVIORAL_1 of MUX21_483 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_482 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_482;

architecture SYN_BEHAVIORAL_1 of MUX21_482 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_481 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_481;

architecture SYN_BEHAVIORAL_1 of MUX21_481 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_480 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_480;

architecture SYN_BEHAVIORAL_1 of MUX21_480 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_479 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_479;

architecture SYN_BEHAVIORAL_1 of MUX21_479 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_478 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_478;

architecture SYN_BEHAVIORAL_1 of MUX21_478 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_477 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_477;

architecture SYN_BEHAVIORAL_1 of MUX21_477 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_476 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_476;

architecture SYN_BEHAVIORAL_1 of MUX21_476 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_475 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_475;

architecture SYN_BEHAVIORAL_1 of MUX21_475 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_474 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_474;

architecture SYN_BEHAVIORAL_1 of MUX21_474 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_473 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_473;

architecture SYN_BEHAVIORAL_1 of MUX21_473 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_472 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_472;

architecture SYN_BEHAVIORAL_1 of MUX21_472 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_471 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_471;

architecture SYN_BEHAVIORAL_1 of MUX21_471 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_470 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_470;

architecture SYN_BEHAVIORAL_1 of MUX21_470 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_469 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_469;

architecture SYN_BEHAVIORAL_1 of MUX21_469 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_468 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_468;

architecture SYN_BEHAVIORAL_1 of MUX21_468 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_467 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_467;

architecture SYN_BEHAVIORAL_1 of MUX21_467 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_466 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_466;

architecture SYN_BEHAVIORAL_1 of MUX21_466 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_465 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_465;

architecture SYN_BEHAVIORAL_1 of MUX21_465 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_464 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_464;

architecture SYN_BEHAVIORAL_1 of MUX21_464 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_463 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_463;

architecture SYN_BEHAVIORAL_1 of MUX21_463 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_462 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_462;

architecture SYN_BEHAVIORAL_1 of MUX21_462 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_461 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_461;

architecture SYN_BEHAVIORAL_1 of MUX21_461 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_460 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_460;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_460 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_459 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_459;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_459 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_458 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_458;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_458 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_457 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_457;

architecture SYN_BEHAVIORAL_1_architecture4 of MUX21_457 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_456 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_456;

architecture SYN_BEHAVIORAL_1 of MUX21_456 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_455 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_455;

architecture SYN_BEHAVIORAL_1 of MUX21_455 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_454 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_454;

architecture SYN_BEHAVIORAL_1 of MUX21_454 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_453 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_453;

architecture SYN_BEHAVIORAL_1 of MUX21_453 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_452 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_452;

architecture SYN_BEHAVIORAL_1 of MUX21_452 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_451 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_451;

architecture SYN_BEHAVIORAL_1 of MUX21_451 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_450 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_450;

architecture SYN_BEHAVIORAL_1 of MUX21_450 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_449 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_449;

architecture SYN_BEHAVIORAL_1 of MUX21_449 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_448 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_448;

architecture SYN_BEHAVIORAL_1 of MUX21_448 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_447 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_447;

architecture SYN_BEHAVIORAL_1 of MUX21_447 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_446 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_446;

architecture SYN_BEHAVIORAL_1 of MUX21_446 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_445 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_445;

architecture SYN_BEHAVIORAL_1 of MUX21_445 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_444 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_444;

architecture SYN_BEHAVIORAL_1 of MUX21_444 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_443 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_443;

architecture SYN_BEHAVIORAL_1 of MUX21_443 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_442 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_442;

architecture SYN_BEHAVIORAL_1 of MUX21_442 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_441 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_441;

architecture SYN_BEHAVIORAL_1 of MUX21_441 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_440 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_440;

architecture SYN_BEHAVIORAL_1 of MUX21_440 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_439 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_439;

architecture SYN_BEHAVIORAL_1 of MUX21_439 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_438 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_438;

architecture SYN_BEHAVIORAL_1 of MUX21_438 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_437 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_437;

architecture SYN_BEHAVIORAL_1 of MUX21_437 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_436 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_436;

architecture SYN_BEHAVIORAL_1 of MUX21_436 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_435 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_435;

architecture SYN_BEHAVIORAL_1 of MUX21_435 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_434 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_434;

architecture SYN_BEHAVIORAL_1 of MUX21_434 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_433 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_433;

architecture SYN_BEHAVIORAL_1 of MUX21_433 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_432 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_432;

architecture SYN_BEHAVIORAL_1 of MUX21_432 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_431 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_431;

architecture SYN_BEHAVIORAL_1 of MUX21_431 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_430 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_430;

architecture SYN_BEHAVIORAL_1 of MUX21_430 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_429 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_429;

architecture SYN_BEHAVIORAL_1 of MUX21_429 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_428 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_428;

architecture SYN_BEHAVIORAL_1 of MUX21_428 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_427 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_427;

architecture SYN_BEHAVIORAL_1 of MUX21_427 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_426 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_426;

architecture SYN_BEHAVIORAL_1 of MUX21_426 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_425 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_425;

architecture SYN_BEHAVIORAL_1 of MUX21_425 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_424 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_424;

architecture SYN_BEHAVIORAL_1 of MUX21_424 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_423 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_423;

architecture SYN_BEHAVIORAL_1 of MUX21_423 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_422 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_422;

architecture SYN_BEHAVIORAL_1 of MUX21_422 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_421 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_421;

architecture SYN_BEHAVIORAL_1 of MUX21_421 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_420 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_420;

architecture SYN_BEHAVIORAL_1 of MUX21_420 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_419 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_419;

architecture SYN_BEHAVIORAL_1 of MUX21_419 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_418 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_418;

architecture SYN_BEHAVIORAL_1 of MUX21_418 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_417 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_417;

architecture SYN_BEHAVIORAL_1 of MUX21_417 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_416 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_416;

architecture SYN_BEHAVIORAL_1 of MUX21_416 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_415 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_415;

architecture SYN_BEHAVIORAL_1 of MUX21_415 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_414 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_414;

architecture SYN_BEHAVIORAL_1 of MUX21_414 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_413 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_413;

architecture SYN_BEHAVIORAL_1 of MUX21_413 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_412 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_412;

architecture SYN_BEHAVIORAL_1 of MUX21_412 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_411 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_411;

architecture SYN_BEHAVIORAL_1 of MUX21_411 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_410 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_410;

architecture SYN_BEHAVIORAL_1 of MUX21_410 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_409 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_409;

architecture SYN_BEHAVIORAL_1 of MUX21_409 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_408 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_408;

architecture SYN_BEHAVIORAL_1 of MUX21_408 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_407 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_407;

architecture SYN_BEHAVIORAL_1 of MUX21_407 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_406 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_406;

architecture SYN_BEHAVIORAL_1 of MUX21_406 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_405 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_405;

architecture SYN_BEHAVIORAL_1 of MUX21_405 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_404 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_404;

architecture SYN_BEHAVIORAL_1 of MUX21_404 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_403 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_403;

architecture SYN_BEHAVIORAL_1 of MUX21_403 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_402 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_402;

architecture SYN_BEHAVIORAL_1 of MUX21_402 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_401 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_401;

architecture SYN_BEHAVIORAL_1 of MUX21_401 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_400 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_400;

architecture SYN_BEHAVIORAL_1 of MUX21_400 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_399 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_399;

architecture SYN_BEHAVIORAL_1 of MUX21_399 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_398 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_398;

architecture SYN_BEHAVIORAL_1 of MUX21_398 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_397 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_397;

architecture SYN_BEHAVIORAL_1 of MUX21_397 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_396 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_396;

architecture SYN_BEHAVIORAL_1 of MUX21_396 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_395 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_395;

architecture SYN_BEHAVIORAL_1 of MUX21_395 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_394 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_394;

architecture SYN_BEHAVIORAL_1 of MUX21_394 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_393 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_393;

architecture SYN_BEHAVIORAL_1 of MUX21_393 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_392 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_392;

architecture SYN_BEHAVIORAL_1 of MUX21_392 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_391 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_391;

architecture SYN_BEHAVIORAL_1 of MUX21_391 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_390 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_390;

architecture SYN_BEHAVIORAL_1 of MUX21_390 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_389 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_389;

architecture SYN_BEHAVIORAL_1 of MUX21_389 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_388 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_388;

architecture SYN_BEHAVIORAL_1 of MUX21_388 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_387 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_387;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_387 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U2 : INV_X1 port map( A => S, ZN => n2);
   U3 : INV_X1 port map( A => n4, ZN => Y);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_386 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_386;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_386 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U2 : INV_X1 port map( A => S, ZN => n2);
   U3 : INV_X1 port map( A => n4, ZN => Y);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_385 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_385;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_385 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_384 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_384;

architecture SYN_BEHAVIORAL_1 of MUX21_384 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_383 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_383;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_383 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_382 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_382;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_382 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_381 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_381;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_381 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_380 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_380;

architecture SYN_BEHAVIORAL_1 of MUX21_380 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_379 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_379;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_379 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_378 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_378;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_378 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_377 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_377;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_377 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U2 : INV_X1 port map( A => S, ZN => n2);
   U3 : INV_X1 port map( A => n4, ZN => Y);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_376 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_376;

architecture SYN_BEHAVIORAL_1 of MUX21_376 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_375 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_375;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_375 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U2 : INV_X1 port map( A => S, ZN => n2);
   U3 : INV_X1 port map( A => n4, ZN => Y);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_374 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_374;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_374 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U2 : INV_X1 port map( A => S, ZN => n2);
   U3 : INV_X1 port map( A => n4, ZN => Y);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_373 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_373;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_373 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U2 : INV_X1 port map( A => S, ZN => n2);
   U3 : INV_X1 port map( A => n4, ZN => Y);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_372 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_372;

architecture SYN_BEHAVIORAL_1 of MUX21_372 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_371 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_371;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_371 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U2 : INV_X1 port map( A => S, ZN => n2);
   U3 : INV_X1 port map( A => n4, ZN => Y);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_370 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_370;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_370 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U2 : INV_X1 port map( A => S, ZN => n2);
   U3 : INV_X1 port map( A => n4, ZN => Y);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_369 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_369;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_369 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U2 : INV_X1 port map( A => S, ZN => n2);
   U3 : INV_X1 port map( A => n4, ZN => Y);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_368 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_368;

architecture SYN_BEHAVIORAL_1 of MUX21_368 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_367 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_367;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_367 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U2 : INV_X1 port map( A => S, ZN => n2);
   U3 : INV_X1 port map( A => n4, ZN => Y);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_366 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_366;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_366 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U2 : INV_X1 port map( A => S, ZN => n2);
   U3 : INV_X1 port map( A => n4, ZN => Y);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_365 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_365;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_365 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U2 : INV_X1 port map( A => S, ZN => n2);
   U3 : INV_X1 port map( A => n4, ZN => Y);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_364 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_364;

architecture SYN_BEHAVIORAL_1 of MUX21_364 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_363 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_363;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_363 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U2 : INV_X1 port map( A => S, ZN => n2);
   U3 : INV_X1 port map( A => n4, ZN => Y);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_362 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_362;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_362 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U2 : INV_X1 port map( A => S, ZN => n2);
   U3 : INV_X1 port map( A => n4, ZN => Y);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_361 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_361;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_361 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_360 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_360;

architecture SYN_BEHAVIORAL_1 of MUX21_360 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_359 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_359;

architecture SYN_BEHAVIORAL_1 of MUX21_359 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_358 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_358;

architecture SYN_BEHAVIORAL_1 of MUX21_358 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_357 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_357;

architecture SYN_BEHAVIORAL_1 of MUX21_357 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_356 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_356;

architecture SYN_BEHAVIORAL_1 of MUX21_356 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_355 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_355;

architecture SYN_BEHAVIORAL_1 of MUX21_355 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_354 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_354;

architecture SYN_BEHAVIORAL_1 of MUX21_354 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_353 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_353;

architecture SYN_BEHAVIORAL_1 of MUX21_353 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_352 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_352;

architecture SYN_BEHAVIORAL_1 of MUX21_352 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_351 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_351;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_351 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_350 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_350;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_350 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_349 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_349;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_349 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_348 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_348;

architecture SYN_BEHAVIORAL_1_architecture4 of MUX21_348 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_347 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_347;

architecture SYN_BEHAVIORAL_1_architecture5 of MUX21_347 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture5;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_346 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_346;

architecture SYN_BEHAVIORAL_1_architecture6 of MUX21_346 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture6;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_345 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_345;

architecture SYN_BEHAVIORAL_1_architecture7 of MUX21_345 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture7;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_344 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_344;

architecture SYN_BEHAVIORAL_1 of MUX21_344 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_343 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_343;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_343 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_342 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_342;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_342 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_341 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_341;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_341 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_340 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_340;

architecture SYN_BEHAVIORAL_1_architecture4 of MUX21_340 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_339 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_339;

architecture SYN_BEHAVIORAL_1_architecture5 of MUX21_339 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture5;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_338 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_338;

architecture SYN_BEHAVIORAL_1_architecture6 of MUX21_338 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture6;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_337 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_337;

architecture SYN_BEHAVIORAL_1_architecture7 of MUX21_337 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture7;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_336 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_336;

architecture SYN_BEHAVIORAL_1 of MUX21_336 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_335 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_335;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_335 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_334 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_334;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_334 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_333 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_333;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_333 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_332 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_332;

architecture SYN_BEHAVIORAL_1_architecture4 of MUX21_332 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_331 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_331;

architecture SYN_BEHAVIORAL_1_architecture5 of MUX21_331 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture5;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_330 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_330;

architecture SYN_BEHAVIORAL_1_architecture6 of MUX21_330 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture6;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_329 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_329;

architecture SYN_BEHAVIORAL_1_architecture7 of MUX21_329 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture7;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_328 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_328;

architecture SYN_BEHAVIORAL_1 of MUX21_328 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_327 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_327;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_327 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_326 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_326;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_326 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_325 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_325;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_325 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_324 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_324;

architecture SYN_BEHAVIORAL_1_architecture4 of MUX21_324 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_323 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_323;

architecture SYN_BEHAVIORAL_1_architecture5 of MUX21_323 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture5;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_322 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_322;

architecture SYN_BEHAVIORAL_1_architecture6 of MUX21_322 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture6;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_321 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_321;

architecture SYN_BEHAVIORAL_1_architecture7 of MUX21_321 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture7;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_320 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_320;

architecture SYN_BEHAVIORAL_1 of MUX21_320 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_319 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_319;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_319 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_318 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_318;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_318 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_317 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_317;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_317 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_316 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_316;

architecture SYN_BEHAVIORAL_1_architecture4 of MUX21_316 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_315 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_315;

architecture SYN_BEHAVIORAL_1_architecture5 of MUX21_315 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture5;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_314 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_314;

architecture SYN_BEHAVIORAL_1_architecture6 of MUX21_314 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture6;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_313 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_313;

architecture SYN_BEHAVIORAL_1_architecture7 of MUX21_313 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture7;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_312 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_312;

architecture SYN_BEHAVIORAL_1 of MUX21_312 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_311 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_311;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_311 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_310 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_310;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_310 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_309 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_309;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_309 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_308 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_308;

architecture SYN_BEHAVIORAL_1_architecture4 of MUX21_308 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_307 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_307;

architecture SYN_BEHAVIORAL_1_architecture5 of MUX21_307 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture5;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_306 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_306;

architecture SYN_BEHAVIORAL_1_architecture6 of MUX21_306 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture6;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_305 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_305;

architecture SYN_BEHAVIORAL_1_architecture7 of MUX21_305 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture7;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_304 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_304;

architecture SYN_BEHAVIORAL_1 of MUX21_304 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_303 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_303;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_303 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_302 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_302;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_302 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_301 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_301;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_301 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_300 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_300;

architecture SYN_BEHAVIORAL_1_architecture4 of MUX21_300 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_299 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_299;

architecture SYN_BEHAVIORAL_1_architecture5 of MUX21_299 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture5;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_298 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_298;

architecture SYN_BEHAVIORAL_1_architecture6 of MUX21_298 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture6;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_297 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_297;

architecture SYN_BEHAVIORAL_1_architecture7 of MUX21_297 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture7;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_296 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_296;

architecture SYN_BEHAVIORAL_1 of MUX21_296 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_295 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_295;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_295 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_294 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_294;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_294 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_293 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_293;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_293 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_292 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_292;

architecture SYN_BEHAVIORAL_1_architecture4 of MUX21_292 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_291 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_291;

architecture SYN_BEHAVIORAL_1_architecture5 of MUX21_291 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture5;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_290 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_290;

architecture SYN_BEHAVIORAL_1_architecture6 of MUX21_290 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture6;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_289 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_289;

architecture SYN_BEHAVIORAL_1_architecture7 of MUX21_289 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture7;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_288 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_288;

architecture SYN_BEHAVIORAL_1 of MUX21_288 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_287 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_287;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_287 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_286 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_286;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_286 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_285 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_285;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_285 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_284 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_284;

architecture SYN_BEHAVIORAL_1_architecture4 of MUX21_284 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_283 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_283;

architecture SYN_BEHAVIORAL_1_architecture5 of MUX21_283 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture5;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_282 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_282;

architecture SYN_BEHAVIORAL_1_architecture6 of MUX21_282 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture6;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_281 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_281;

architecture SYN_BEHAVIORAL_1_architecture7 of MUX21_281 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture7;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_280 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_280;

architecture SYN_BEHAVIORAL_1 of MUX21_280 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_279 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_279;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_279 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_278 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_278;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_278 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_277 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_277;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_277 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_276 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_276;

architecture SYN_BEHAVIORAL_1_architecture4 of MUX21_276 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_275 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_275;

architecture SYN_BEHAVIORAL_1_architecture5 of MUX21_275 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture5;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_274 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_274;

architecture SYN_BEHAVIORAL_1_architecture6 of MUX21_274 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture6;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_273 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_273;

architecture SYN_BEHAVIORAL_1_architecture7 of MUX21_273 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture7;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_272 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_272;

architecture SYN_BEHAVIORAL_1 of MUX21_272 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_271 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_271;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_271 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_270 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_270;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_270 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_269 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_269;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_269 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_268 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_268;

architecture SYN_BEHAVIORAL_1_architecture4 of MUX21_268 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_267 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_267;

architecture SYN_BEHAVIORAL_1_architecture5 of MUX21_267 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture5;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_266 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_266;

architecture SYN_BEHAVIORAL_1_architecture6 of MUX21_266 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture6;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_265 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_265;

architecture SYN_BEHAVIORAL_1_architecture7 of MUX21_265 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture7;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_264 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_264;

architecture SYN_BEHAVIORAL_1 of MUX21_264 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_263 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_263;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_263 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_262 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_262;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_262 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_261 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_261;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_261 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_260 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_260;

architecture SYN_BEHAVIORAL_1_architecture4 of MUX21_260 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_259 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_259;

architecture SYN_BEHAVIORAL_1_architecture5 of MUX21_259 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture5;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_258 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_258;

architecture SYN_BEHAVIORAL_1_architecture6 of MUX21_258 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture6;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_257 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_257;

architecture SYN_BEHAVIORAL_1_architecture7 of MUX21_257 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture7;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_256 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_256;

architecture SYN_BEHAVIORAL_1 of MUX21_256 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_255 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_255;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_255 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_254 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_254;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_254 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_253 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_253;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_253 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_252 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_252;

architecture SYN_BEHAVIORAL_1_architecture4 of MUX21_252 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_251 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_251;

architecture SYN_BEHAVIORAL_1_architecture5 of MUX21_251 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture5;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_250 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_250;

architecture SYN_BEHAVIORAL_1_architecture6 of MUX21_250 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture6;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_249 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_249;

architecture SYN_BEHAVIORAL_1_architecture7 of MUX21_249 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture7;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_248 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_248;

architecture SYN_BEHAVIORAL_1 of MUX21_248 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_247 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_247;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_247 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_246 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_246;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_246 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_245 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_245;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_245 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_244 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_244;

architecture SYN_BEHAVIORAL_1_architecture4 of MUX21_244 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_243 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_243;

architecture SYN_BEHAVIORAL_1_architecture5 of MUX21_243 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture5;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_242 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_242;

architecture SYN_BEHAVIORAL_1_architecture6 of MUX21_242 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture6;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_241 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_241;

architecture SYN_BEHAVIORAL_1_architecture7 of MUX21_241 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture7;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_240 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_240;

architecture SYN_BEHAVIORAL_1 of MUX21_240 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_239 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_239;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_239 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_238 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_238;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_238 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_237 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_237;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_237 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_236 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_236;

architecture SYN_BEHAVIORAL_1_architecture4 of MUX21_236 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_235 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_235;

architecture SYN_BEHAVIORAL_1_architecture5 of MUX21_235 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture5;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_234 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_234;

architecture SYN_BEHAVIORAL_1_architecture6 of MUX21_234 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture6;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_233 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_233;

architecture SYN_BEHAVIORAL_1_architecture7 of MUX21_233 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture7;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_232 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_232;

architecture SYN_BEHAVIORAL_1 of MUX21_232 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_231 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_231;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_231 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_230 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_230;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_230 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_229 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_229;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_229 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_228 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_228;

architecture SYN_BEHAVIORAL_1_architecture4 of MUX21_228 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_227 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_227;

architecture SYN_BEHAVIORAL_1_architecture5 of MUX21_227 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture5;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_226 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_226;

architecture SYN_BEHAVIORAL_1_architecture6 of MUX21_226 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture6;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_225 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_225;

architecture SYN_BEHAVIORAL_1_architecture7 of MUX21_225 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture7;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_224 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_224;

architecture SYN_BEHAVIORAL_1 of MUX21_224 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_223 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_223;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_223 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_222 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_222;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_222 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_221 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_221;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_221 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_220 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_220;

architecture SYN_BEHAVIORAL_1 of MUX21_220 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_219 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_219;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_219 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_218 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_218;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_218 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_217 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_217;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_217 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_216 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_216;

architecture SYN_BEHAVIORAL_1 of MUX21_216 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_215 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_215;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_215 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_214 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_214;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_214 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_213 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_213;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_213 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_212 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_212;

architecture SYN_BEHAVIORAL_1 of MUX21_212 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_211 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_211;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_211 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_210 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_210;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_210 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_209 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_209;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_209 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_208 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_208;

architecture SYN_BEHAVIORAL_1 of MUX21_208 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_207 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_207;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_207 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_206 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_206;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_206 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_205 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_205;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_205 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_204 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_204;

architecture SYN_BEHAVIORAL_1 of MUX21_204 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_203 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_203;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_203 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_202 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_202;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_202 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_201 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_201;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_201 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_200 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_200;

architecture SYN_BEHAVIORAL_1 of MUX21_200 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_199 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_199;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_199 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_198 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_198;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_198 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_197 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_197;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_197 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_196 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_196;

architecture SYN_BEHAVIORAL_1 of MUX21_196 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_195 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_195;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_195 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_194 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_194;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_194 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_193 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_193;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_193 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_192 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_192;

architecture SYN_BEHAVIORAL_1 of MUX21_192 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_191 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_191;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_191 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_190 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_190;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_190 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_189 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_189;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_189 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_188 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_188;

architecture SYN_BEHAVIORAL_1 of MUX21_188 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_187 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_187;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_187 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_186 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_186;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_186 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_185 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_185;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_185 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_184 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_184;

architecture SYN_BEHAVIORAL_1 of MUX21_184 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_183 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_183;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_183 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_182 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_182;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_182 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_181 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_181;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_181 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_180 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_180;

architecture SYN_BEHAVIORAL_1 of MUX21_180 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_179 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_179;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_179 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_178 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_178;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_178 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_177 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_177;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_177 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_176 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_176;

architecture SYN_BEHAVIORAL_1 of MUX21_176 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_175 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_175;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_175 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_174 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_174;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_174 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_173 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_173;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_173 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_172 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_172;

architecture SYN_BEHAVIORAL_1 of MUX21_172 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_171 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_171;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_171 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_170 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_170;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_170 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_169 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_169;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_169 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_168 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_168;

architecture SYN_BEHAVIORAL_1 of MUX21_168 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_167 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_167;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_167 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_166 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_166;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_166 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_165 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_165;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_165 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_164 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_164;

architecture SYN_BEHAVIORAL_1 of MUX21_164 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_163 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_163;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_163 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_162 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_162;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_162 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_161 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_161;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_161 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_160 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_160;

architecture SYN_BEHAVIORAL_1 of MUX21_160 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_159 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_159;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_159 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_158 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_158;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_158 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_157 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_157;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_157 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_156 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_156;

architecture SYN_BEHAVIORAL_1 of MUX21_156 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_155 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_155;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_155 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_154 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_154;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_154 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_153 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_153;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_153 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_152 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_152;

architecture SYN_BEHAVIORAL_1 of MUX21_152 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_151 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_151;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_151 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_150 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_150;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_150 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_149 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_149;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_149 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_148 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_148;

architecture SYN_BEHAVIORAL_1 of MUX21_148 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_147 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_147;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_147 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_146 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_146;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_146 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_145 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_145;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_145 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_144 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_144;

architecture SYN_BEHAVIORAL_1 of MUX21_144 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_143 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_143;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_143 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_142 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_142;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_142 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_141 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_141;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_141 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_140 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_140;

architecture SYN_BEHAVIORAL_1 of MUX21_140 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_139 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_139;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_139 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_138 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_138;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_138 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_137 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_137;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_137 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_136 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_136;

architecture SYN_BEHAVIORAL_1 of MUX21_136 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_135 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_135;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_135 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_134 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_134;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_134 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_133 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_133;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_133 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_132 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_132;

architecture SYN_BEHAVIORAL_1 of MUX21_132 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_131 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_131;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_131 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_130 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_130;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_130 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_129 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_129;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_129 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_128 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_128;

architecture SYN_BEHAVIORAL_1 of MUX21_128 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_127 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_127;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_127 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_126 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_126;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_126 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_125 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_125;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_125 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_124 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_124;

architecture SYN_BEHAVIORAL_1 of MUX21_124 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_123 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_123;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_123 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_122 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_122;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_122 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_121 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_121;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_121 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_120 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_120;

architecture SYN_BEHAVIORAL_1 of MUX21_120 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_119 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_119;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_119 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_118 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_118;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_118 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_117 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_117;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_117 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_116 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_116;

architecture SYN_BEHAVIORAL_1 of MUX21_116 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_115 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_115;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_115 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_114 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_114;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_114 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_113 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_113;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_113 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_112 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_112;

architecture SYN_BEHAVIORAL_1 of MUX21_112 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_111 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_111;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_111 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_110 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_110;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_110 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_109 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_109;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_109 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_108 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_108;

architecture SYN_BEHAVIORAL_1 of MUX21_108 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_107 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_107;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_107 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_106 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_106;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_106 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_105 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_105;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_105 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_104 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_104;

architecture SYN_BEHAVIORAL_1 of MUX21_104 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_103 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_103;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_103 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_102 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_102;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_102 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_101 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_101;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_101 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_100 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_100;

architecture SYN_BEHAVIORAL_1 of MUX21_100 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_99 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_99;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_99 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_98 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_98;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_98 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_97 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_97;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_97 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_96 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_96;

architecture SYN_BEHAVIORAL_1 of MUX21_96 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_95 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_95;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_95 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_94 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_94;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_94 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_93 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_93;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_93 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_92 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_92;

architecture SYN_BEHAVIORAL_1 of MUX21_92 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_91 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_91;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_91 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_90 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_90;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_90 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_89 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_89;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_89 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_88 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_88;

architecture SYN_BEHAVIORAL_1 of MUX21_88 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_87 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_87;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_87 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_86 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_86;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_86 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_85 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_85;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_85 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_84 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_84;

architecture SYN_BEHAVIORAL_1 of MUX21_84 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_83 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_83;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_83 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_82 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_82;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_82 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_81 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_81;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_81 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_80 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_80;

architecture SYN_BEHAVIORAL_1 of MUX21_80 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_79 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_79;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_79 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_78 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_78;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_78 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_77 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_77;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_77 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_76 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_76;

architecture SYN_BEHAVIORAL_1 of MUX21_76 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_75 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_75;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_75 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_74 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_74;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_74 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_73 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_73;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_73 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_72 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_72;

architecture SYN_BEHAVIORAL_1 of MUX21_72 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_71 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_71;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_71 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_70 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_70;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_70 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_69 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_69;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_69 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_68 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_68;

architecture SYN_BEHAVIORAL_1 of MUX21_68 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_67 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_67;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_67 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_66 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_66;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_66 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_65 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_65;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_65 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => S, ZN => n2);
   U2 : INV_X1 port map( A => n4, ZN => Y);
   U3 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_64 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_64;

architecture SYN_BEHAVIORAL_1 of MUX21_64 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_63 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_63;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_63 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_62 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_62;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_62 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_61 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_61;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_61 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_60 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_60;

architecture SYN_BEHAVIORAL_1 of MUX21_60 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_59 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_59;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_59 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_58 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_58;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_58 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_57 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_57;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_57 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_56 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_56;

architecture SYN_BEHAVIORAL_1 of MUX21_56 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_55 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_55;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_55 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_54 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_54;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_54 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_53 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_53;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_53 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_52 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_52;

architecture SYN_BEHAVIORAL_1 of MUX21_52 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_51 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_51;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_51 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_50 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_50;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_50 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_49 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_49;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_49 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_48 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_48;

architecture SYN_BEHAVIORAL_1 of MUX21_48 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_47 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_47;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_47 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_46 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_46;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_46 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_45 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_45;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_45 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_44 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_44;

architecture SYN_BEHAVIORAL_1 of MUX21_44 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_43 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_43;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_43 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_42 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_42;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_42 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_41 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_41;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_41 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_40 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_40;

architecture SYN_BEHAVIORAL_1 of MUX21_40 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_39 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_39;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_39 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_38 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_38;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_38 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_37 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_37;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_37 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_36 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_36;

architecture SYN_BEHAVIORAL_1 of MUX21_36 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_35 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_35;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_35 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_34 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_34;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_34 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_33 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_33;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_33 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_32 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_32;

architecture SYN_BEHAVIORAL_1 of MUX21_32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_31 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_31;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_31 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_30 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_30;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_30 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_29 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_29;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_29 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_28 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_28;

architecture SYN_BEHAVIORAL_1 of MUX21_28 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_27 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_27;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_27 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_26 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_26;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_26 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_25 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_25;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_25 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_24 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_24;

architecture SYN_BEHAVIORAL_1 of MUX21_24 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_23 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_23;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_23 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_22 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_22;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_22 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_21 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_21;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_21 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_20 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_20;

architecture SYN_BEHAVIORAL_1 of MUX21_20 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_19 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_19;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_19 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_18 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_18;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_18 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_17 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_17;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_17 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_16 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_16;

architecture SYN_BEHAVIORAL_1 of MUX21_16 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_15 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_15;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_15 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_14 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_14;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_14 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_13 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_13;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_13 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_12 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_12;

architecture SYN_BEHAVIORAL_1 of MUX21_12 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_11 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_11;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_11 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_10 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_10;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_10 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_9 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_9;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_9 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_8 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_8;

architecture SYN_BEHAVIORAL_1 of MUX21_8 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_7 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_7;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_7 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_6 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_6;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_5 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_5;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_4 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_4;

architecture SYN_BEHAVIORAL_1 of MUX21_4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_3 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_3;

architecture SYN_BEHAVIORAL_1_architecture of MUX21_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_2 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_2;

architecture SYN_BEHAVIORAL_1_architecture2 of MUX21_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_1 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_1;

architecture SYN_BEHAVIORAL_1_architecture3 of MUX21_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n4, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n2, B1 => S, B2 => B, ZN => n4);
   U3 : INV_X1 port map( A => S, ZN => n2);

end SYN_BEHAVIORAL_1_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT32_5 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX21_GENERIC_NBIT32_5;

architecture SYN_structural of MUX21_GENERIC_NBIT32_5 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX21_531
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_532
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_533
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_534
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_535
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_536
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_537
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_538
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_539
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_540
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_541
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_542
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_543
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_544
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_545
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_546
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_547
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_548
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_549
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_550
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_551
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_552
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_553
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_554
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_555
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_556
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_557
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_558
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_559
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_560
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_561
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_562
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   MUXES_0 : MUX21_562 port map( A => A(0), B => B(0), S => n1, Y => Y(0));
   MUXES_1 : MUX21_561 port map( A => A(1), B => B(1), S => n1, Y => Y(1));
   MUXES_2 : MUX21_560 port map( A => A(2), B => B(2), S => n1, Y => Y(2));
   MUXES_3 : MUX21_559 port map( A => A(3), B => B(3), S => n1, Y => Y(3));
   MUXES_4 : MUX21_558 port map( A => A(4), B => B(4), S => n1, Y => Y(4));
   MUXES_5 : MUX21_557 port map( A => A(5), B => B(5), S => n1, Y => Y(5));
   MUXES_6 : MUX21_556 port map( A => A(6), B => B(6), S => n1, Y => Y(6));
   MUXES_7 : MUX21_555 port map( A => A(7), B => B(7), S => n1, Y => Y(7));
   MUXES_8 : MUX21_554 port map( A => A(8), B => B(8), S => n1, Y => Y(8));
   MUXES_9 : MUX21_553 port map( A => A(9), B => B(9), S => n1, Y => Y(9));
   MUXES_10 : MUX21_552 port map( A => A(10), B => B(10), S => n1, Y => Y(10));
   MUXES_11 : MUX21_551 port map( A => A(11), B => B(11), S => n1, Y => Y(11));
   MUXES_12 : MUX21_550 port map( A => A(12), B => B(12), S => n2, Y => Y(12));
   MUXES_13 : MUX21_549 port map( A => A(13), B => B(13), S => n2, Y => Y(13));
   MUXES_14 : MUX21_548 port map( A => A(14), B => B(14), S => n2, Y => Y(14));
   MUXES_15 : MUX21_547 port map( A => A(15), B => B(15), S => n2, Y => Y(15));
   MUXES_16 : MUX21_546 port map( A => A(16), B => B(16), S => n2, Y => Y(16));
   MUXES_17 : MUX21_545 port map( A => A(17), B => B(17), S => n2, Y => Y(17));
   MUXES_18 : MUX21_544 port map( A => A(18), B => B(18), S => n2, Y => Y(18));
   MUXES_19 : MUX21_543 port map( A => A(19), B => B(19), S => n2, Y => Y(19));
   MUXES_20 : MUX21_542 port map( A => A(20), B => B(20), S => n2, Y => Y(20));
   MUXES_21 : MUX21_541 port map( A => A(21), B => B(21), S => n2, Y => Y(21));
   MUXES_22 : MUX21_540 port map( A => A(22), B => B(22), S => n2, Y => Y(22));
   MUXES_23 : MUX21_539 port map( A => A(23), B => B(23), S => n2, Y => Y(23));
   MUXES_24 : MUX21_538 port map( A => A(24), B => B(24), S => n3, Y => Y(24));
   MUXES_25 : MUX21_537 port map( A => A(25), B => B(25), S => n3, Y => Y(25));
   MUXES_26 : MUX21_536 port map( A => A(26), B => B(26), S => n3, Y => Y(26));
   MUXES_27 : MUX21_535 port map( A => A(27), B => B(27), S => n3, Y => Y(27));
   MUXES_28 : MUX21_534 port map( A => A(28), B => B(28), S => n3, Y => Y(28));
   MUXES_29 : MUX21_533 port map( A => A(29), B => B(29), S => n3, Y => Y(29));
   MUXES_30 : MUX21_532 port map( A => A(30), B => B(30), S => n3, Y => Y(30));
   MUXES_31 : MUX21_531 port map( A => A(31), B => B(31), S => n3, Y => Y(31));
   U1 : BUF_X1 port map( A => SEL, Z => n2);
   U2 : BUF_X1 port map( A => SEL, Z => n1);
   U3 : BUF_X1 port map( A => SEL, Z => n3);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT32_4 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX21_GENERIC_NBIT32_4;

architecture SYN_structural of MUX21_GENERIC_NBIT32_4 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX21_499
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_500
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_501
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_502
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_503
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_504
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_505
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_506
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_507
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_508
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_509
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_510
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_511
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_512
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_513
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_514
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_515
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_516
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_517
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_518
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_519
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_520
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_521
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_522
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_523
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_524
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_525
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_526
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_527
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_528
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_529
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_530
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   MUXES_0 : MUX21_530 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_529 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_528 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_527 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));
   MUXES_4 : MUX21_526 port map( A => A(4), B => B(4), S => SEL, Y => Y(4));
   MUXES_5 : MUX21_525 port map( A => A(5), B => B(5), S => n2, Y => Y(5));
   MUXES_6 : MUX21_524 port map( A => A(6), B => B(6), S => n1, Y => Y(6));
   MUXES_7 : MUX21_523 port map( A => A(7), B => B(7), S => n1, Y => Y(7));
   MUXES_8 : MUX21_522 port map( A => A(8), B => B(8), S => n1, Y => Y(8));
   MUXES_9 : MUX21_521 port map( A => A(9), B => B(9), S => n1, Y => Y(9));
   MUXES_10 : MUX21_520 port map( A => A(10), B => B(10), S => n2, Y => Y(10));
   MUXES_11 : MUX21_519 port map( A => A(11), B => B(11), S => n1, Y => Y(11));
   MUXES_12 : MUX21_518 port map( A => A(12), B => B(12), S => n1, Y => Y(12));
   MUXES_13 : MUX21_517 port map( A => A(13), B => B(13), S => n1, Y => Y(13));
   MUXES_14 : MUX21_516 port map( A => A(14), B => B(14), S => n1, Y => Y(14));
   MUXES_15 : MUX21_515 port map( A => A(15), B => B(15), S => n1, Y => Y(15));
   MUXES_16 : MUX21_514 port map( A => A(16), B => B(16), S => n1, Y => Y(16));
   MUXES_17 : MUX21_513 port map( A => A(17), B => B(17), S => n1, Y => Y(17));
   MUXES_18 : MUX21_512 port map( A => A(18), B => B(18), S => n1, Y => Y(18));
   MUXES_19 : MUX21_511 port map( A => A(19), B => B(19), S => n1, Y => Y(19));
   MUXES_20 : MUX21_510 port map( A => A(20), B => B(20), S => n1, Y => Y(20));
   MUXES_21 : MUX21_509 port map( A => A(21), B => B(21), S => n1, Y => Y(21));
   MUXES_22 : MUX21_508 port map( A => A(22), B => B(22), S => n1, Y => Y(22));
   MUXES_23 : MUX21_507 port map( A => A(23), B => B(23), S => n1, Y => Y(23));
   MUXES_24 : MUX21_506 port map( A => A(24), B => B(24), S => n2, Y => Y(24));
   MUXES_25 : MUX21_505 port map( A => A(25), B => B(25), S => n2, Y => Y(25));
   MUXES_26 : MUX21_504 port map( A => A(26), B => B(26), S => n2, Y => Y(26));
   MUXES_27 : MUX21_503 port map( A => A(27), B => B(27), S => n1, Y => Y(27));
   MUXES_28 : MUX21_502 port map( A => A(28), B => B(28), S => n2, Y => Y(28));
   MUXES_29 : MUX21_501 port map( A => A(29), B => B(29), S => n1, Y => Y(29));
   MUXES_30 : MUX21_500 port map( A => A(30), B => B(30), S => SEL, Y => Y(30))
                           ;
   MUXES_31 : MUX21_499 port map( A => A(31), B => B(31), S => SEL, Y => Y(31))
                           ;
   U1 : BUF_X2 port map( A => SEL, Z => n1);
   U2 : CLKBUF_X1 port map( A => SEL, Z => n2);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT32_3 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX21_GENERIC_NBIT32_3;

architecture SYN_structural of MUX21_GENERIC_NBIT32_3 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX21_467
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_468
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_469
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_470
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_471
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_472
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_473
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_474
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_475
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_476
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_477
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_478
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_479
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_480
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_481
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_482
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_483
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_484
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_485
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_486
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_487
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_488
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_489
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_490
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_491
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_492
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_493
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_494
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_495
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_496
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_497
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_498
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   MUXES_0 : MUX21_498 port map( A => A(0), B => B(0), S => n1, Y => Y(0));
   MUXES_1 : MUX21_497 port map( A => A(1), B => B(1), S => n1, Y => Y(1));
   MUXES_2 : MUX21_496 port map( A => A(2), B => B(2), S => n1, Y => Y(2));
   MUXES_3 : MUX21_495 port map( A => A(3), B => B(3), S => n1, Y => Y(3));
   MUXES_4 : MUX21_494 port map( A => A(4), B => B(4), S => n1, Y => Y(4));
   MUXES_5 : MUX21_493 port map( A => A(5), B => B(5), S => n1, Y => Y(5));
   MUXES_6 : MUX21_492 port map( A => A(6), B => B(6), S => n1, Y => Y(6));
   MUXES_7 : MUX21_491 port map( A => A(7), B => B(7), S => n1, Y => Y(7));
   MUXES_8 : MUX21_490 port map( A => A(8), B => B(8), S => n1, Y => Y(8));
   MUXES_9 : MUX21_489 port map( A => A(9), B => B(9), S => n1, Y => Y(9));
   MUXES_10 : MUX21_488 port map( A => A(10), B => B(10), S => n1, Y => Y(10));
   MUXES_11 : MUX21_487 port map( A => A(11), B => B(11), S => n1, Y => Y(11));
   MUXES_12 : MUX21_486 port map( A => A(12), B => B(12), S => n2, Y => Y(12));
   MUXES_13 : MUX21_485 port map( A => A(13), B => B(13), S => n2, Y => Y(13));
   MUXES_14 : MUX21_484 port map( A => A(14), B => B(14), S => n2, Y => Y(14));
   MUXES_15 : MUX21_483 port map( A => A(15), B => B(15), S => n2, Y => Y(15));
   MUXES_16 : MUX21_482 port map( A => A(16), B => B(16), S => n2, Y => Y(16));
   MUXES_17 : MUX21_481 port map( A => A(17), B => B(17), S => n2, Y => Y(17));
   MUXES_18 : MUX21_480 port map( A => A(18), B => B(18), S => n2, Y => Y(18));
   MUXES_19 : MUX21_479 port map( A => A(19), B => B(19), S => n2, Y => Y(19));
   MUXES_20 : MUX21_478 port map( A => A(20), B => B(20), S => n2, Y => Y(20));
   MUXES_21 : MUX21_477 port map( A => A(21), B => B(21), S => n2, Y => Y(21));
   MUXES_22 : MUX21_476 port map( A => A(22), B => B(22), S => n2, Y => Y(22));
   MUXES_23 : MUX21_475 port map( A => A(23), B => B(23), S => n2, Y => Y(23));
   MUXES_24 : MUX21_474 port map( A => A(24), B => B(24), S => n3, Y => Y(24));
   MUXES_25 : MUX21_473 port map( A => A(25), B => B(25), S => n3, Y => Y(25));
   MUXES_26 : MUX21_472 port map( A => A(26), B => B(26), S => n3, Y => Y(26));
   MUXES_27 : MUX21_471 port map( A => A(27), B => B(27), S => n3, Y => Y(27));
   MUXES_28 : MUX21_470 port map( A => A(28), B => B(28), S => n3, Y => Y(28));
   MUXES_29 : MUX21_469 port map( A => A(29), B => B(29), S => n3, Y => Y(29));
   MUXES_30 : MUX21_468 port map( A => A(30), B => B(30), S => n3, Y => Y(30));
   MUXES_31 : MUX21_467 port map( A => A(31), B => B(31), S => n3, Y => Y(31));
   U1 : BUF_X1 port map( A => SEL, Z => n2);
   U2 : BUF_X1 port map( A => SEL, Z => n1);
   U3 : BUF_X1 port map( A => SEL, Z => n3);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT32_2 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX21_GENERIC_NBIT32_2;

architecture SYN_structural of MUX21_GENERIC_NBIT32_2 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX21_425
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_426
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_427
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_428
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_429
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_430
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_431
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_432
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_433
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_434
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_435
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_436
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_437
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_438
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_439
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_440
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_441
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_442
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_443
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_444
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_445
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_446
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_447
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_448
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_449
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_450
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_451
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_452
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_453
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_454
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_455
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_456
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   MUXES_0 : MUX21_456 port map( A => A(0), B => B(0), S => n1, Y => Y(0));
   MUXES_1 : MUX21_455 port map( A => A(1), B => B(1), S => n1, Y => Y(1));
   MUXES_2 : MUX21_454 port map( A => A(2), B => B(2), S => n1, Y => Y(2));
   MUXES_3 : MUX21_453 port map( A => A(3), B => B(3), S => n1, Y => Y(3));
   MUXES_4 : MUX21_452 port map( A => A(4), B => B(4), S => n1, Y => Y(4));
   MUXES_5 : MUX21_451 port map( A => A(5), B => B(5), S => n1, Y => Y(5));
   MUXES_6 : MUX21_450 port map( A => A(6), B => B(6), S => n1, Y => Y(6));
   MUXES_7 : MUX21_449 port map( A => A(7), B => B(7), S => n1, Y => Y(7));
   MUXES_8 : MUX21_448 port map( A => A(8), B => B(8), S => n1, Y => Y(8));
   MUXES_9 : MUX21_447 port map( A => A(9), B => B(9), S => n1, Y => Y(9));
   MUXES_10 : MUX21_446 port map( A => A(10), B => B(10), S => n1, Y => Y(10));
   MUXES_11 : MUX21_445 port map( A => A(11), B => B(11), S => n1, Y => Y(11));
   MUXES_12 : MUX21_444 port map( A => A(12), B => B(12), S => n2, Y => Y(12));
   MUXES_13 : MUX21_443 port map( A => A(13), B => B(13), S => n2, Y => Y(13));
   MUXES_14 : MUX21_442 port map( A => A(14), B => B(14), S => n2, Y => Y(14));
   MUXES_15 : MUX21_441 port map( A => A(15), B => B(15), S => n2, Y => Y(15));
   MUXES_16 : MUX21_440 port map( A => A(16), B => B(16), S => n2, Y => Y(16));
   MUXES_17 : MUX21_439 port map( A => A(17), B => B(17), S => n2, Y => Y(17));
   MUXES_18 : MUX21_438 port map( A => A(18), B => B(18), S => n2, Y => Y(18));
   MUXES_19 : MUX21_437 port map( A => A(19), B => B(19), S => n2, Y => Y(19));
   MUXES_20 : MUX21_436 port map( A => A(20), B => B(20), S => n2, Y => Y(20));
   MUXES_21 : MUX21_435 port map( A => A(21), B => B(21), S => n2, Y => Y(21));
   MUXES_22 : MUX21_434 port map( A => A(22), B => B(22), S => n2, Y => Y(22));
   MUXES_23 : MUX21_433 port map( A => A(23), B => B(23), S => n2, Y => Y(23));
   MUXES_24 : MUX21_432 port map( A => A(24), B => B(24), S => n3, Y => Y(24));
   MUXES_25 : MUX21_431 port map( A => A(25), B => B(25), S => n3, Y => Y(25));
   MUXES_26 : MUX21_430 port map( A => A(26), B => B(26), S => n3, Y => Y(26));
   MUXES_27 : MUX21_429 port map( A => A(27), B => B(27), S => n3, Y => Y(27));
   MUXES_28 : MUX21_428 port map( A => A(28), B => B(28), S => n3, Y => Y(28));
   MUXES_29 : MUX21_427 port map( A => A(29), B => B(29), S => n3, Y => Y(29));
   MUXES_30 : MUX21_426 port map( A => A(30), B => B(30), S => n3, Y => Y(30));
   MUXES_31 : MUX21_425 port map( A => A(31), B => B(31), S => n3, Y => Y(31));
   U1 : BUF_X1 port map( A => SEL, Z => n1);
   U2 : BUF_X1 port map( A => SEL, Z => n2);
   U3 : BUF_X1 port map( A => SEL, Z => n3);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT32_1 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX21_GENERIC_NBIT32_1;

architecture SYN_structural of MUX21_GENERIC_NBIT32_1 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX21_393
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_394
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_395
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_396
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_397
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_398
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_399
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_400
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_401
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_402
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_403
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_404
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_405
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_406
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_407
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_408
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_409
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_410
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_411
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_412
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_413
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_414
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_415
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_416
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_417
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_418
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_419
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_420
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_421
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_422
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_423
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_424
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   MUXES_0 : MUX21_424 port map( A => A(0), B => B(0), S => n1, Y => Y(0));
   MUXES_1 : MUX21_423 port map( A => A(1), B => B(1), S => n1, Y => Y(1));
   MUXES_2 : MUX21_422 port map( A => A(2), B => B(2), S => n1, Y => Y(2));
   MUXES_3 : MUX21_421 port map( A => A(3), B => B(3), S => n1, Y => Y(3));
   MUXES_4 : MUX21_420 port map( A => A(4), B => B(4), S => n1, Y => Y(4));
   MUXES_5 : MUX21_419 port map( A => A(5), B => B(5), S => n1, Y => Y(5));
   MUXES_6 : MUX21_418 port map( A => A(6), B => B(6), S => n1, Y => Y(6));
   MUXES_7 : MUX21_417 port map( A => A(7), B => B(7), S => n1, Y => Y(7));
   MUXES_8 : MUX21_416 port map( A => A(8), B => B(8), S => n1, Y => Y(8));
   MUXES_9 : MUX21_415 port map( A => A(9), B => B(9), S => n1, Y => Y(9));
   MUXES_10 : MUX21_414 port map( A => A(10), B => B(10), S => n1, Y => Y(10));
   MUXES_11 : MUX21_413 port map( A => A(11), B => B(11), S => n1, Y => Y(11));
   MUXES_12 : MUX21_412 port map( A => A(12), B => B(12), S => n2, Y => Y(12));
   MUXES_13 : MUX21_411 port map( A => A(13), B => B(13), S => n2, Y => Y(13));
   MUXES_14 : MUX21_410 port map( A => A(14), B => B(14), S => n2, Y => Y(14));
   MUXES_15 : MUX21_409 port map( A => A(15), B => B(15), S => n2, Y => Y(15));
   MUXES_16 : MUX21_408 port map( A => A(16), B => B(16), S => n2, Y => Y(16));
   MUXES_17 : MUX21_407 port map( A => A(17), B => B(17), S => n2, Y => Y(17));
   MUXES_18 : MUX21_406 port map( A => A(18), B => B(18), S => n2, Y => Y(18));
   MUXES_19 : MUX21_405 port map( A => A(19), B => B(19), S => n2, Y => Y(19));
   MUXES_20 : MUX21_404 port map( A => A(20), B => B(20), S => n2, Y => Y(20));
   MUXES_21 : MUX21_403 port map( A => A(21), B => B(21), S => n2, Y => Y(21));
   MUXES_22 : MUX21_402 port map( A => A(22), B => B(22), S => n2, Y => Y(22));
   MUXES_23 : MUX21_401 port map( A => A(23), B => B(23), S => n2, Y => Y(23));
   MUXES_24 : MUX21_400 port map( A => A(24), B => B(24), S => n3, Y => Y(24));
   MUXES_25 : MUX21_399 port map( A => A(25), B => B(25), S => n3, Y => Y(25));
   MUXES_26 : MUX21_398 port map( A => A(26), B => B(26), S => n3, Y => Y(26));
   MUXES_27 : MUX21_397 port map( A => A(27), B => B(27), S => n3, Y => Y(27));
   MUXES_28 : MUX21_396 port map( A => A(28), B => B(28), S => n3, Y => Y(28));
   MUXES_29 : MUX21_395 port map( A => A(29), B => B(29), S => n3, Y => Y(29));
   MUXES_30 : MUX21_394 port map( A => A(30), B => B(30), S => n3, Y => Y(30));
   MUXES_31 : MUX21_393 port map( A => A(31), B => B(31), S => n3, Y => Y(31));
   U1 : BUF_X1 port map( A => SEL, Z => n2);
   U2 : BUF_X1 port map( A => SEL, Z => n1);
   U3 : BUF_X1 port map( A => SEL, Z => n3);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX81_0 is

   port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
         downto 0);  Y : out std_logic);

end MUX81_0;

architecture SYN_BEHAVIORAL_1 of MUX81_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n1
      , n2, n3, n4, n5, n6 : std_logic;

begin
   
   U20 : NAND3_X1 port map( A1 => S(1), A2 => n6, A3 => H, ZN => n19);
   U21 : NAND3_X1 port map( A1 => S(0), A2 => n2, A3 => F, ZN => n17);
   U1 : INV_X1 port map( A => n15, ZN => n5);
   U2 : NOR2_X1 port map( A1 => n1, A2 => S(2), ZN => n15);
   U3 : INV_X1 port map( A => n10, ZN => n4);
   U4 : INV_X1 port map( A => n20, ZN => n6);
   U5 : NAND2_X1 port map( A1 => n7, A2 => n8, ZN => Y);
   U6 : NAND4_X1 port map( A1 => A, A2 => n1, A3 => n2, A4 => n3, ZN => n8);
   U7 : AOI22_X1 port map( A1 => n9, A2 => n4, B1 => B, B2 => n10, ZN => n7);
   U8 : OAI21_X1 port map( B1 => n11, B2 => n12, A => n13, ZN => n9);
   U9 : NAND2_X1 port map( A1 => C, A2 => n12, ZN => n13);
   U10 : AOI22_X1 port map( A1 => n14, A2 => n5, B1 => D, B2 => n15, ZN => n11)
                           ;
   U11 : NOR3_X1 port map( A1 => S(0), A2 => S(2), A3 => n2, ZN => n12);
   U12 : NAND4_X1 port map( A1 => n16, A2 => n17, A3 => n18, A4 => n19, ZN => 
                           n14);
   U13 : NAND4_X1 port map( A1 => E, A2 => S(2), A3 => n1, A4 => n2, ZN => n16)
                           ;
   U14 : NAND2_X1 port map( A1 => G, A2 => n20, ZN => n18);
   U15 : NOR3_X1 port map( A1 => S(1), A2 => S(2), A3 => n1, ZN => n10);
   U16 : NOR2_X1 port map( A1 => n2, A2 => S(0), ZN => n20);
   U17 : INV_X1 port map( A => S(0), ZN => n1);
   U18 : INV_X1 port map( A => S(1), ZN => n2);
   U19 : INV_X1 port map( A => S(2), ZN => n3);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_GENERIC_NBIT8_0 is

   port( A, B, C, D : in std_logic_vector (7 downto 0);  SEL : in 
         std_logic_vector (1 downto 0);  Y : out std_logic_vector (7 downto 0)
         );

end MUX41_GENERIC_NBIT8_0;

architecture SYN_structural of MUX41_GENERIC_NBIT8_0 is

   component MUX41_25
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_26
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_27
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_28
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_29
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_30
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_31
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_32
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX41_32 port map( A => A(0), B => B(0), C => C(0), D => D(0), 
                           S(1) => SEL(1), S(0) => SEL(0), Y => Y(0));
   MUXES_1 : MUX41_31 port map( A => A(1), B => B(1), C => C(1), D => D(1), 
                           S(1) => SEL(1), S(0) => SEL(0), Y => Y(1));
   MUXES_2 : MUX41_30 port map( A => A(2), B => B(2), C => C(2), D => D(2), 
                           S(1) => SEL(1), S(0) => SEL(0), Y => Y(2));
   MUXES_3 : MUX41_29 port map( A => A(3), B => B(3), C => C(3), D => D(3), 
                           S(1) => SEL(1), S(0) => SEL(0), Y => Y(3));
   MUXES_4 : MUX41_28 port map( A => A(4), B => B(4), C => C(4), D => D(4), 
                           S(1) => SEL(1), S(0) => SEL(0), Y => Y(4));
   MUXES_5 : MUX41_27 port map( A => A(5), B => B(5), C => C(5), D => D(5), 
                           S(1) => SEL(1), S(0) => SEL(0), Y => Y(5));
   MUXES_6 : MUX41_26 port map( A => A(6), B => B(6), C => C(6), D => D(6), 
                           S(1) => SEL(1), S(0) => SEL(0), Y => Y(6));
   MUXES_7 : MUX41_25 port map( A => A(7), B => B(7), C => C(7), D => D(7), 
                           S(1) => SEL(1), S(0) => SEL(0), Y => Y(7));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT8_0 is

   port( A, B : in std_logic_vector (7 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (7 downto 0));

end MUX21_GENERIC_NBIT8_0;

architecture SYN_structural of MUX21_GENERIC_NBIT8_0 is

   component MUX21_353
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_354
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_355
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_356
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_357
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_358
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_359
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_360
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_360 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_359 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_358 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_357 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));
   MUXES_4 : MUX21_356 port map( A => A(4), B => B(4), S => SEL, Y => Y(4));
   MUXES_5 : MUX21_355 port map( A => A(5), B => B(5), S => SEL, Y => Y(5));
   MUXES_6 : MUX21_354 port map( A => A(6), B => B(6), S => SEL, Y => Y(6));
   MUXES_7 : MUX21_353 port map( A => A(7), B => B(7), S => SEL, Y => Y(7));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FA_0 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_0;

architecture SYN_BEHAVIORAL of FA_0 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => Ci, B => n2, Z => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => Co);
   U2 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n2, B2 => Ci, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity sum_generator_n_bit64_n_CSB16_0 is

   port( A, B : in std_logic_vector (63 downto 0);  C_in : in std_logic_vector 
         (15 downto 0);  S : out std_logic_vector (63 downto 0));

end sum_generator_n_bit64_n_CSB16_0;

architecture SYN_STRUCTURAL of sum_generator_n_bit64_n_CSB16_0 is

   component carry_select_block_n4_33
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_n4_34
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_n4_35
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_n4_36
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_n4_37
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_n4_38
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_n4_39
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_n4_40
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_n4_41
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_n4_42
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_n4_43
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_n4_44
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_n4_45
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_n4_46
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_n4_47
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_n4_48
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;

begin
   
   csb_0 : carry_select_block_n4_48 port map( A(3) => A(3), A(2) => A(2), A(1) 
                           => A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), 
                           B(1) => B(1), B(0) => B(0), C_sel => C_in(0), S(3) 
                           => S(3), S(2) => S(2), S(1) => S(1), S(0) => S(0));
   csb_1 : carry_select_block_n4_47 port map( A(3) => A(7), A(2) => A(6), A(1) 
                           => A(5), A(0) => A(4), B(3) => B(7), B(2) => B(6), 
                           B(1) => B(5), B(0) => B(4), C_sel => C_in(1), S(3) 
                           => S(7), S(2) => S(6), S(1) => S(5), S(0) => S(4));
   csb_2 : carry_select_block_n4_46 port map( A(3) => A(11), A(2) => A(10), 
                           A(1) => A(9), A(0) => A(8), B(3) => B(11), B(2) => 
                           B(10), B(1) => B(9), B(0) => B(8), C_sel => C_in(2),
                           S(3) => S(11), S(2) => S(10), S(1) => S(9), S(0) => 
                           S(8));
   csb_3 : carry_select_block_n4_45 port map( A(3) => A(15), A(2) => A(14), 
                           A(1) => A(13), A(0) => A(12), B(3) => B(15), B(2) =>
                           B(14), B(1) => B(13), B(0) => B(12), C_sel => 
                           C_in(3), S(3) => S(15), S(2) => S(14), S(1) => S(13)
                           , S(0) => S(12));
   csb_4 : carry_select_block_n4_44 port map( A(3) => A(19), A(2) => A(18), 
                           A(1) => A(17), A(0) => A(16), B(3) => B(19), B(2) =>
                           B(18), B(1) => B(17), B(0) => B(16), C_sel => 
                           C_in(4), S(3) => S(19), S(2) => S(18), S(1) => S(17)
                           , S(0) => S(16));
   csb_5 : carry_select_block_n4_43 port map( A(3) => A(23), A(2) => A(22), 
                           A(1) => A(21), A(0) => A(20), B(3) => B(23), B(2) =>
                           B(22), B(1) => B(21), B(0) => B(20), C_sel => 
                           C_in(5), S(3) => S(23), S(2) => S(22), S(1) => S(21)
                           , S(0) => S(20));
   csb_6 : carry_select_block_n4_42 port map( A(3) => A(27), A(2) => A(26), 
                           A(1) => A(25), A(0) => A(24), B(3) => B(27), B(2) =>
                           B(26), B(1) => B(25), B(0) => B(24), C_sel => 
                           C_in(6), S(3) => S(27), S(2) => S(26), S(1) => S(25)
                           , S(0) => S(24));
   csb_7 : carry_select_block_n4_41 port map( A(3) => A(31), A(2) => A(30), 
                           A(1) => A(29), A(0) => A(28), B(3) => B(31), B(2) =>
                           B(30), B(1) => B(29), B(0) => B(28), C_sel => 
                           C_in(7), S(3) => S(31), S(2) => S(30), S(1) => S(29)
                           , S(0) => S(28));
   csb_8 : carry_select_block_n4_40 port map( A(3) => A(35), A(2) => A(34), 
                           A(1) => A(33), A(0) => A(32), B(3) => B(35), B(2) =>
                           B(34), B(1) => B(33), B(0) => B(32), C_sel => 
                           C_in(8), S(3) => S(35), S(2) => S(34), S(1) => S(33)
                           , S(0) => S(32));
   csb_9 : carry_select_block_n4_39 port map( A(3) => A(39), A(2) => A(38), 
                           A(1) => A(37), A(0) => A(36), B(3) => B(39), B(2) =>
                           B(38), B(1) => B(37), B(0) => B(36), C_sel => 
                           C_in(9), S(3) => S(39), S(2) => S(38), S(1) => S(37)
                           , S(0) => S(36));
   csb_10 : carry_select_block_n4_38 port map( A(3) => A(43), A(2) => A(42), 
                           A(1) => A(41), A(0) => A(40), B(3) => B(43), B(2) =>
                           B(42), B(1) => B(41), B(0) => B(40), C_sel => 
                           C_in(10), S(3) => S(43), S(2) => S(42), S(1) => 
                           S(41), S(0) => S(40));
   csb_11 : carry_select_block_n4_37 port map( A(3) => A(47), A(2) => A(46), 
                           A(1) => A(45), A(0) => A(44), B(3) => B(47), B(2) =>
                           B(46), B(1) => B(45), B(0) => B(44), C_sel => 
                           C_in(11), S(3) => S(47), S(2) => S(46), S(1) => 
                           S(45), S(0) => S(44));
   csb_12 : carry_select_block_n4_36 port map( A(3) => A(51), A(2) => A(50), 
                           A(1) => A(49), A(0) => A(48), B(3) => B(51), B(2) =>
                           B(50), B(1) => B(49), B(0) => B(48), C_sel => 
                           C_in(12), S(3) => S(51), S(2) => S(50), S(1) => 
                           S(49), S(0) => S(48));
   csb_13 : carry_select_block_n4_35 port map( A(3) => A(55), A(2) => A(54), 
                           A(1) => A(53), A(0) => A(52), B(3) => B(55), B(2) =>
                           B(54), B(1) => B(53), B(0) => B(52), C_sel => 
                           C_in(13), S(3) => S(55), S(2) => S(54), S(1) => 
                           S(53), S(0) => S(52));
   csb_14 : carry_select_block_n4_34 port map( A(3) => A(59), A(2) => A(58), 
                           A(1) => A(57), A(0) => A(56), B(3) => B(59), B(2) =>
                           B(58), B(1) => B(57), B(0) => B(56), C_sel => 
                           C_in(14), S(3) => S(59), S(2) => S(58), S(1) => 
                           S(57), S(0) => S(56));
   csb_15 : carry_select_block_n4_33 port map( A(3) => A(63), A(2) => A(62), 
                           A(1) => A(61), A(0) => A(60), B(3) => B(63), B(2) =>
                           B(62), B(1) => B(61), B(0) => B(60), C_sel => 
                           C_in(15), S(3) => S(63), S(2) => S(62), S(1) => 
                           S(61), S(0) => S(60));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity CARRY_GENERATOR_NBIT64_NBIT_PER_BLOCK4_0 is

   port( A, B : in std_logic_vector (63 downto 0);  Cin : in std_logic;  Co : 
         out std_logic_vector (15 downto 0));

end CARRY_GENERATOR_NBIT64_NBIT_PER_BLOCK4_0;

architecture SYN_structural of CARRY_GENERATOR_NBIT64_NBIT_PER_BLOCK4_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component G_BLOCK_35
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component G_BLOCK_36
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component G_BLOCK_37
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component G_BLOCK_38
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component G_BLOCK_39
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component G_BLOCK_40
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component G_BLOCK_41
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component G_BLOCK_42
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component G_BLOCK_43
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component G_BLOCK_44
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component G_BLOCK_45
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component G_BLOCK_46
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component PG_BLOCK_127
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_128
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_129
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_130
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component G_BLOCK_47
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component G_BLOCK_48
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component PG_BLOCK_131
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_132
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_133
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_134
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_135
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_136
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component G_BLOCK_49
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component PG_BLOCK_137
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_138
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_139
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_140
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_141
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_142
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_143
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component G_BLOCK_50
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component PG_BLOCK_144
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_145
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_146
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_147
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_148
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_149
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_150
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_151
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_152
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_153
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_154
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_155
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_156
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_157
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_158
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component G_BLOCK_51
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component PG_BLOCK_159
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_160
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_161
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_162
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_163
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_164
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_165
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_166
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_167
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_168
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_169
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_170
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_171
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_172
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_173
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_174
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_175
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_176
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_177
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_178
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_179
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_180
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_181
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_182
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_183
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_184
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_185
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_186
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_187
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_188
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_189
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component pg_net_127
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_128
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_129
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_130
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_131
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_132
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_133
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_134
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_135
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_136
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_137
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_138
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_139
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_140
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_141
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_142
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_143
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_144
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_145
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_146
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_147
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_148
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_149
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_150
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_151
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_152
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_153
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_154
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_155
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_156
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_157
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_158
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_159
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_160
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_161
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_162
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_163
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_164
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_165
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_166
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_167
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_168
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_169
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_170
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_171
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_172
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_173
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_174
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_175
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_176
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_177
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_178
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_179
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_180
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_181
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_182
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_183
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_184
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_185
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_186
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_187
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_188
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_189
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   signal Co_15_port, Co_14_port, Co_13_port, Co_12_port, Co_11_port, 
      Co_10_port, Co_9_port, Co_8_port, Co_7_port, Co_6_port, Co_5_port, 
      Co_4_port, Co_3_port, Co_2_port, Co_1_port, Co_0_port, g_vector_5_63_port
      , g_vector_5_59_port, g_vector_5_55_port, g_vector_5_51_port, 
      g_vector_4_63_port, g_vector_4_59_port, g_vector_4_47_port, 
      g_vector_4_43_port, g_vector_4_31_port, g_vector_4_27_port, 
      g_vector_3_63_port, g_vector_3_55_port, g_vector_3_47_port, 
      g_vector_3_39_port, g_vector_3_31_port, g_vector_3_23_port, 
      g_vector_3_15_port, g_vector_2_63_port, g_vector_2_59_port, 
      g_vector_2_55_port, g_vector_2_51_port, g_vector_2_47_port, 
      g_vector_2_43_port, g_vector_2_39_port, g_vector_2_35_port, 
      g_vector_2_31_port, g_vector_2_27_port, g_vector_2_23_port, 
      g_vector_2_19_port, g_vector_2_15_port, g_vector_2_11_port, 
      g_vector_2_7_port, g_vector_1_63_port, g_vector_1_61_port, 
      g_vector_1_59_port, g_vector_1_57_port, g_vector_1_55_port, 
      g_vector_1_53_port, g_vector_1_51_port, g_vector_1_49_port, 
      g_vector_1_47_port, g_vector_1_45_port, g_vector_1_43_port, 
      g_vector_1_41_port, g_vector_1_39_port, g_vector_1_37_port, 
      g_vector_1_35_port, g_vector_1_33_port, g_vector_1_31_port, 
      g_vector_1_29_port, g_vector_1_27_port, g_vector_1_25_port, 
      g_vector_1_23_port, g_vector_1_21_port, g_vector_1_19_port, 
      g_vector_1_17_port, g_vector_1_15_port, g_vector_1_13_port, 
      g_vector_1_11_port, g_vector_1_9_port, g_vector_1_7_port, 
      g_vector_1_5_port, g_vector_1_3_port, g_vector_1_1_port, 
      g_vector_0_63_port, g_vector_0_62_port, g_vector_0_61_port, 
      g_vector_0_60_port, g_vector_0_59_port, g_vector_0_58_port, 
      g_vector_0_57_port, g_vector_0_56_port, g_vector_0_55_port, 
      g_vector_0_54_port, g_vector_0_53_port, g_vector_0_52_port, 
      g_vector_0_51_port, g_vector_0_50_port, g_vector_0_49_port, 
      g_vector_0_48_port, g_vector_0_47_port, g_vector_0_46_port, 
      g_vector_0_45_port, g_vector_0_44_port, g_vector_0_43_port, 
      g_vector_0_42_port, g_vector_0_41_port, g_vector_0_40_port, 
      g_vector_0_39_port, g_vector_0_38_port, g_vector_0_37_port, 
      g_vector_0_36_port, g_vector_0_35_port, g_vector_0_34_port, 
      g_vector_0_33_port, g_vector_0_32_port, g_vector_0_31_port, 
      g_vector_0_30_port, g_vector_0_29_port, g_vector_0_28_port, 
      g_vector_0_27_port, g_vector_0_26_port, g_vector_0_25_port, 
      g_vector_0_24_port, g_vector_0_23_port, g_vector_0_22_port, 
      g_vector_0_21_port, g_vector_0_20_port, g_vector_0_19_port, 
      g_vector_0_18_port, g_vector_0_17_port, g_vector_0_16_port, 
      g_vector_0_15_port, g_vector_0_14_port, g_vector_0_13_port, 
      g_vector_0_12_port, g_vector_0_11_port, g_vector_0_10_port, 
      g_vector_0_9_port, g_vector_0_8_port, g_vector_0_7_port, 
      g_vector_0_6_port, g_vector_0_5_port, g_vector_0_4_port, 
      g_vector_0_3_port, g_vector_0_2_port, g_vector_0_1_port, 
      g_vector_0_0_port, p_vector_5_63_port, p_vector_5_59_port, 
      p_vector_5_55_port, p_vector_5_51_port, p_vector_4_63_port, 
      p_vector_4_59_port, p_vector_4_47_port, p_vector_4_43_port, 
      p_vector_4_31_port, p_vector_4_27_port, p_vector_3_63_port, 
      p_vector_3_55_port, p_vector_3_47_port, p_vector_3_39_port, 
      p_vector_3_31_port, p_vector_3_23_port, p_vector_3_15_port, 
      p_vector_2_63_port, p_vector_2_59_port, p_vector_2_55_port, 
      p_vector_2_51_port, p_vector_2_47_port, p_vector_2_43_port, 
      p_vector_2_39_port, p_vector_2_35_port, p_vector_2_31_port, 
      p_vector_2_27_port, p_vector_2_23_port, p_vector_2_19_port, 
      p_vector_2_15_port, p_vector_2_11_port, p_vector_2_7_port, 
      p_vector_1_63_port, p_vector_1_61_port, p_vector_1_59_port, 
      p_vector_1_57_port, p_vector_1_55_port, p_vector_1_53_port, 
      p_vector_1_51_port, p_vector_1_49_port, p_vector_1_47_port, 
      p_vector_1_45_port, p_vector_1_43_port, p_vector_1_41_port, 
      p_vector_1_39_port, p_vector_1_37_port, p_vector_1_35_port, 
      p_vector_1_33_port, p_vector_1_31_port, p_vector_1_29_port, 
      p_vector_1_27_port, p_vector_1_25_port, p_vector_1_23_port, 
      p_vector_1_21_port, p_vector_1_19_port, p_vector_1_17_port, 
      p_vector_1_15_port, p_vector_1_13_port, p_vector_1_11_port, 
      p_vector_1_9_port, p_vector_1_7_port, p_vector_1_5_port, 
      p_vector_1_3_port, p_vector_0_63_port, p_vector_0_62_port, 
      p_vector_0_61_port, p_vector_0_60_port, p_vector_0_59_port, 
      p_vector_0_58_port, p_vector_0_57_port, p_vector_0_56_port, 
      p_vector_0_55_port, p_vector_0_54_port, p_vector_0_53_port, 
      p_vector_0_52_port, p_vector_0_51_port, p_vector_0_50_port, 
      p_vector_0_49_port, p_vector_0_48_port, p_vector_0_47_port, 
      p_vector_0_46_port, p_vector_0_45_port, p_vector_0_44_port, 
      p_vector_0_43_port, p_vector_0_42_port, p_vector_0_41_port, 
      p_vector_0_40_port, p_vector_0_39_port, p_vector_0_38_port, 
      p_vector_0_37_port, p_vector_0_36_port, p_vector_0_35_port, 
      p_vector_0_34_port, p_vector_0_33_port, p_vector_0_32_port, 
      p_vector_0_31_port, p_vector_0_30_port, p_vector_0_29_port, 
      p_vector_0_28_port, p_vector_0_27_port, p_vector_0_26_port, 
      p_vector_0_25_port, p_vector_0_24_port, p_vector_0_23_port, 
      p_vector_0_22_port, p_vector_0_21_port, p_vector_0_20_port, 
      p_vector_0_19_port, p_vector_0_18_port, p_vector_0_17_port, 
      p_vector_0_16_port, p_vector_0_15_port, p_vector_0_14_port, 
      p_vector_0_13_port, p_vector_0_12_port, p_vector_0_11_port, 
      p_vector_0_10_port, p_vector_0_9_port, p_vector_0_8_port, 
      p_vector_0_7_port, p_vector_0_6_port, p_vector_0_5_port, 
      p_vector_0_4_port, p_vector_0_3_port, p_vector_0_2_port, 
      p_vector_0_1_port, n3, n1, n2 : std_logic;

begin
   Co <= ( Co_15_port, Co_14_port, Co_13_port, Co_12_port, Co_11_port, 
      Co_10_port, Co_9_port, Co_8_port, Co_7_port, Co_6_port, Co_5_port, 
      Co_4_port, Co_3_port, Co_2_port, Co_1_port, Co_0_port );
   
   pg_network_63 : pg_net_189 port map( a => A(63), b => B(63), p => 
                           p_vector_0_63_port, g => g_vector_0_63_port);
   pg_network_62 : pg_net_188 port map( a => A(62), b => B(62), p => 
                           p_vector_0_62_port, g => g_vector_0_62_port);
   pg_network_61 : pg_net_187 port map( a => A(61), b => B(61), p => 
                           p_vector_0_61_port, g => g_vector_0_61_port);
   pg_network_60 : pg_net_186 port map( a => A(60), b => B(60), p => 
                           p_vector_0_60_port, g => g_vector_0_60_port);
   pg_network_59 : pg_net_185 port map( a => A(59), b => B(59), p => 
                           p_vector_0_59_port, g => g_vector_0_59_port);
   pg_network_58 : pg_net_184 port map( a => A(58), b => B(58), p => 
                           p_vector_0_58_port, g => g_vector_0_58_port);
   pg_network_57 : pg_net_183 port map( a => A(57), b => B(57), p => 
                           p_vector_0_57_port, g => g_vector_0_57_port);
   pg_network_56 : pg_net_182 port map( a => A(56), b => B(56), p => 
                           p_vector_0_56_port, g => g_vector_0_56_port);
   pg_network_55 : pg_net_181 port map( a => A(55), b => B(55), p => 
                           p_vector_0_55_port, g => g_vector_0_55_port);
   pg_network_54 : pg_net_180 port map( a => A(54), b => B(54), p => 
                           p_vector_0_54_port, g => g_vector_0_54_port);
   pg_network_53 : pg_net_179 port map( a => A(53), b => B(53), p => 
                           p_vector_0_53_port, g => g_vector_0_53_port);
   pg_network_52 : pg_net_178 port map( a => A(52), b => B(52), p => 
                           p_vector_0_52_port, g => g_vector_0_52_port);
   pg_network_51 : pg_net_177 port map( a => A(51), b => B(51), p => 
                           p_vector_0_51_port, g => g_vector_0_51_port);
   pg_network_50 : pg_net_176 port map( a => A(50), b => B(50), p => 
                           p_vector_0_50_port, g => g_vector_0_50_port);
   pg_network_49 : pg_net_175 port map( a => A(49), b => B(49), p => 
                           p_vector_0_49_port, g => g_vector_0_49_port);
   pg_network_48 : pg_net_174 port map( a => A(48), b => B(48), p => 
                           p_vector_0_48_port, g => g_vector_0_48_port);
   pg_network_47 : pg_net_173 port map( a => A(47), b => B(47), p => 
                           p_vector_0_47_port, g => g_vector_0_47_port);
   pg_network_46 : pg_net_172 port map( a => A(46), b => B(46), p => 
                           p_vector_0_46_port, g => g_vector_0_46_port);
   pg_network_45 : pg_net_171 port map( a => A(45), b => B(45), p => 
                           p_vector_0_45_port, g => g_vector_0_45_port);
   pg_network_44 : pg_net_170 port map( a => A(44), b => B(44), p => 
                           p_vector_0_44_port, g => g_vector_0_44_port);
   pg_network_43 : pg_net_169 port map( a => A(43), b => B(43), p => 
                           p_vector_0_43_port, g => g_vector_0_43_port);
   pg_network_42 : pg_net_168 port map( a => A(42), b => B(42), p => 
                           p_vector_0_42_port, g => g_vector_0_42_port);
   pg_network_41 : pg_net_167 port map( a => A(41), b => B(41), p => 
                           p_vector_0_41_port, g => g_vector_0_41_port);
   pg_network_40 : pg_net_166 port map( a => A(40), b => B(40), p => 
                           p_vector_0_40_port, g => g_vector_0_40_port);
   pg_network_39 : pg_net_165 port map( a => A(39), b => B(39), p => 
                           p_vector_0_39_port, g => g_vector_0_39_port);
   pg_network_38 : pg_net_164 port map( a => A(38), b => B(38), p => 
                           p_vector_0_38_port, g => g_vector_0_38_port);
   pg_network_37 : pg_net_163 port map( a => A(37), b => B(37), p => 
                           p_vector_0_37_port, g => g_vector_0_37_port);
   pg_network_36 : pg_net_162 port map( a => A(36), b => B(36), p => 
                           p_vector_0_36_port, g => g_vector_0_36_port);
   pg_network_35 : pg_net_161 port map( a => A(35), b => B(35), p => 
                           p_vector_0_35_port, g => g_vector_0_35_port);
   pg_network_34 : pg_net_160 port map( a => A(34), b => B(34), p => 
                           p_vector_0_34_port, g => g_vector_0_34_port);
   pg_network_33 : pg_net_159 port map( a => A(33), b => B(33), p => 
                           p_vector_0_33_port, g => g_vector_0_33_port);
   pg_network_32 : pg_net_158 port map( a => A(32), b => B(32), p => 
                           p_vector_0_32_port, g => g_vector_0_32_port);
   pg_network_31 : pg_net_157 port map( a => A(31), b => B(31), p => 
                           p_vector_0_31_port, g => g_vector_0_31_port);
   pg_network_30 : pg_net_156 port map( a => A(30), b => B(30), p => 
                           p_vector_0_30_port, g => g_vector_0_30_port);
   pg_network_29 : pg_net_155 port map( a => A(29), b => B(29), p => 
                           p_vector_0_29_port, g => g_vector_0_29_port);
   pg_network_28 : pg_net_154 port map( a => A(28), b => B(28), p => 
                           p_vector_0_28_port, g => g_vector_0_28_port);
   pg_network_27 : pg_net_153 port map( a => A(27), b => B(27), p => 
                           p_vector_0_27_port, g => g_vector_0_27_port);
   pg_network_26 : pg_net_152 port map( a => A(26), b => B(26), p => 
                           p_vector_0_26_port, g => g_vector_0_26_port);
   pg_network_25 : pg_net_151 port map( a => A(25), b => B(25), p => 
                           p_vector_0_25_port, g => g_vector_0_25_port);
   pg_network_24 : pg_net_150 port map( a => A(24), b => B(24), p => 
                           p_vector_0_24_port, g => g_vector_0_24_port);
   pg_network_23 : pg_net_149 port map( a => A(23), b => B(23), p => 
                           p_vector_0_23_port, g => g_vector_0_23_port);
   pg_network_22 : pg_net_148 port map( a => A(22), b => B(22), p => 
                           p_vector_0_22_port, g => g_vector_0_22_port);
   pg_network_21 : pg_net_147 port map( a => A(21), b => B(21), p => 
                           p_vector_0_21_port, g => g_vector_0_21_port);
   pg_network_20 : pg_net_146 port map( a => A(20), b => B(20), p => 
                           p_vector_0_20_port, g => g_vector_0_20_port);
   pg_network_19 : pg_net_145 port map( a => A(19), b => B(19), p => 
                           p_vector_0_19_port, g => g_vector_0_19_port);
   pg_network_18 : pg_net_144 port map( a => A(18), b => B(18), p => 
                           p_vector_0_18_port, g => g_vector_0_18_port);
   pg_network_17 : pg_net_143 port map( a => A(17), b => B(17), p => 
                           p_vector_0_17_port, g => g_vector_0_17_port);
   pg_network_16 : pg_net_142 port map( a => A(16), b => B(16), p => 
                           p_vector_0_16_port, g => g_vector_0_16_port);
   pg_network_15 : pg_net_141 port map( a => A(15), b => B(15), p => 
                           p_vector_0_15_port, g => g_vector_0_15_port);
   pg_network_14 : pg_net_140 port map( a => A(14), b => B(14), p => 
                           p_vector_0_14_port, g => g_vector_0_14_port);
   pg_network_13 : pg_net_139 port map( a => A(13), b => B(13), p => 
                           p_vector_0_13_port, g => g_vector_0_13_port);
   pg_network_12 : pg_net_138 port map( a => A(12), b => B(12), p => 
                           p_vector_0_12_port, g => g_vector_0_12_port);
   pg_network_11 : pg_net_137 port map( a => A(11), b => B(11), p => 
                           p_vector_0_11_port, g => g_vector_0_11_port);
   pg_network_10 : pg_net_136 port map( a => A(10), b => B(10), p => 
                           p_vector_0_10_port, g => g_vector_0_10_port);
   pg_network_9 : pg_net_135 port map( a => A(9), b => B(9), p => 
                           p_vector_0_9_port, g => g_vector_0_9_port);
   pg_network_8 : pg_net_134 port map( a => A(8), b => B(8), p => 
                           p_vector_0_8_port, g => g_vector_0_8_port);
   pg_network_7 : pg_net_133 port map( a => A(7), b => B(7), p => 
                           p_vector_0_7_port, g => g_vector_0_7_port);
   pg_network_6 : pg_net_132 port map( a => A(6), b => B(6), p => 
                           p_vector_0_6_port, g => g_vector_0_6_port);
   pg_network_5 : pg_net_131 port map( a => A(5), b => B(5), p => 
                           p_vector_0_5_port, g => g_vector_0_5_port);
   pg_network_4 : pg_net_130 port map( a => A(4), b => B(4), p => 
                           p_vector_0_4_port, g => g_vector_0_4_port);
   pg_network_3 : pg_net_129 port map( a => A(3), b => B(3), p => 
                           p_vector_0_3_port, g => g_vector_0_3_port);
   pg_network_2 : pg_net_128 port map( a => A(2), b => B(2), p => 
                           p_vector_0_2_port, g => g_vector_0_2_port);
   pg_network_1 : pg_net_127 port map( a => A(1), b => B(1), p => 
                           p_vector_0_1_port, g => g_vector_0_1_port);
   std_PG_1_63 : PG_BLOCK_189 port map( p2 => p_vector_0_63_port, g2 => 
                           g_vector_0_63_port, p1 => p_vector_0_62_port, g1 => 
                           g_vector_0_62_port, PG_P => p_vector_1_63_port, PG_G
                           => g_vector_1_63_port);
   std_PG_1_61 : PG_BLOCK_188 port map( p2 => p_vector_0_61_port, g2 => 
                           g_vector_0_61_port, p1 => p_vector_0_60_port, g1 => 
                           g_vector_0_60_port, PG_P => p_vector_1_61_port, PG_G
                           => g_vector_1_61_port);
   std_PG_1_59 : PG_BLOCK_187 port map( p2 => p_vector_0_59_port, g2 => 
                           g_vector_0_59_port, p1 => p_vector_0_58_port, g1 => 
                           g_vector_0_58_port, PG_P => p_vector_1_59_port, PG_G
                           => g_vector_1_59_port);
   std_PG_1_57 : PG_BLOCK_186 port map( p2 => p_vector_0_57_port, g2 => 
                           g_vector_0_57_port, p1 => p_vector_0_56_port, g1 => 
                           g_vector_0_56_port, PG_P => p_vector_1_57_port, PG_G
                           => g_vector_1_57_port);
   std_PG_1_55 : PG_BLOCK_185 port map( p2 => p_vector_0_55_port, g2 => 
                           g_vector_0_55_port, p1 => p_vector_0_54_port, g1 => 
                           g_vector_0_54_port, PG_P => p_vector_1_55_port, PG_G
                           => g_vector_1_55_port);
   std_PG_1_53 : PG_BLOCK_184 port map( p2 => p_vector_0_53_port, g2 => 
                           g_vector_0_53_port, p1 => p_vector_0_52_port, g1 => 
                           g_vector_0_52_port, PG_P => p_vector_1_53_port, PG_G
                           => g_vector_1_53_port);
   std_PG_1_51 : PG_BLOCK_183 port map( p2 => p_vector_0_51_port, g2 => 
                           g_vector_0_51_port, p1 => p_vector_0_50_port, g1 => 
                           g_vector_0_50_port, PG_P => p_vector_1_51_port, PG_G
                           => g_vector_1_51_port);
   std_PG_1_49 : PG_BLOCK_182 port map( p2 => p_vector_0_49_port, g2 => 
                           g_vector_0_49_port, p1 => p_vector_0_48_port, g1 => 
                           g_vector_0_48_port, PG_P => p_vector_1_49_port, PG_G
                           => g_vector_1_49_port);
   std_PG_1_47 : PG_BLOCK_181 port map( p2 => p_vector_0_47_port, g2 => 
                           g_vector_0_47_port, p1 => p_vector_0_46_port, g1 => 
                           g_vector_0_46_port, PG_P => p_vector_1_47_port, PG_G
                           => g_vector_1_47_port);
   std_PG_1_45 : PG_BLOCK_180 port map( p2 => p_vector_0_45_port, g2 => 
                           g_vector_0_45_port, p1 => p_vector_0_44_port, g1 => 
                           g_vector_0_44_port, PG_P => p_vector_1_45_port, PG_G
                           => g_vector_1_45_port);
   std_PG_1_43 : PG_BLOCK_179 port map( p2 => p_vector_0_43_port, g2 => 
                           g_vector_0_43_port, p1 => p_vector_0_42_port, g1 => 
                           g_vector_0_42_port, PG_P => p_vector_1_43_port, PG_G
                           => g_vector_1_43_port);
   std_PG_1_41 : PG_BLOCK_178 port map( p2 => p_vector_0_41_port, g2 => 
                           g_vector_0_41_port, p1 => p_vector_0_40_port, g1 => 
                           g_vector_0_40_port, PG_P => p_vector_1_41_port, PG_G
                           => g_vector_1_41_port);
   std_PG_1_39 : PG_BLOCK_177 port map( p2 => p_vector_0_39_port, g2 => 
                           g_vector_0_39_port, p1 => p_vector_0_38_port, g1 => 
                           g_vector_0_38_port, PG_P => p_vector_1_39_port, PG_G
                           => g_vector_1_39_port);
   std_PG_1_37 : PG_BLOCK_176 port map( p2 => p_vector_0_37_port, g2 => 
                           g_vector_0_37_port, p1 => p_vector_0_36_port, g1 => 
                           g_vector_0_36_port, PG_P => p_vector_1_37_port, PG_G
                           => g_vector_1_37_port);
   std_PG_1_35 : PG_BLOCK_175 port map( p2 => p_vector_0_35_port, g2 => 
                           g_vector_0_35_port, p1 => p_vector_0_34_port, g1 => 
                           g_vector_0_34_port, PG_P => p_vector_1_35_port, PG_G
                           => g_vector_1_35_port);
   std_PG_1_33 : PG_BLOCK_174 port map( p2 => p_vector_0_33_port, g2 => 
                           g_vector_0_33_port, p1 => p_vector_0_32_port, g1 => 
                           g_vector_0_32_port, PG_P => p_vector_1_33_port, PG_G
                           => g_vector_1_33_port);
   std_PG_1_31 : PG_BLOCK_173 port map( p2 => p_vector_0_31_port, g2 => 
                           g_vector_0_31_port, p1 => p_vector_0_30_port, g1 => 
                           g_vector_0_30_port, PG_P => p_vector_1_31_port, PG_G
                           => g_vector_1_31_port);
   std_PG_1_29 : PG_BLOCK_172 port map( p2 => p_vector_0_29_port, g2 => 
                           g_vector_0_29_port, p1 => p_vector_0_28_port, g1 => 
                           g_vector_0_28_port, PG_P => p_vector_1_29_port, PG_G
                           => g_vector_1_29_port);
   std_PG_1_27 : PG_BLOCK_171 port map( p2 => p_vector_0_27_port, g2 => 
                           g_vector_0_27_port, p1 => p_vector_0_26_port, g1 => 
                           g_vector_0_26_port, PG_P => p_vector_1_27_port, PG_G
                           => g_vector_1_27_port);
   std_PG_1_25 : PG_BLOCK_170 port map( p2 => p_vector_0_25_port, g2 => 
                           g_vector_0_25_port, p1 => p_vector_0_24_port, g1 => 
                           g_vector_0_24_port, PG_P => p_vector_1_25_port, PG_G
                           => g_vector_1_25_port);
   std_PG_1_23 : PG_BLOCK_169 port map( p2 => p_vector_0_23_port, g2 => 
                           g_vector_0_23_port, p1 => p_vector_0_22_port, g1 => 
                           g_vector_0_22_port, PG_P => p_vector_1_23_port, PG_G
                           => g_vector_1_23_port);
   std_PG_1_21 : PG_BLOCK_168 port map( p2 => p_vector_0_21_port, g2 => 
                           g_vector_0_21_port, p1 => p_vector_0_20_port, g1 => 
                           g_vector_0_20_port, PG_P => p_vector_1_21_port, PG_G
                           => g_vector_1_21_port);
   std_PG_1_19 : PG_BLOCK_167 port map( p2 => p_vector_0_19_port, g2 => 
                           g_vector_0_19_port, p1 => p_vector_0_18_port, g1 => 
                           g_vector_0_18_port, PG_P => p_vector_1_19_port, PG_G
                           => g_vector_1_19_port);
   std_PG_1_17 : PG_BLOCK_166 port map( p2 => p_vector_0_17_port, g2 => 
                           g_vector_0_17_port, p1 => p_vector_0_16_port, g1 => 
                           g_vector_0_16_port, PG_P => p_vector_1_17_port, PG_G
                           => g_vector_1_17_port);
   std_PG_1_15 : PG_BLOCK_165 port map( p2 => p_vector_0_15_port, g2 => 
                           g_vector_0_15_port, p1 => p_vector_0_14_port, g1 => 
                           g_vector_0_14_port, PG_P => p_vector_1_15_port, PG_G
                           => g_vector_1_15_port);
   std_PG_1_13 : PG_BLOCK_164 port map( p2 => p_vector_0_13_port, g2 => 
                           g_vector_0_13_port, p1 => p_vector_0_12_port, g1 => 
                           g_vector_0_12_port, PG_P => p_vector_1_13_port, PG_G
                           => g_vector_1_13_port);
   std_PG_1_11 : PG_BLOCK_163 port map( p2 => p_vector_0_11_port, g2 => 
                           g_vector_0_11_port, p1 => p_vector_0_10_port, g1 => 
                           g_vector_0_10_port, PG_P => p_vector_1_11_port, PG_G
                           => g_vector_1_11_port);
   std_PG_1_9 : PG_BLOCK_162 port map( p2 => p_vector_0_9_port, g2 => 
                           g_vector_0_9_port, p1 => p_vector_0_8_port, g1 => 
                           g_vector_0_8_port, PG_P => p_vector_1_9_port, PG_G 
                           => g_vector_1_9_port);
   std_PG_1_7 : PG_BLOCK_161 port map( p2 => p_vector_0_7_port, g2 => 
                           g_vector_0_7_port, p1 => p_vector_0_6_port, g1 => 
                           g_vector_0_6_port, PG_P => p_vector_1_7_port, PG_G 
                           => g_vector_1_7_port);
   std_PG_1_5 : PG_BLOCK_160 port map( p2 => p_vector_0_5_port, g2 => 
                           g_vector_0_5_port, p1 => p_vector_0_4_port, g1 => 
                           g_vector_0_4_port, PG_P => p_vector_1_5_port, PG_G 
                           => g_vector_1_5_port);
   std_PG_1_3 : PG_BLOCK_159 port map( p2 => p_vector_0_3_port, g2 => 
                           g_vector_0_3_port, p1 => p_vector_0_2_port, g1 => 
                           g_vector_0_2_port, PG_P => p_vector_1_3_port, PG_G 
                           => g_vector_1_3_port);
   std_G_1_1 : G_BLOCK_51 port map( p2 => p_vector_0_1_port, g2 => 
                           g_vector_0_1_port, g1 => g_vector_0_0_port, G => 
                           g_vector_1_1_port);
   std_PG_2_63 : PG_BLOCK_158 port map( p2 => p_vector_1_63_port, g2 => 
                           g_vector_1_63_port, p1 => p_vector_1_61_port, g1 => 
                           g_vector_1_61_port, PG_P => p_vector_2_63_port, PG_G
                           => g_vector_2_63_port);
   std_PG_2_59 : PG_BLOCK_157 port map( p2 => p_vector_1_59_port, g2 => 
                           g_vector_1_59_port, p1 => p_vector_1_57_port, g1 => 
                           g_vector_1_57_port, PG_P => p_vector_2_59_port, PG_G
                           => g_vector_2_59_port);
   std_PG_2_55 : PG_BLOCK_156 port map( p2 => p_vector_1_55_port, g2 => 
                           g_vector_1_55_port, p1 => p_vector_1_53_port, g1 => 
                           g_vector_1_53_port, PG_P => p_vector_2_55_port, PG_G
                           => g_vector_2_55_port);
   std_PG_2_51 : PG_BLOCK_155 port map( p2 => p_vector_1_51_port, g2 => 
                           g_vector_1_51_port, p1 => p_vector_1_49_port, g1 => 
                           g_vector_1_49_port, PG_P => p_vector_2_51_port, PG_G
                           => g_vector_2_51_port);
   std_PG_2_47 : PG_BLOCK_154 port map( p2 => p_vector_1_47_port, g2 => 
                           g_vector_1_47_port, p1 => p_vector_1_45_port, g1 => 
                           g_vector_1_45_port, PG_P => p_vector_2_47_port, PG_G
                           => g_vector_2_47_port);
   std_PG_2_43 : PG_BLOCK_153 port map( p2 => p_vector_1_43_port, g2 => 
                           g_vector_1_43_port, p1 => p_vector_1_41_port, g1 => 
                           g_vector_1_41_port, PG_P => p_vector_2_43_port, PG_G
                           => g_vector_2_43_port);
   std_PG_2_39 : PG_BLOCK_152 port map( p2 => p_vector_1_39_port, g2 => 
                           g_vector_1_39_port, p1 => p_vector_1_37_port, g1 => 
                           g_vector_1_37_port, PG_P => p_vector_2_39_port, PG_G
                           => g_vector_2_39_port);
   std_PG_2_35 : PG_BLOCK_151 port map( p2 => p_vector_1_35_port, g2 => 
                           g_vector_1_35_port, p1 => p_vector_1_33_port, g1 => 
                           g_vector_1_33_port, PG_P => p_vector_2_35_port, PG_G
                           => g_vector_2_35_port);
   std_PG_2_31 : PG_BLOCK_150 port map( p2 => p_vector_1_31_port, g2 => 
                           g_vector_1_31_port, p1 => p_vector_1_29_port, g1 => 
                           g_vector_1_29_port, PG_P => p_vector_2_31_port, PG_G
                           => g_vector_2_31_port);
   std_PG_2_27 : PG_BLOCK_149 port map( p2 => p_vector_1_27_port, g2 => 
                           g_vector_1_27_port, p1 => p_vector_1_25_port, g1 => 
                           g_vector_1_25_port, PG_P => p_vector_2_27_port, PG_G
                           => g_vector_2_27_port);
   std_PG_2_23 : PG_BLOCK_148 port map( p2 => p_vector_1_23_port, g2 => 
                           g_vector_1_23_port, p1 => p_vector_1_21_port, g1 => 
                           g_vector_1_21_port, PG_P => p_vector_2_23_port, PG_G
                           => g_vector_2_23_port);
   std_PG_2_19 : PG_BLOCK_147 port map( p2 => p_vector_1_19_port, g2 => 
                           g_vector_1_19_port, p1 => p_vector_1_17_port, g1 => 
                           g_vector_1_17_port, PG_P => p_vector_2_19_port, PG_G
                           => g_vector_2_19_port);
   std_PG_2_15 : PG_BLOCK_146 port map( p2 => p_vector_1_15_port, g2 => 
                           g_vector_1_15_port, p1 => p_vector_1_13_port, g1 => 
                           g_vector_1_13_port, PG_P => p_vector_2_15_port, PG_G
                           => g_vector_2_15_port);
   std_PG_2_11 : PG_BLOCK_145 port map( p2 => p_vector_1_11_port, g2 => 
                           g_vector_1_11_port, p1 => p_vector_1_9_port, g1 => 
                           g_vector_1_9_port, PG_P => p_vector_2_11_port, PG_G 
                           => g_vector_2_11_port);
   std_PG_2_7 : PG_BLOCK_144 port map( p2 => p_vector_1_7_port, g2 => 
                           g_vector_1_7_port, p1 => p_vector_1_5_port, g1 => 
                           g_vector_1_5_port, PG_P => p_vector_2_7_port, PG_G 
                           => g_vector_2_7_port);
   std_G_2_3 : G_BLOCK_50 port map( p2 => p_vector_1_3_port, g2 => 
                           g_vector_1_3_port, g1 => g_vector_1_1_port, G => 
                           Co_0_port);
   std_PG_3_63 : PG_BLOCK_143 port map( p2 => p_vector_2_63_port, g2 => 
                           g_vector_2_63_port, p1 => p_vector_2_59_port, g1 => 
                           g_vector_2_59_port, PG_P => p_vector_3_63_port, PG_G
                           => g_vector_3_63_port);
   std_PG_3_55 : PG_BLOCK_142 port map( p2 => p_vector_2_55_port, g2 => 
                           g_vector_2_55_port, p1 => p_vector_2_51_port, g1 => 
                           g_vector_2_51_port, PG_P => p_vector_3_55_port, PG_G
                           => g_vector_3_55_port);
   std_PG_3_47 : PG_BLOCK_141 port map( p2 => p_vector_2_47_port, g2 => 
                           g_vector_2_47_port, p1 => p_vector_2_43_port, g1 => 
                           g_vector_2_43_port, PG_P => p_vector_3_47_port, PG_G
                           => g_vector_3_47_port);
   std_PG_3_39 : PG_BLOCK_140 port map( p2 => p_vector_2_39_port, g2 => 
                           g_vector_2_39_port, p1 => p_vector_2_35_port, g1 => 
                           g_vector_2_35_port, PG_P => p_vector_3_39_port, PG_G
                           => g_vector_3_39_port);
   std_PG_3_31 : PG_BLOCK_139 port map( p2 => p_vector_2_31_port, g2 => 
                           g_vector_2_31_port, p1 => p_vector_2_27_port, g1 => 
                           g_vector_2_27_port, PG_P => p_vector_3_31_port, PG_G
                           => g_vector_3_31_port);
   std_PG_3_23 : PG_BLOCK_138 port map( p2 => p_vector_2_23_port, g2 => 
                           g_vector_2_23_port, p1 => p_vector_2_19_port, g1 => 
                           g_vector_2_19_port, PG_P => p_vector_3_23_port, PG_G
                           => g_vector_3_23_port);
   std_PG_3_15 : PG_BLOCK_137 port map( p2 => p_vector_2_15_port, g2 => 
                           g_vector_2_15_port, p1 => p_vector_2_11_port, g1 => 
                           g_vector_2_11_port, PG_P => p_vector_3_15_port, PG_G
                           => g_vector_3_15_port);
   std_G_3_7 : G_BLOCK_49 port map( p2 => p_vector_2_7_port, g2 => 
                           g_vector_2_7_port, g1 => Co_0_port, G => Co_1_port);
   std_PG_4_63 : PG_BLOCK_136 port map( p2 => p_vector_3_63_port, g2 => 
                           g_vector_3_63_port, p1 => p_vector_3_55_port, g1 => 
                           g_vector_3_55_port, PG_P => p_vector_4_63_port, PG_G
                           => g_vector_4_63_port);
   add_PG_4_63_1 : PG_BLOCK_135 port map( p2 => p_vector_2_59_port, g2 => 
                           g_vector_2_59_port, p1 => p_vector_3_55_port, g1 => 
                           g_vector_3_55_port, PG_P => p_vector_4_59_port, PG_G
                           => g_vector_4_59_port);
   std_PG_4_47 : PG_BLOCK_134 port map( p2 => p_vector_3_47_port, g2 => 
                           g_vector_3_47_port, p1 => p_vector_3_39_port, g1 => 
                           g_vector_3_39_port, PG_P => p_vector_4_47_port, PG_G
                           => g_vector_4_47_port);
   add_PG_4_47_1 : PG_BLOCK_133 port map( p2 => p_vector_2_43_port, g2 => 
                           g_vector_2_43_port, p1 => p_vector_3_39_port, g1 => 
                           g_vector_3_39_port, PG_P => p_vector_4_43_port, PG_G
                           => g_vector_4_43_port);
   std_PG_4_31 : PG_BLOCK_132 port map( p2 => p_vector_3_31_port, g2 => 
                           g_vector_3_31_port, p1 => p_vector_3_23_port, g1 => 
                           g_vector_3_23_port, PG_P => p_vector_4_31_port, PG_G
                           => g_vector_4_31_port);
   add_PG_4_31_1 : PG_BLOCK_131 port map( p2 => p_vector_2_27_port, g2 => 
                           g_vector_2_27_port, p1 => p_vector_3_23_port, g1 => 
                           g_vector_3_23_port, PG_P => p_vector_4_27_port, PG_G
                           => g_vector_4_27_port);
   std_G_4_15 : G_BLOCK_48 port map( p2 => p_vector_3_15_port, g2 => 
                           g_vector_3_15_port, g1 => Co_1_port, G => Co_3_port)
                           ;
   add_G_4_15_1 : G_BLOCK_47 port map( p2 => p_vector_2_11_port, g2 => 
                           g_vector_2_11_port, g1 => Co_1_port, G => Co_2_port)
                           ;
   std_PG_5_63 : PG_BLOCK_130 port map( p2 => p_vector_4_63_port, g2 => 
                           g_vector_4_63_port, p1 => p_vector_4_47_port, g1 => 
                           g_vector_4_47_port, PG_P => p_vector_5_63_port, PG_G
                           => g_vector_5_63_port);
   add_PG_5_63_1 : PG_BLOCK_129 port map( p2 => p_vector_4_59_port, g2 => 
                           g_vector_4_59_port, p1 => p_vector_4_47_port, g1 => 
                           g_vector_4_47_port, PG_P => p_vector_5_59_port, PG_G
                           => g_vector_5_59_port);
   add_PG_5_63_2 : PG_BLOCK_128 port map( p2 => p_vector_3_55_port, g2 => 
                           g_vector_3_55_port, p1 => p_vector_4_47_port, g1 => 
                           g_vector_4_47_port, PG_P => p_vector_5_55_port, PG_G
                           => g_vector_5_55_port);
   add_PG_5_63_3 : PG_BLOCK_127 port map( p2 => p_vector_2_51_port, g2 => 
                           g_vector_2_51_port, p1 => p_vector_4_47_port, g1 => 
                           g_vector_4_47_port, PG_P => p_vector_5_51_port, PG_G
                           => g_vector_5_51_port);
   std_G_5_31 : G_BLOCK_46 port map( p2 => p_vector_4_31_port, g2 => 
                           g_vector_4_31_port, g1 => Co_3_port, G => Co_7_port)
                           ;
   add_G_5_31_1 : G_BLOCK_45 port map( p2 => p_vector_4_27_port, g2 => 
                           g_vector_4_27_port, g1 => Co_3_port, G => Co_6_port)
                           ;
   add_G_5_31_2 : G_BLOCK_44 port map( p2 => p_vector_3_23_port, g2 => 
                           g_vector_3_23_port, g1 => Co_3_port, G => Co_5_port)
                           ;
   add_G_5_31_3 : G_BLOCK_43 port map( p2 => p_vector_2_19_port, g2 => 
                           g_vector_2_19_port, g1 => Co_3_port, G => Co_4_port)
                           ;
   std_G_6_63 : G_BLOCK_42 port map( p2 => p_vector_5_63_port, g2 => 
                           g_vector_5_63_port, g1 => Co_7_port, G => Co_15_port
                           );
   add_G_6_63_1 : G_BLOCK_41 port map( p2 => p_vector_5_59_port, g2 => 
                           g_vector_5_59_port, g1 => Co_7_port, G => Co_14_port
                           );
   add_G_6_63_2 : G_BLOCK_40 port map( p2 => p_vector_5_55_port, g2 => 
                           g_vector_5_55_port, g1 => Co_7_port, G => Co_13_port
                           );
   add_G_6_63_3 : G_BLOCK_39 port map( p2 => p_vector_5_51_port, g2 => 
                           g_vector_5_51_port, g1 => Co_7_port, G => Co_12_port
                           );
   add_G_6_63_4 : G_BLOCK_38 port map( p2 => p_vector_4_47_port, g2 => 
                           g_vector_4_47_port, g1 => Co_7_port, G => Co_11_port
                           );
   add_G_6_63_5 : G_BLOCK_37 port map( p2 => p_vector_4_43_port, g2 => 
                           g_vector_4_43_port, g1 => Co_7_port, G => Co_10_port
                           );
   add_G_6_63_6 : G_BLOCK_36 port map( p2 => p_vector_3_39_port, g2 => 
                           g_vector_3_39_port, g1 => Co_7_port, G => Co_9_port)
                           ;
   add_G_6_63_7 : G_BLOCK_35 port map( p2 => p_vector_2_35_port, g2 => 
                           g_vector_2_35_port, g1 => Co_7_port, G => Co_8_port)
                           ;
   U1 : OAI21_X1 port map( B1 => n2, B2 => n1, A => n3, ZN => g_vector_0_0_port
                           );
   U2 : OAI21_X1 port map( B1 => A(0), B2 => B(0), A => Cin, ZN => n3);
   U3 : INV_X1 port map( A => A(0), ZN => n2);
   U4 : INV_X1 port map( A => B(0), ZN => n1);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand41_0 is

   port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);

end nand41_0;

architecture SYN_behavioral of nand41_0 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND4_X1 port map( A1 => in4, A2 => in3, A3 => in2, A4 => in1, ZN => o)
                           ;

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nand31_0 is

   port( in1, in2, in3 : in std_logic;  o : out std_logic);

end nand31_0;

architecture SYN_behavioral of nand31_0 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND3_X1 port map( A1 => in2, A2 => in1, A3 => in3, ZN => o);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX81_GENERIC_NBIT32 is

   port( A, B, C, D, E, F, G, H : in std_logic_vector (31 downto 0);  SEL : in 
         std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end MUX81_GENERIC_NBIT32;

architecture SYN_structural of MUX81_GENERIC_NBIT32 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX81_1
      port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
            downto 0);  Y : out std_logic);
   end component;
   
   component MUX81_2
      port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
            downto 0);  Y : out std_logic);
   end component;
   
   component MUX81_3
      port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
            downto 0);  Y : out std_logic);
   end component;
   
   component MUX81_4
      port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
            downto 0);  Y : out std_logic);
   end component;
   
   component MUX81_5
      port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
            downto 0);  Y : out std_logic);
   end component;
   
   component MUX81_6
      port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
            downto 0);  Y : out std_logic);
   end component;
   
   component MUX81_7
      port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
            downto 0);  Y : out std_logic);
   end component;
   
   component MUX81_8
      port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
            downto 0);  Y : out std_logic);
   end component;
   
   component MUX81_9
      port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
            downto 0);  Y : out std_logic);
   end component;
   
   component MUX81_10
      port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
            downto 0);  Y : out std_logic);
   end component;
   
   component MUX81_11
      port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
            downto 0);  Y : out std_logic);
   end component;
   
   component MUX81_12
      port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
            downto 0);  Y : out std_logic);
   end component;
   
   component MUX81_13
      port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
            downto 0);  Y : out std_logic);
   end component;
   
   component MUX81_14
      port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
            downto 0);  Y : out std_logic);
   end component;
   
   component MUX81_15
      port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
            downto 0);  Y : out std_logic);
   end component;
   
   component MUX81_16
      port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
            downto 0);  Y : out std_logic);
   end component;
   
   component MUX81_17
      port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
            downto 0);  Y : out std_logic);
   end component;
   
   component MUX81_18
      port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
            downto 0);  Y : out std_logic);
   end component;
   
   component MUX81_19
      port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
            downto 0);  Y : out std_logic);
   end component;
   
   component MUX81_20
      port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
            downto 0);  Y : out std_logic);
   end component;
   
   component MUX81_21
      port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
            downto 0);  Y : out std_logic);
   end component;
   
   component MUX81_22
      port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
            downto 0);  Y : out std_logic);
   end component;
   
   component MUX81_23
      port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
            downto 0);  Y : out std_logic);
   end component;
   
   component MUX81_24
      port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
            downto 0);  Y : out std_logic);
   end component;
   
   component MUX81_25
      port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
            downto 0);  Y : out std_logic);
   end component;
   
   component MUX81_26
      port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
            downto 0);  Y : out std_logic);
   end component;
   
   component MUX81_27
      port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
            downto 0);  Y : out std_logic);
   end component;
   
   component MUX81_28
      port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
            downto 0);  Y : out std_logic);
   end component;
   
   component MUX81_29
      port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
            downto 0);  Y : out std_logic);
   end component;
   
   component MUX81_30
      port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
            downto 0);  Y : out std_logic);
   end component;
   
   component MUX81_31
      port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
            downto 0);  Y : out std_logic);
   end component;
   
   component MUX81_0
      port( A, B, C, D, E, F, G, H : in std_logic;  S : in std_logic_vector (2 
            downto 0);  Y : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9 : std_logic;

begin
   
   MUXES_0 : MUX81_0 port map( A => A(0), B => B(0), C => C(0), D => D(0), E =>
                           E(0), F => F(0), G => G(0), H => H(0), S(2) => n9, 
                           S(1) => n6, S(0) => n3, Y => Y(0));
   MUXES_1 : MUX81_31 port map( A => A(1), B => B(1), C => C(1), D => D(1), E 
                           => E(1), F => F(1), G => G(1), H => H(1), S(2) => n7
                           , S(1) => n4, S(0) => n1, Y => Y(1));
   MUXES_2 : MUX81_30 port map( A => A(2), B => B(2), C => C(2), D => D(2), E 
                           => E(2), F => F(2), G => G(2), H => H(2), S(2) => n7
                           , S(1) => n4, S(0) => n1, Y => Y(2));
   MUXES_3 : MUX81_29 port map( A => A(3), B => B(3), C => C(3), D => D(3), E 
                           => E(3), F => F(3), G => G(3), H => H(3), S(2) => n7
                           , S(1) => n4, S(0) => n1, Y => Y(3));
   MUXES_4 : MUX81_28 port map( A => A(4), B => B(4), C => C(4), D => D(4), E 
                           => E(4), F => F(4), G => G(4), H => H(4), S(2) => n7
                           , S(1) => n4, S(0) => n1, Y => Y(4));
   MUXES_5 : MUX81_27 port map( A => A(5), B => B(5), C => C(5), D => D(5), E 
                           => E(5), F => F(5), G => G(5), H => H(5), S(2) => n7
                           , S(1) => n4, S(0) => n1, Y => Y(5));
   MUXES_6 : MUX81_26 port map( A => A(6), B => B(6), C => C(6), D => D(6), E 
                           => E(6), F => F(6), G => G(6), H => H(6), S(2) => n7
                           , S(1) => n4, S(0) => n1, Y => Y(6));
   MUXES_7 : MUX81_25 port map( A => A(7), B => B(7), C => C(7), D => D(7), E 
                           => E(7), F => F(7), G => G(7), H => H(7), S(2) => n7
                           , S(1) => n4, S(0) => n1, Y => Y(7));
   MUXES_8 : MUX81_24 port map( A => A(8), B => B(8), C => C(8), D => D(8), E 
                           => E(8), F => F(8), G => G(8), H => H(8), S(2) => n7
                           , S(1) => n4, S(0) => n1, Y => Y(8));
   MUXES_9 : MUX81_23 port map( A => A(9), B => B(9), C => C(9), D => D(9), E 
                           => E(9), F => F(9), G => G(9), H => H(9), S(2) => n7
                           , S(1) => n4, S(0) => n1, Y => Y(9));
   MUXES_10 : MUX81_22 port map( A => A(10), B => B(10), C => C(10), D => D(10)
                           , E => E(10), F => F(10), G => G(10), H => H(10), 
                           S(2) => n7, S(1) => n4, S(0) => n1, Y => Y(10));
   MUXES_11 : MUX81_21 port map( A => A(11), B => B(11), C => C(11), D => D(11)
                           , E => E(11), F => F(11), G => G(11), H => H(11), 
                           S(2) => n7, S(1) => n4, S(0) => n1, Y => Y(11));
   MUXES_12 : MUX81_20 port map( A => A(12), B => B(12), C => C(12), D => D(12)
                           , E => E(12), F => F(12), G => G(12), H => H(12), 
                           S(2) => n8, S(1) => n4, S(0) => n1, Y => Y(12));
   MUXES_13 : MUX81_19 port map( A => A(13), B => B(13), C => C(13), D => D(13)
                           , E => E(13), F => F(13), G => G(13), H => H(13), 
                           S(2) => n8, S(1) => n5, S(0) => n2, Y => Y(13));
   MUXES_14 : MUX81_18 port map( A => A(14), B => B(14), C => C(14), D => D(14)
                           , E => E(14), F => F(14), G => G(14), H => H(14), 
                           S(2) => n8, S(1) => n5, S(0) => n2, Y => Y(14));
   MUXES_15 : MUX81_17 port map( A => A(15), B => B(15), C => C(15), D => D(15)
                           , E => E(15), F => F(15), G => G(15), H => H(15), 
                           S(2) => n8, S(1) => n5, S(0) => n2, Y => Y(15));
   MUXES_16 : MUX81_16 port map( A => A(16), B => B(16), C => C(16), D => D(16)
                           , E => E(16), F => F(16), G => G(16), H => H(16), 
                           S(2) => n8, S(1) => n5, S(0) => n2, Y => Y(16));
   MUXES_17 : MUX81_15 port map( A => A(17), B => B(17), C => C(17), D => D(17)
                           , E => E(17), F => F(17), G => G(17), H => H(17), 
                           S(2) => n8, S(1) => n5, S(0) => n2, Y => Y(17));
   MUXES_18 : MUX81_14 port map( A => A(18), B => B(18), C => C(18), D => D(18)
                           , E => E(18), F => F(18), G => G(18), H => H(18), 
                           S(2) => n8, S(1) => n5, S(0) => n2, Y => Y(18));
   MUXES_19 : MUX81_13 port map( A => A(19), B => B(19), C => C(19), D => D(19)
                           , E => E(19), F => F(19), G => G(19), H => H(19), 
                           S(2) => n8, S(1) => n5, S(0) => n2, Y => Y(19));
   MUXES_20 : MUX81_12 port map( A => A(20), B => B(20), C => C(20), D => D(20)
                           , E => E(20), F => F(20), G => G(20), H => H(20), 
                           S(2) => n8, S(1) => n5, S(0) => n2, Y => Y(20));
   MUXES_21 : MUX81_11 port map( A => A(21), B => B(21), C => C(21), D => D(21)
                           , E => E(21), F => F(21), G => G(21), H => H(21), 
                           S(2) => n8, S(1) => n5, S(0) => n2, Y => Y(21));
   MUXES_22 : MUX81_10 port map( A => A(22), B => B(22), C => C(22), D => D(22)
                           , E => E(22), F => F(22), G => G(22), H => H(22), 
                           S(2) => n8, S(1) => n5, S(0) => n2, Y => Y(22));
   MUXES_23 : MUX81_9 port map( A => A(23), B => B(23), C => C(23), D => D(23),
                           E => E(23), F => F(23), G => G(23), H => H(23), S(2)
                           => n9, S(1) => n5, S(0) => n2, Y => Y(23));
   MUXES_24 : MUX81_8 port map( A => A(24), B => B(24), C => C(24), D => D(24),
                           E => E(24), F => F(24), G => G(24), H => H(24), S(2)
                           => n9, S(1) => n5, S(0) => n2, Y => Y(24));
   MUXES_25 : MUX81_7 port map( A => A(25), B => B(25), C => C(25), D => D(25),
                           E => E(25), F => F(25), G => G(25), H => H(25), S(2)
                           => n9, S(1) => n6, S(0) => n3, Y => Y(25));
   MUXES_26 : MUX81_6 port map( A => A(26), B => B(26), C => C(26), D => D(26),
                           E => E(26), F => F(26), G => G(26), H => H(26), S(2)
                           => n9, S(1) => n6, S(0) => n3, Y => Y(26));
   MUXES_27 : MUX81_5 port map( A => A(27), B => B(27), C => C(27), D => D(27),
                           E => E(27), F => F(27), G => G(27), H => H(27), S(2)
                           => n9, S(1) => n6, S(0) => n3, Y => Y(27));
   MUXES_28 : MUX81_4 port map( A => A(28), B => B(28), C => C(28), D => D(28),
                           E => E(28), F => F(28), G => G(28), H => H(28), S(2)
                           => n9, S(1) => n6, S(0) => n3, Y => Y(28));
   MUXES_29 : MUX81_3 port map( A => A(29), B => B(29), C => C(29), D => D(29),
                           E => E(29), F => F(29), G => G(29), H => H(29), S(2)
                           => n9, S(1) => n6, S(0) => n3, Y => Y(29));
   MUXES_30 : MUX81_2 port map( A => A(30), B => B(30), C => C(30), D => D(30),
                           E => E(30), F => F(30), G => G(30), H => H(30), S(2)
                           => n9, S(1) => n6, S(0) => n3, Y => Y(30));
   MUXES_31 : MUX81_1 port map( A => A(31), B => B(31), C => C(31), D => D(31),
                           E => E(31), F => F(31), G => G(31), H => H(31), S(2)
                           => n9, S(1) => n6, S(0) => n3, Y => Y(31));
   U1 : BUF_X2 port map( A => SEL(0), Z => n2);
   U2 : BUF_X2 port map( A => SEL(0), Z => n1);
   U3 : BUF_X1 port map( A => SEL(1), Z => n6);
   U4 : BUF_X2 port map( A => SEL(0), Z => n3);
   U5 : BUF_X2 port map( A => SEL(1), Z => n5);
   U6 : BUF_X2 port map( A => SEL(1), Z => n4);
   U7 : BUF_X1 port map( A => SEL(2), Z => n8);
   U8 : BUF_X1 port map( A => SEL(2), Z => n7);
   U9 : BUF_X1 port map( A => SEL(2), Z => n9);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity mask_shifter_NBITS40 is

   port( R1 : in std_logic_vector (39 downto 0);  LnR : in std_logic;  mask_sh0
         , mask_sh1, mask_sh2, mask_sh3, mask_sh4, mask_sh5, mask_sh6, mask_sh7
         : out std_logic_vector (31 downto 0));

end mask_shifter_NBITS40;

architecture SYN_structural of mask_shifter_NBITS40 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, 
      n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36
      , n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, 
      n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65
      , n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n1, n2, n3,
      n4, n5, n6, n7, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95 : std_logic;

begin
   mask_sh4 <= ( R1(35), R1(34), R1(33), R1(32), R1(31), R1(30), R1(29), R1(28)
      , R1(27), R1(26), R1(25), R1(24), R1(23), R1(22), R1(21), R1(20), R1(19),
      R1(18), R1(17), R1(16), R1(15), R1(14), R1(13), R1(12), R1(11), R1(10), 
      R1(9), R1(8), R1(7), R1(6), R1(5), R1(4) );
   
   U1 : NAND2_X1 port map( A1 => n58, A2 => n62, ZN => mask_sh6(13));
   U2 : NAND2_X1 port map( A1 => n60, A2 => n64, ZN => mask_sh6(12));
   U3 : NAND2_X1 port map( A1 => n61, A2 => n66, ZN => mask_sh6(11));
   U4 : NAND2_X1 port map( A1 => n50, A2 => n53, ZN => mask_sh6(17));
   U5 : NAND2_X1 port map( A1 => n30, A2 => n51, ZN => mask_sh2(22));
   U6 : NAND2_X1 port map( A1 => n32, A2 => n53, ZN => mask_sh2(21));
   U7 : NAND2_X1 port map( A1 => n52, A2 => n55, ZN => mask_sh6(16));
   U8 : NAND2_X1 port map( A1 => n54, A2 => n57, ZN => mask_sh6(15));
   U9 : NAND2_X1 port map( A1 => n56, A2 => n59, ZN => mask_sh6(14));
   U10 : NAND2_X1 port map( A1 => n34, A2 => n55, ZN => mask_sh2(20));
   U11 : NAND2_X1 port map( A1 => n37, A2 => n57, ZN => mask_sh2(19));
   U12 : NAND2_X1 port map( A1 => n39, A2 => n59, ZN => mask_sh2(18));
   U13 : NAND2_X1 port map( A1 => n34, A2 => n51, ZN => mask_sh3(21));
   U14 : NAND2_X1 port map( A1 => n37, A2 => n53, ZN => mask_sh3(20));
   U15 : NAND2_X1 port map( A1 => n39, A2 => n55, ZN => mask_sh3(19));
   U16 : NAND2_X1 port map( A1 => n26, A2 => n47, ZN => mask_sh2(24));
   U17 : NAND2_X1 port map( A1 => n28, A2 => n49, ZN => mask_sh2(23));
   U18 : NAND2_X1 port map( A1 => n30, A2 => n47, ZN => mask_sh3(23));
   U19 : NAND2_X1 port map( A1 => n32, A2 => n49, ZN => mask_sh3(22));
   U20 : NAND2_X1 port map( A1 => n22, A2 => n42, ZN => mask_sh2(26));
   U21 : NAND2_X1 port map( A1 => n23, A2 => n44, ZN => mask_sh2(25));
   U22 : NAND2_X1 port map( A1 => n34, A2 => n38, ZN => mask_sh6(24));
   U23 : NAND2_X1 port map( A1 => n26, A2 => n42, ZN => mask_sh3(25));
   U24 : NAND2_X1 port map( A1 => n28, A2 => n44, ZN => mask_sh3(24));
   U25 : NAND2_X1 port map( A1 => n37, A2 => n40, ZN => mask_sh6(23));
   U26 : NAND2_X1 port map( A1 => n22, A2 => n38, ZN => mask_sh3(27));
   U27 : NAND2_X1 port map( A1 => n23, A2 => n40, ZN => mask_sh3(26));
   U28 : NAND2_X1 port map( A1 => n8, A2 => n13, ZN => mask_sh6(8));
   U29 : NAND2_X1 port map( A1 => n10, A2 => n14, ZN => mask_sh6(7));
   U30 : NAND2_X1 port map( A1 => n8, A2 => n46, ZN => mask_sh3(5));
   U31 : NAND2_X1 port map( A1 => n11, A2 => n54, ZN => mask_sh3(12));
   U32 : NAND2_X1 port map( A1 => n16, A2 => n60, ZN => mask_sh3(9));
   U33 : NAND2_X1 port map( A1 => n14, A2 => n58, ZN => mask_sh3(10));
   U34 : NAND2_X1 port map( A1 => n20, A2 => n63, ZN => mask_sh3(7));
   U35 : NAND2_X1 port map( A1 => n18, A2 => n61, ZN => mask_sh3(8));
   U36 : NAND2_X1 port map( A1 => n24, A2 => n65, ZN => mask_sh3(6));
   U37 : NAND2_X1 port map( A1 => n13, A2 => n56, ZN => mask_sh3(11));
   U38 : NAND2_X1 port map( A1 => n38, A2 => n70, ZN => mask_sh2(28));
   U39 : NAND2_X1 port map( A1 => n40, A2 => n68, ZN => mask_sh2(27));
   U40 : NAND2_X1 port map( A1 => n36, A2 => n73, ZN => mask_sh2(29));
   U41 : NAND2_X1 port map( A1 => n36, A2 => n68, ZN => mask_sh3(28));
   U42 : NAND2_X1 port map( A1 => n30, A2 => n35, ZN => mask_sh6(26));
   U43 : NAND2_X1 port map( A1 => n22, A2 => n27, ZN => mask_sh6(30));
   U44 : NAND2_X1 port map( A1 => n23, A2 => n29, ZN => mask_sh6(29));
   U45 : NAND2_X1 port map( A1 => n26, A2 => n31, ZN => mask_sh6(28));
   U46 : NAND2_X1 port map( A1 => n28, A2 => n33, ZN => mask_sh6(27));
   U47 : NAND2_X1 port map( A1 => n54, A2 => n62, ZN => mask_sh5(14));
   U48 : NAND2_X1 port map( A1 => n56, A2 => n64, ZN => mask_sh5(13));
   U49 : NAND2_X1 port map( A1 => n58, A2 => n66, ZN => mask_sh5(12));
   U50 : NAND2_X1 port map( A1 => n65, A2 => n66, ZN => mask_sh7(10));
   U51 : NAND2_X1 port map( A1 => n43, A2 => n51, ZN => mask_sh5(19));
   U52 : NAND2_X1 port map( A1 => n45, A2 => n53, ZN => mask_sh5(18));
   U53 : NAND2_X1 port map( A1 => n48, A2 => n55, ZN => mask_sh5(17));
   U54 : NAND2_X1 port map( A1 => n50, A2 => n57, ZN => mask_sh5(16));
   U55 : NAND2_X1 port map( A1 => n52, A2 => n59, ZN => mask_sh5(15));
   U56 : NAND2_X1 port map( A1 => n39, A2 => n47, ZN => mask_sh5(21));
   U57 : NAND2_X1 port map( A1 => n41, A2 => n49, ZN => mask_sh5(20));
   U58 : NAND2_X1 port map( A1 => n34, A2 => n42, ZN => mask_sh5(23));
   U59 : NAND2_X1 port map( A1 => n37, A2 => n44, ZN => mask_sh5(22));
   U60 : NAND2_X1 port map( A1 => n30, A2 => n38, ZN => mask_sh5(25));
   U61 : NAND2_X1 port map( A1 => n32, A2 => n40, ZN => mask_sh5(24));
   U62 : NAND2_X1 port map( A1 => n8, A2 => n16, ZN => mask_sh5(7));
   U63 : NAND2_X1 port map( A1 => n12, A2 => n20, ZN => mask_sh5(5));
   U64 : NAND2_X1 port map( A1 => n8, A2 => n9, ZN => mask_sh7(9));
   U65 : NAND2_X1 port map( A1 => n10, A2 => n18, ZN => mask_sh5(6));
   U66 : NAND2_X1 port map( A1 => n9, A2 => n60, ZN => mask_sh5(11));
   U67 : NAND2_X1 port map( A1 => n47, A2 => n48, ZN => mask_sh7(19));
   U68 : NAND2_X1 port map( A1 => n49, A2 => n50, ZN => mask_sh7(18));
   U69 : NAND2_X1 port map( A1 => n13, A2 => n63, ZN => mask_sh5(9));
   U70 : NAND2_X1 port map( A1 => n42, A2 => n43, ZN => mask_sh7(21));
   U71 : NAND2_X1 port map( A1 => n44, A2 => n45, ZN => mask_sh7(20));
   U72 : NAND2_X1 port map( A1 => n11, A2 => n61, ZN => mask_sh5(10));
   U73 : NAND2_X1 port map( A1 => n14, A2 => n65, ZN => mask_sh5(8));
   U74 : NAND2_X1 port map( A1 => n40, A2 => n41, ZN => mask_sh7(22));
   U75 : NAND2_X1 port map( A1 => n26, A2 => n35, ZN => mask_sh5(27));
   U76 : NAND2_X1 port map( A1 => n34, A2 => n35, ZN => mask_sh7(25));
   U77 : NAND2_X1 port map( A1 => n22, A2 => n31, ZN => mask_sh5(29));
   U78 : NAND2_X1 port map( A1 => n23, A2 => n33, ZN => mask_sh5(28));
   U79 : NAND2_X1 port map( A1 => n32, A2 => n33, ZN => mask_sh7(26));
   U80 : NAND2_X1 port map( A1 => n68, A2 => n29, ZN => mask_sh5(30));
   U81 : NAND2_X1 port map( A1 => n70, A2 => n27, ZN => mask_sh5(31));
   U82 : NAND2_X1 port map( A1 => n41, A2 => n62, ZN => mask_sh2(17));
   U83 : NAND2_X1 port map( A1 => n43, A2 => n64, ZN => mask_sh2(16));
   U84 : NAND2_X1 port map( A1 => n45, A2 => n66, ZN => mask_sh2(15));
   U85 : NAND2_X1 port map( A1 => n45, A2 => n62, ZN => mask_sh3(16));
   U86 : NAND2_X1 port map( A1 => n48, A2 => n64, ZN => mask_sh3(15));
   U87 : NAND2_X1 port map( A1 => n50, A2 => n66, ZN => mask_sh3(14));
   U88 : NAND2_X1 port map( A1 => n41, A2 => n57, ZN => mask_sh3(18));
   U89 : NAND2_X1 port map( A1 => n43, A2 => n59, ZN => mask_sh3(17));
   U90 : NAND2_X1 port map( A1 => n13, A2 => n52, ZN => mask_sh2(12));
   U91 : NAND2_X1 port map( A1 => n14, A2 => n54, ZN => mask_sh2(11));
   U92 : NAND2_X1 port map( A1 => n20, A2 => n60, ZN => mask_sh2(8));
   U93 : NAND2_X1 port map( A1 => n9, A2 => n48, ZN => mask_sh2(14));
   U94 : NAND2_X1 port map( A1 => n11, A2 => n50, ZN => mask_sh2(13));
   U95 : NAND2_X1 port map( A1 => n18, A2 => n58, ZN => mask_sh2(9));
   U96 : NAND2_X1 port map( A1 => n46, A2 => n63, ZN => mask_sh2(6));
   U97 : NAND2_X1 port map( A1 => n9, A2 => n52, ZN => mask_sh3(13));
   U98 : NAND2_X1 port map( A1 => n24, A2 => n61, ZN => mask_sh2(7));
   U99 : NAND2_X1 port map( A1 => n16, A2 => n56, ZN => mask_sh2(10));
   U100 : NAND2_X1 port map( A1 => n35, A2 => n72, ZN => mask_sh2(30));
   U101 : NAND2_X1 port map( A1 => n35, A2 => n70, ZN => mask_sh3(29));
   U102 : NAND2_X1 port map( A1 => n33, A2 => n76, ZN => mask_sh2(31));
   U103 : NAND2_X1 port map( A1 => n33, A2 => n73, ZN => mask_sh3(30));
   U104 : NAND2_X1 port map( A1 => n31, A2 => n72, ZN => mask_sh3(31));
   U105 : NAND2_X1 port map( A1 => R1(19), A2 => n78, ZN => n62);
   U106 : NAND2_X1 port map( A1 => R1(18), A2 => n78, ZN => n64);
   U107 : NAND2_X1 port map( A1 => R1(17), A2 => n78, ZN => n66);
   U108 : NAND2_X1 port map( A1 => R1(24), A2 => n7, ZN => n51);
   U109 : NAND2_X1 port map( A1 => R1(23), A2 => n78, ZN => n53);
   U110 : NAND2_X1 port map( A1 => R1(22), A2 => n78, ZN => n55);
   U111 : NAND2_X1 port map( A1 => R1(21), A2 => n78, ZN => n57);
   U112 : NAND2_X1 port map( A1 => R1(20), A2 => n78, ZN => n59);
   U113 : NAND2_X1 port map( A1 => R1(26), A2 => n7, ZN => n47);
   U114 : NAND2_X1 port map( A1 => R1(25), A2 => n78, ZN => n49);
   U115 : NAND2_X1 port map( A1 => n89, A2 => R1(16), ZN => n56);
   U116 : NAND2_X1 port map( A1 => R1(18), A2 => n79, ZN => n52);
   U117 : NAND2_X1 port map( A1 => R1(17), A2 => n87, ZN => n54);
   U118 : NAND2_X1 port map( A1 => R1(14), A2 => n87, ZN => n60);
   U119 : NAND2_X1 port map( A1 => R1(28), A2 => n7, ZN => n42);
   U120 : NAND2_X1 port map( A1 => R1(27), A2 => n78, ZN => n44);
   U121 : NAND2_X1 port map( A1 => R1(30), A2 => n7, ZN => n38);
   U122 : NAND2_X1 port map( A1 => R1(20), A2 => n79, ZN => n48);
   U123 : NAND2_X1 port map( A1 => R1(19), A2 => n80, ZN => n50);
   U124 : NAND2_X1 port map( A1 => R1(15), A2 => n86, ZN => n58);
   U125 : NAND2_X1 port map( A1 => R1(12), A2 => n85, ZN => n63);
   U126 : NAND2_X1 port map( A1 => R1(29), A2 => n78, ZN => n40);
   U127 : NAND2_X1 port map( A1 => R1(31), A2 => n7, ZN => n36);
   U128 : NAND2_X1 port map( A1 => R1(22), A2 => n81, ZN => n43);
   U129 : NAND2_X1 port map( A1 => R1(21), A2 => n80, ZN => n45);
   U130 : NAND2_X1 port map( A1 => R1(13), A2 => n86, ZN => n61);
   U131 : NAND2_X1 port map( A1 => R1(11), A2 => n84, ZN => n65);
   U132 : NAND2_X1 port map( A1 => R1(14), A2 => n78, ZN => n13);
   U133 : NAND2_X1 port map( A1 => R1(12), A2 => n78, ZN => n16);
   U134 : NAND2_X1 port map( A1 => R1(8), A2 => n78, ZN => n46);
   U135 : NAND2_X1 port map( A1 => R1(24), A2 => n81, ZN => n39);
   U136 : NAND2_X1 port map( A1 => R1(23), A2 => n81, ZN => n41);
   U137 : NAND2_X1 port map( A1 => R1(10), A2 => n7, ZN => n20);
   U138 : NAND2_X1 port map( A1 => R1(16), A2 => n78, ZN => n9);
   U139 : NAND2_X1 port map( A1 => R1(15), A2 => n78, ZN => n11);
   U140 : NAND2_X1 port map( A1 => R1(13), A2 => n78, ZN => n14);
   U141 : NAND2_X1 port map( A1 => R1(11), A2 => n78, ZN => n18);
   U142 : NAND2_X1 port map( A1 => R1(9), A2 => n7, ZN => n24);
   U143 : NAND2_X1 port map( A1 => R1(25), A2 => n82, ZN => n37);
   U144 : NAND2_X1 port map( A1 => R1(32), A2 => n82, ZN => n22);
   U145 : NAND2_X1 port map( A1 => R1(31), A2 => n83, ZN => n23);
   U146 : NAND2_X1 port map( A1 => R1(9), A2 => n83, ZN => n10);
   U147 : NAND2_X1 port map( A1 => R1(8), A2 => n80, ZN => n12);
   U148 : NAND2_X1 port map( A1 => R1(30), A2 => n84, ZN => n26);
   U149 : NAND2_X1 port map( A1 => R1(29), A2 => n83, ZN => n28);
   U150 : NAND2_X1 port map( A1 => R1(28), A2 => n82, ZN => n30);
   U151 : NAND2_X1 port map( A1 => R1(27), A2 => n81, ZN => n32);
   U152 : NAND2_X1 port map( A1 => R1(26), A2 => n82, ZN => n34);
   U153 : NAND2_X1 port map( A1 => R1(10), A2 => n86, ZN => n8);
   U154 : NAND2_X1 port map( A1 => R1(32), A2 => n7, ZN => n35);
   U155 : NAND2_X1 port map( A1 => R1(33), A2 => n84, ZN => n68);
   U156 : NAND2_X1 port map( A1 => R1(33), A2 => n7, ZN => n33);
   U157 : NAND2_X1 port map( A1 => R1(34), A2 => n84, ZN => n70);
   U158 : NAND2_X1 port map( A1 => R1(34), A2 => n7, ZN => n31);
   U159 : NAND2_X1 port map( A1 => R1(36), A2 => n7, ZN => n27);
   U160 : NAND2_X1 port map( A1 => R1(35), A2 => n7, ZN => n29);
   U161 : OAI21_X1 port map( B1 => n88, B2 => n93, A => n68, ZN => mask_sh6(31)
                           );
   U162 : NAND2_X1 port map( A1 => n43, A2 => n47, ZN => mask_sh6(20));
   U163 : NAND2_X1 port map( A1 => n45, A2 => n49, ZN => mask_sh6(19));
   U164 : NAND2_X1 port map( A1 => n10, A2 => n67, ZN => mask_sh3(4));
   U165 : NAND2_X1 port map( A1 => n12, A2 => n16, ZN => mask_sh6(6));
   U166 : NAND2_X1 port map( A1 => n9, A2 => n63, ZN => mask_sh6(10));
   U167 : NAND2_X1 port map( A1 => n11, A2 => n65, ZN => mask_sh6(9));
   U168 : NAND2_X1 port map( A1 => n46, A2 => n21, ZN => mask_sh6(2));
   U169 : NAND2_X1 port map( A1 => n20, A2 => n17, ZN => mask_sh6(4));
   U170 : NAND2_X1 port map( A1 => n18, A2 => n15, ZN => mask_sh6(5));
   U171 : NAND2_X1 port map( A1 => n12, A2 => n69, ZN => mask_sh3(3));
   U172 : NAND2_X1 port map( A1 => n24, A2 => n19, ZN => mask_sh6(3));
   U173 : INV_X1 port map( A => R1(37), ZN => n93);
   U174 : NAND2_X1 port map( A1 => n39, A2 => n42, ZN => mask_sh6(22));
   U175 : NAND2_X1 port map( A1 => n41, A2 => n44, ZN => mask_sh6(21));
   U176 : NAND2_X1 port map( A1 => n48, A2 => n51, ZN => mask_sh6(18));
   U177 : NAND2_X1 port map( A1 => n32, A2 => n36, ZN => mask_sh6(25));
   U178 : NAND2_X1 port map( A1 => n46, A2 => n17, ZN => mask_sh5(3));
   U179 : NAND2_X1 port map( A1 => n14, A2 => n15, ZN => mask_sh7(6));
   U180 : NAND2_X1 port map( A1 => n24, A2 => n15, ZN => mask_sh5(4));
   U181 : NAND2_X1 port map( A1 => R1(36), A2 => n85, ZN => n72);
   U182 : NAND2_X1 port map( A1 => R1(35), A2 => n85, ZN => n73);
   U183 : OAI21_X1 port map( B1 => n95, B2 => n78, A => n36, ZN => mask_sh0(31)
                           );
   U184 : INV_X1 port map( A => R1(39), ZN => n95);
   U185 : OAI21_X1 port map( B1 => n78, B2 => n94, A => n38, ZN => mask_sh0(30)
                           );
   U186 : NAND2_X1 port map( A1 => n40, A2 => n76, ZN => mask_sh0(29));
   U187 : NAND2_X1 port map( A1 => n42, A2 => n72, ZN => mask_sh0(28));
   U188 : NAND2_X1 port map( A1 => n44, A2 => n73, ZN => mask_sh0(27));
   U189 : NAND2_X1 port map( A1 => n47, A2 => n70, ZN => mask_sh0(26));
   U190 : NAND2_X1 port map( A1 => n49, A2 => n68, ZN => mask_sh0(25));
   U191 : NAND2_X1 port map( A1 => n22, A2 => n51, ZN => mask_sh0(24));
   U192 : NAND2_X1 port map( A1 => n23, A2 => n53, ZN => mask_sh0(23));
   U193 : NAND2_X1 port map( A1 => n26, A2 => n55, ZN => mask_sh0(22));
   U194 : NAND2_X1 port map( A1 => n28, A2 => n57, ZN => mask_sh0(21));
   U195 : NAND2_X1 port map( A1 => n30, A2 => n59, ZN => mask_sh0(20));
   U196 : NAND2_X1 port map( A1 => n32, A2 => n62, ZN => mask_sh0(19));
   U197 : NAND2_X1 port map( A1 => n34, A2 => n64, ZN => mask_sh0(18));
   U198 : NAND2_X1 port map( A1 => n9, A2 => n39, ZN => mask_sh0(16));
   U199 : NAND2_X1 port map( A1 => n11, A2 => n41, ZN => mask_sh0(15));
   U200 : NAND2_X1 port map( A1 => n13, A2 => n43, ZN => mask_sh0(14));
   U201 : NAND2_X1 port map( A1 => n14, A2 => n45, ZN => mask_sh0(13));
   U202 : NAND2_X1 port map( A1 => n16, A2 => n48, ZN => mask_sh0(12));
   U203 : NAND2_X1 port map( A1 => n18, A2 => n50, ZN => mask_sh0(11));
   U204 : NAND2_X1 port map( A1 => n20, A2 => n52, ZN => mask_sh0(10));
   U205 : NAND2_X1 port map( A1 => n24, A2 => n54, ZN => mask_sh0(9));
   U206 : NAND2_X1 port map( A1 => n46, A2 => n56, ZN => mask_sh0(8));
   U207 : NAND2_X1 port map( A1 => n58, A2 => n67, ZN => mask_sh0(7));
   U208 : NAND2_X1 port map( A1 => n60, A2 => n69, ZN => mask_sh0(6));
   U209 : NAND2_X1 port map( A1 => n61, A2 => n71, ZN => mask_sh0(5));
   U210 : NAND2_X1 port map( A1 => n63, A2 => n74, ZN => mask_sh0(4));
   U211 : NAND2_X1 port map( A1 => n65, A2 => n75, ZN => mask_sh0(3));
   U212 : NAND2_X1 port map( A1 => n8, A2 => n77, ZN => mask_sh0(2));
   U213 : OAI21_X1 port map( B1 => n7, B2 => n92, A => n69, ZN => mask_sh6(0));
   U214 : NAND2_X1 port map( A1 => R1(37), A2 => n85, ZN => n76);
   U215 : NAND2_X1 port map( A1 => n37, A2 => n66, ZN => mask_sh0(17));
   U216 : NAND2_X1 port map( A1 => n65, A2 => n67, ZN => mask_sh2(5));
   U217 : NAND2_X1 port map( A1 => n67, A2 => n25, ZN => mask_sh6(1));
   U218 : NAND2_X1 port map( A1 => n8, A2 => n69, ZN => mask_sh2(4));
   U219 : NAND2_X1 port map( A1 => n10, A2 => n71, ZN => mask_sh2(3));
   U220 : NAND2_X1 port map( A1 => n12, A2 => n74, ZN => mask_sh2(2));
   U221 : NAND2_X1 port map( A1 => n15, A2 => n71, ZN => mask_sh3(2));
   U222 : NAND2_X1 port map( A1 => n15, A2 => n75, ZN => mask_sh2(1));
   U223 : NAND2_X1 port map( A1 => n67, A2 => n19, ZN => mask_sh5(2));
   U224 : NAND2_X1 port map( A1 => n17, A2 => n74, ZN => mask_sh3(1));
   U225 : NAND2_X1 port map( A1 => n19, A2 => n75, ZN => mask_sh3(0));
   U226 : NAND2_X1 port map( A1 => n17, A2 => n77, ZN => mask_sh2(0));
   U227 : NAND2_X1 port map( A1 => n69, A2 => n21, ZN => mask_sh5(1));
   U228 : NAND2_X1 port map( A1 => n71, A2 => n25, ZN => mask_sh5(0));
   U229 : INV_X1 port map( A => n88, ZN => n7);
   U230 : INV_X1 port map( A => n89, ZN => n78);
   U231 : NAND2_X1 port map( A1 => R1(7), A2 => n7, ZN => n67);
   U232 : NAND2_X1 port map( A1 => n28, A2 => n36, ZN => mask_sh5(26));
   U233 : NAND2_X1 port map( A1 => n36, A2 => n37, ZN => mask_sh7(24));
   U234 : NAND2_X1 port map( A1 => n38, A2 => n39, ZN => mask_sh7(23));
   U235 : NAND2_X1 port map( A1 => n51, A2 => n52, ZN => mask_sh7(17));
   U236 : NAND2_X1 port map( A1 => n53, A2 => n54, ZN => mask_sh7(16));
   U237 : NAND2_X1 port map( A1 => n55, A2 => n56, ZN => mask_sh7(15));
   U238 : NAND2_X1 port map( A1 => n57, A2 => n58, ZN => mask_sh7(14));
   U239 : NAND2_X1 port map( A1 => n59, A2 => n60, ZN => mask_sh7(13));
   U240 : NAND2_X1 port map( A1 => n61, A2 => n62, ZN => mask_sh7(12));
   U241 : NAND2_X1 port map( A1 => n63, A2 => n64, ZN => mask_sh7(11));
   U242 : NAND2_X1 port map( A1 => n10, A2 => n11, ZN => mask_sh7(8));
   U243 : NAND2_X1 port map( A1 => n12, A2 => n13, ZN => mask_sh7(7));
   U244 : NAND2_X1 port map( A1 => n16, A2 => n17, ZN => mask_sh7(5));
   U245 : NAND2_X1 port map( A1 => n18, A2 => n19, ZN => mask_sh7(4));
   U246 : NAND2_X1 port map( A1 => n20, A2 => n21, ZN => mask_sh7(3));
   U247 : NAND2_X1 port map( A1 => n24, A2 => n25, ZN => mask_sh7(2));
   U248 : OAI21_X1 port map( B1 => n78, B2 => n92, A => n46, ZN => mask_sh7(1))
                           ;
   U249 : OAI21_X1 port map( B1 => n88, B2 => n94, A => n22, ZN => mask_sh7(31)
                           );
   U250 : OAI21_X1 port map( B1 => n87, B2 => n93, A => n23, ZN => mask_sh7(30)
                           );
   U251 : NAND2_X1 port map( A1 => n26, A2 => n27, ZN => mask_sh7(29));
   U252 : NAND2_X1 port map( A1 => n28, A2 => n29, ZN => mask_sh7(28));
   U253 : NAND2_X1 port map( A1 => n30, A2 => n31, ZN => mask_sh7(27));
   U254 : OAI21_X1 port map( B1 => n78, B2 => n91, A => n67, ZN => mask_sh7(0))
                           ;
   U255 : NAND2_X1 port map( A1 => n23, A2 => n49, ZN => mask_sh1(24));
   U256 : NAND2_X1 port map( A1 => n26, A2 => n51, ZN => mask_sh1(23));
   U257 : NAND2_X1 port map( A1 => n28, A2 => n53, ZN => mask_sh1(22));
   U258 : NAND2_X1 port map( A1 => n30, A2 => n55, ZN => mask_sh1(21));
   U259 : NAND2_X1 port map( A1 => n32, A2 => n57, ZN => mask_sh1(20));
   U260 : NAND2_X1 port map( A1 => n34, A2 => n59, ZN => mask_sh1(19));
   U261 : NAND2_X1 port map( A1 => n37, A2 => n62, ZN => mask_sh1(18));
   U262 : NAND2_X1 port map( A1 => n39, A2 => n64, ZN => mask_sh1(17));
   U263 : NAND2_X1 port map( A1 => n41, A2 => n66, ZN => mask_sh1(16));
   U264 : NAND2_X1 port map( A1 => n9, A2 => n43, ZN => mask_sh1(15));
   U265 : NAND2_X1 port map( A1 => n11, A2 => n45, ZN => mask_sh1(14));
   U266 : NAND2_X1 port map( A1 => n13, A2 => n48, ZN => mask_sh1(13));
   U267 : NAND2_X1 port map( A1 => n14, A2 => n50, ZN => mask_sh1(12));
   U268 : NAND2_X1 port map( A1 => n16, A2 => n52, ZN => mask_sh1(11));
   U269 : NAND2_X1 port map( A1 => n18, A2 => n54, ZN => mask_sh1(10));
   U270 : NAND2_X1 port map( A1 => n20, A2 => n56, ZN => mask_sh1(9));
   U271 : NAND2_X1 port map( A1 => n24, A2 => n58, ZN => mask_sh1(8));
   U272 : NAND2_X1 port map( A1 => n46, A2 => n60, ZN => mask_sh1(7));
   U273 : NAND2_X1 port map( A1 => n61, A2 => n67, ZN => mask_sh1(6));
   U274 : NAND2_X1 port map( A1 => n63, A2 => n69, ZN => mask_sh1(5));
   U275 : NAND2_X1 port map( A1 => n65, A2 => n71, ZN => mask_sh1(4));
   U276 : NAND2_X1 port map( A1 => n8, A2 => n74, ZN => mask_sh1(3));
   U277 : NAND2_X1 port map( A1 => n10, A2 => n75, ZN => mask_sh1(2));
   U278 : NAND2_X1 port map( A1 => n12, A2 => n77, ZN => mask_sh1(1));
   U279 : OAI21_X1 port map( B1 => n7, B2 => n94, A => n35, ZN => mask_sh1(31))
                           ;
   U280 : NAND2_X1 port map( A1 => n36, A2 => n76, ZN => mask_sh1(30));
   U281 : NAND2_X1 port map( A1 => n38, A2 => n72, ZN => mask_sh1(29));
   U282 : NAND2_X1 port map( A1 => n40, A2 => n73, ZN => mask_sh1(28));
   U283 : NAND2_X1 port map( A1 => n42, A2 => n70, ZN => mask_sh1(27));
   U284 : NAND2_X1 port map( A1 => n44, A2 => n68, ZN => mask_sh1(26));
   U285 : NAND2_X1 port map( A1 => n22, A2 => n47, ZN => mask_sh1(25));
   U286 : OAI21_X1 port map( B1 => n88, B2 => n90, A => n12, ZN => mask_sh0(0))
                           ;
   U287 : INV_X1 port map( A => R1(38), ZN => n94);
   U288 : NAND2_X1 port map( A1 => R1(6), A2 => n7, ZN => n69);
   U289 : NAND2_X1 port map( A1 => R1(7), A2 => n86, ZN => n15);
   U290 : NAND2_X1 port map( A1 => R1(5), A2 => n7, ZN => n71);
   U291 : NAND2_X1 port map( A1 => R1(6), A2 => n83, ZN => n17);
   U292 : NAND2_X1 port map( A1 => R1(4), A2 => n7, ZN => n74);
   U293 : NAND2_X1 port map( A1 => R1(3), A2 => n7, ZN => n75);
   U294 : NAND2_X1 port map( A1 => R1(5), A2 => n80, ZN => n19);
   U295 : NAND2_X1 port map( A1 => R1(2), A2 => n7, ZN => n77);
   U296 : OAI21_X1 port map( B1 => n88, B2 => n91, A => n10, ZN => mask_sh0(1))
                           ;
   U297 : NAND2_X1 port map( A1 => R1(4), A2 => n79, ZN => n21);
   U298 : NAND2_X1 port map( A1 => R1(3), A2 => n79, ZN => n25);
   U299 : OAI21_X1 port map( B1 => n87, B2 => n91, A => n15, ZN => mask_sh1(0))
                           ;
   U300 : INV_X1 port map( A => R1(2), ZN => n92);
   U301 : BUF_X1 port map( A => n4, Z => n88);
   U302 : BUF_X1 port map( A => n2, Z => n82);
   U303 : BUF_X1 port map( A => n1, Z => n81);
   U304 : BUF_X1 port map( A => n1, Z => n79);
   U305 : BUF_X1 port map( A => n3, Z => n85);
   U306 : BUF_X1 port map( A => n2, Z => n84);
   U307 : BUF_X1 port map( A => n3, Z => n86);
   U308 : BUF_X1 port map( A => n2, Z => n83);
   U309 : BUF_X1 port map( A => n1, Z => n80);
   U310 : BUF_X1 port map( A => n3, Z => n87);
   U311 : BUF_X1 port map( A => n4, Z => n89);
   U312 : INV_X1 port map( A => R1(1), ZN => n91);
   U313 : INV_X1 port map( A => R1(0), ZN => n90);
   U314 : BUF_X1 port map( A => n5, Z => n3);
   U315 : BUF_X1 port map( A => n6, Z => n2);
   U316 : BUF_X1 port map( A => n6, Z => n1);
   U317 : BUF_X1 port map( A => n5, Z => n4);
   U318 : BUF_X1 port map( A => LnR, Z => n5);
   U319 : BUF_X1 port map( A => LnR, Z => n6);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_GENERIC_NBIT40 is

   port( A, B, C, D : in std_logic_vector (39 downto 0);  SEL : in 
         std_logic_vector (1 downto 0);  Y : out std_logic_vector (39 downto 0)
         );

end MUX41_GENERIC_NBIT40;

architecture SYN_structural of MUX41_GENERIC_NBIT40 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX41_33
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_34
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_35
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_36
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_37
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_38
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_39
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_40
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_41
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_42
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_43
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_44
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_45
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_46
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_47
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_48
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_49
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_50
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_51
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_52
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_53
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_54
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_55
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_56
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_57
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_58
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_59
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_60
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_61
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_62
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_63
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_64
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_65
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_66
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_67
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_68
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_69
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_70
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_71
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_72
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12 : std_logic;

begin
   
   MUXES_0 : MUX41_72 port map( A => A(0), B => B(0), C => C(0), D => D(0), 
                           S(1) => n9, S(0) => n3, Y => Y(0));
   MUXES_1 : MUX41_71 port map( A => A(1), B => B(1), C => C(1), D => D(1), 
                           S(1) => n9, S(0) => n3, Y => Y(1));
   MUXES_2 : MUX41_70 port map( A => A(2), B => B(2), C => C(2), D => D(2), 
                           S(1) => n9, S(0) => n3, Y => Y(2));
   MUXES_3 : MUX41_69 port map( A => A(3), B => B(3), C => C(3), D => D(3), 
                           S(1) => n9, S(0) => n3, Y => Y(3));
   MUXES_4 : MUX41_68 port map( A => A(4), B => B(4), C => C(4), D => D(4), 
                           S(1) => n9, S(0) => n3, Y => Y(4));
   MUXES_5 : MUX41_67 port map( A => A(5), B => B(5), C => C(5), D => D(5), 
                           S(1) => n9, S(0) => n3, Y => Y(5));
   MUXES_6 : MUX41_66 port map( A => A(6), B => B(6), C => C(6), D => D(6), 
                           S(1) => n9, S(0) => n3, Y => Y(6));
   MUXES_7 : MUX41_65 port map( A => A(7), B => B(7), C => C(7), D => D(7), 
                           S(1) => n9, S(0) => n3, Y => Y(7));
   MUXES_8 : MUX41_64 port map( A => A(8), B => B(8), C => C(8), D => D(8), 
                           S(1) => n9, S(0) => n3, Y => Y(8));
   MUXES_9 : MUX41_63 port map( A => A(9), B => B(9), C => C(9), D => D(9), 
                           S(1) => n9, S(0) => n3, Y => Y(9));
   MUXES_10 : MUX41_62 port map( A => A(10), B => B(10), C => C(10), D => D(10)
                           , S(1) => n9, S(0) => n3, Y => Y(10));
   MUXES_11 : MUX41_61 port map( A => A(11), B => B(11), C => C(11), D => D(11)
                           , S(1) => n9, S(0) => n4, Y => Y(11));
   MUXES_12 : MUX41_60 port map( A => A(12), B => B(12), C => C(12), D => D(12)
                           , S(1) => n10, S(0) => n4, Y => Y(12));
   MUXES_13 : MUX41_59 port map( A => A(13), B => B(13), C => C(13), D => D(13)
                           , S(1) => n10, S(0) => n4, Y => Y(13));
   MUXES_14 : MUX41_58 port map( A => A(14), B => B(14), C => C(14), D => D(14)
                           , S(1) => n10, S(0) => n4, Y => Y(14));
   MUXES_15 : MUX41_57 port map( A => A(15), B => B(15), C => C(15), D => D(15)
                           , S(1) => n10, S(0) => n4, Y => Y(15));
   MUXES_16 : MUX41_56 port map( A => A(16), B => B(16), C => C(16), D => D(16)
                           , S(1) => n10, S(0) => n4, Y => Y(16));
   MUXES_17 : MUX41_55 port map( A => A(17), B => B(17), C => C(17), D => D(17)
                           , S(1) => n10, S(0) => n4, Y => Y(17));
   MUXES_18 : MUX41_54 port map( A => A(18), B => B(18), C => C(18), D => D(18)
                           , S(1) => n10, S(0) => n4, Y => Y(18));
   MUXES_19 : MUX41_53 port map( A => A(19), B => B(19), C => C(19), D => D(19)
                           , S(1) => n10, S(0) => n4, Y => Y(19));
   MUXES_20 : MUX41_52 port map( A => A(20), B => B(20), C => C(20), D => D(20)
                           , S(1) => n10, S(0) => n4, Y => Y(20));
   MUXES_21 : MUX41_51 port map( A => A(21), B => B(21), C => C(21), D => D(21)
                           , S(1) => n10, S(0) => n4, Y => Y(21));
   MUXES_22 : MUX41_50 port map( A => A(22), B => B(22), C => C(22), D => D(22)
                           , S(1) => n10, S(0) => n5, Y => Y(22));
   MUXES_23 : MUX41_49 port map( A => A(23), B => B(23), C => C(23), D => D(23)
                           , S(1) => n10, S(0) => n5, Y => Y(23));
   MUXES_24 : MUX41_48 port map( A => A(24), B => B(24), C => C(24), D => D(24)
                           , S(1) => n11, S(0) => n5, Y => Y(24));
   MUXES_25 : MUX41_47 port map( A => A(25), B => B(25), C => C(25), D => D(25)
                           , S(1) => n11, S(0) => n5, Y => Y(25));
   MUXES_26 : MUX41_46 port map( A => A(26), B => B(26), C => C(26), D => D(26)
                           , S(1) => n11, S(0) => n5, Y => Y(26));
   MUXES_27 : MUX41_45 port map( A => A(27), B => B(27), C => C(27), D => D(27)
                           , S(1) => n11, S(0) => n5, Y => Y(27));
   MUXES_28 : MUX41_44 port map( A => A(28), B => B(28), C => C(28), D => D(28)
                           , S(1) => n11, S(0) => n5, Y => Y(28));
   MUXES_29 : MUX41_43 port map( A => A(29), B => B(29), C => C(29), D => D(29)
                           , S(1) => n11, S(0) => n5, Y => Y(29));
   MUXES_30 : MUX41_42 port map( A => A(30), B => B(30), C => C(30), D => D(30)
                           , S(1) => n11, S(0) => n5, Y => Y(30));
   MUXES_31 : MUX41_41 port map( A => A(31), B => B(31), C => C(31), D => D(31)
                           , S(1) => n11, S(0) => n5, Y => Y(31));
   MUXES_32 : MUX41_40 port map( A => A(32), B => B(32), C => C(32), D => D(32)
                           , S(1) => n11, S(0) => n5, Y => Y(32));
   MUXES_33 : MUX41_39 port map( A => A(33), B => B(33), C => C(33), D => D(33)
                           , S(1) => n11, S(0) => n6, Y => Y(33));
   MUXES_34 : MUX41_38 port map( A => A(34), B => B(34), C => C(34), D => D(34)
                           , S(1) => n11, S(0) => n6, Y => Y(34));
   MUXES_35 : MUX41_37 port map( A => A(35), B => B(35), C => C(35), D => D(35)
                           , S(1) => n11, S(0) => n6, Y => Y(35));
   MUXES_36 : MUX41_36 port map( A => A(36), B => B(36), C => C(36), D => D(36)
                           , S(1) => n12, S(0) => n6, Y => Y(36));
   MUXES_37 : MUX41_35 port map( A => A(37), B => B(37), C => C(37), D => D(37)
                           , S(1) => n12, S(0) => n6, Y => Y(37));
   MUXES_38 : MUX41_34 port map( A => A(38), B => B(38), C => C(38), D => D(38)
                           , S(1) => n12, S(0) => n6, Y => Y(38));
   MUXES_39 : MUX41_33 port map( A => A(39), B => B(39), C => C(39), D => D(39)
                           , S(1) => n12, S(0) => n6, Y => Y(39));
   U1 : BUF_X1 port map( A => n7, Z => n10);
   U2 : BUF_X1 port map( A => n7, Z => n9);
   U3 : BUF_X1 port map( A => n8, Z => n11);
   U4 : BUF_X1 port map( A => n8, Z => n12);
   U5 : BUF_X1 port map( A => n1, Z => n4);
   U6 : BUF_X1 port map( A => n1, Z => n3);
   U7 : BUF_X1 port map( A => n2, Z => n5);
   U8 : BUF_X1 port map( A => n2, Z => n6);
   U9 : BUF_X1 port map( A => SEL(0), Z => n1);
   U10 : BUF_X1 port map( A => SEL(1), Z => n7);
   U11 : BUF_X1 port map( A => SEL(0), Z => n2);
   U12 : BUF_X1 port map( A => SEL(1), Z => n8);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity mask_generator_NBITS32 is

   port( R1, R2 : in std_logic_vector (31 downto 0);  LnR, AnL, RnS : in 
         std_logic;  mask0, mask8, mask16, mask24 : out std_logic_vector (39 
         downto 0));

end mask_generator_NBITS32;

architecture SYN_structural of mask_generator_NBITS32 is

   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX41_GENERIC_NBIT8_1
      port( A, B, C, D : in std_logic_vector (7 downto 0);  SEL : in 
            std_logic_vector (1 downto 0);  Y : out std_logic_vector (7 downto 
            0));
   end component;
   
   component MUX21_GENERIC_NBIT8_1
      port( A, B : in std_logic_vector (7 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (7 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT8_2
      port( A, B : in std_logic_vector (7 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (7 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT8_3
      port( A, B : in std_logic_vector (7 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (7 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT8_4
      port( A, B : in std_logic_vector (7 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (7 downto 0));
   end component;
   
   component MUX41_GENERIC_NBIT8_2
      port( A, B, C, D : in std_logic_vector (7 downto 0);  SEL : in 
            std_logic_vector (1 downto 0);  Y : out std_logic_vector (7 downto 
            0));
   end component;
   
   component MUX21_GENERIC_NBIT8_5
      port( A, B : in std_logic_vector (7 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (7 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT8_6
      port( A, B : in std_logic_vector (7 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (7 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT8_7
      port( A, B : in std_logic_vector (7 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (7 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT8_8
      port( A, B : in std_logic_vector (7 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (7 downto 0));
   end component;
   
   component MUX41_GENERIC_NBIT8_3
      port( A, B, C, D : in std_logic_vector (7 downto 0);  SEL : in 
            std_logic_vector (1 downto 0);  Y : out std_logic_vector (7 downto 
            0));
   end component;
   
   component MUX21_GENERIC_NBIT8_9
      port( A, B : in std_logic_vector (7 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (7 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT8_10
      port( A, B : in std_logic_vector (7 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (7 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT8_11
      port( A, B : in std_logic_vector (7 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (7 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT8_12
      port( A, B : in std_logic_vector (7 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (7 downto 0));
   end component;
   
   component MUX41_GENERIC_NBIT8_0
      port( A, B, C, D : in std_logic_vector (7 downto 0);  SEL : in 
            std_logic_vector (1 downto 0);  Y : out std_logic_vector (7 downto 
            0));
   end component;
   
   component MUX21_GENERIC_NBIT8_13
      port( A, B : in std_logic_vector (7 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (7 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT8_14
      port( A, B : in std_logic_vector (7 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (7 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT8_15
      port( A, B : in std_logic_vector (7 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (7 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT8_16
      port( A, B : in std_logic_vector (7 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (7 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT8_0
      port( A, B : in std_logic_vector (7 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (7 downto 0));
   end component;
   
   signal X_Logic0_port, mask0_39_port, mask0_38_port, mask0_37_port, 
      mask0_36_port, mask0_35_port, mask0_34_port, mask0_33_port, mask0_32_port
      , mask0_31_port, mask0_30_port, mask0_29_port, mask0_28_port, 
      mask0_27_port, mask0_26_port, mask0_25_port, mask0_24_port, mask0_23_port
      , mask0_22_port, mask0_21_port, mask0_20_port, mask0_19_port, 
      mask0_18_port, mask0_17_port, mask0_16_port, mask0_15_port, mask0_14_port
      , mask0_13_port, mask0_12_port, mask0_11_port, mask0_10_port, 
      mask0_9_port, mask0_8_port, mask0_7_port, mask0_6_port, mask0_5_port, 
      mask0_4_port, mask0_3_port, mask0_2_port, mask0_1_port, mask0_0_port, 
      mask8_39_port, mask8_38_port, mask8_37_port, mask8_36_port, mask8_35_port
      , mask8_34_port, mask8_33_port, mask8_32_port, mask8_31_port, 
      mask8_30_port, mask8_29_port, mask8_28_port, mask8_27_port, mask8_26_port
      , mask8_25_port, mask8_24_port, mask8_23_port, mask8_22_port, 
      mask8_21_port, mask8_20_port, mask8_19_port, mask8_18_port, mask8_17_port
      , mask8_16_port, mask8_15_port, mask8_14_port, mask8_13_port, 
      mask8_12_port, mask8_11_port, mask8_10_port, mask8_9_port, mask8_8_port, 
      mask8_7_port, mask8_6_port, mask8_5_port, mask8_4_port, mask8_3_port, 
      mask8_2_port, mask8_1_port, mask8_0_port, mask16_39_port, mask16_38_port,
      mask16_37_port, mask16_36_port, mask16_35_port, mask16_34_port, 
      mask16_33_port, mask16_32_port, mask16_31_port, mask16_30_port, 
      mask16_29_port, mask16_28_port, mask16_27_port, mask16_26_port, 
      mask16_25_port, mask16_24_port, mask16_23_port, mask16_22_port, 
      mask16_21_port, mask16_20_port, mask16_19_port, mask16_18_port, 
      mask16_17_port, mask16_16_port, mask16_15_port, mask16_14_port, 
      mask16_13_port, mask16_12_port, mask16_11_port, mask16_10_port, 
      mask16_9_port, mask16_8_port, mask16_7_port, mask16_6_port, mask16_5_port
      , mask16_4_port, mask16_3_port, mask16_2_port, mask16_1_port, 
      mask16_0_port, shr_new_block_7_port, shr_new_block_6_port, 
      shr_new_block_5_port, shr_new_block_4_port, shr_new_block_3_port, 
      shr_new_block_2_port, shr_new_block_1_port, shr_new_block_0_port, n1, n2,
      n3, n4, n5, n6, n7, n8, n9 : std_logic;

begin
   mask0 <= ( mask0_39_port, mask0_38_port, mask0_37_port, mask0_36_port, 
      mask0_35_port, mask0_34_port, mask0_33_port, mask0_32_port, mask0_31_port
      , mask0_30_port, mask0_29_port, mask0_28_port, mask0_27_port, 
      mask0_26_port, mask0_25_port, mask0_24_port, mask0_23_port, mask0_22_port
      , mask0_21_port, mask0_20_port, mask0_19_port, mask0_18_port, 
      mask0_17_port, mask0_16_port, mask0_15_port, mask0_14_port, mask0_13_port
      , mask0_12_port, mask0_11_port, mask0_10_port, mask0_9_port, mask0_8_port
      , mask0_7_port, mask0_6_port, mask0_5_port, mask0_4_port, mask0_3_port, 
      mask0_2_port, mask0_1_port, mask0_0_port );
   mask8 <= ( mask8_39_port, mask8_38_port, mask8_37_port, mask8_36_port, 
      mask8_35_port, mask8_34_port, mask8_33_port, mask8_32_port, mask8_31_port
      , mask8_30_port, mask8_29_port, mask8_28_port, mask8_27_port, 
      mask8_26_port, mask8_25_port, mask8_24_port, mask8_23_port, mask8_22_port
      , mask8_21_port, mask8_20_port, mask8_19_port, mask8_18_port, 
      mask8_17_port, mask8_16_port, mask8_15_port, mask8_14_port, mask8_13_port
      , mask8_12_port, mask8_11_port, mask8_10_port, mask8_9_port, mask8_8_port
      , mask8_7_port, mask8_6_port, mask8_5_port, mask8_4_port, mask8_3_port, 
      mask8_2_port, mask8_1_port, mask8_0_port );
   mask16 <= ( mask16_39_port, mask16_38_port, mask16_37_port, mask16_36_port, 
      mask16_35_port, mask16_34_port, mask16_33_port, mask16_32_port, 
      mask16_31_port, mask16_30_port, mask16_29_port, mask16_28_port, 
      mask16_27_port, mask16_26_port, mask16_25_port, mask16_24_port, 
      mask16_23_port, mask16_22_port, mask16_21_port, mask16_20_port, 
      mask16_19_port, mask16_18_port, mask16_17_port, mask16_16_port, 
      mask16_15_port, mask16_14_port, mask16_13_port, mask16_12_port, 
      mask16_11_port, mask16_10_port, mask16_9_port, mask16_8_port, 
      mask16_7_port, mask16_6_port, mask16_5_port, mask16_4_port, mask16_3_port
      , mask16_2_port, mask16_1_port, mask16_0_port );
   
   X_Logic0_port <= '0';
   MUX_shift_type : MUX21_GENERIC_NBIT8_0 port map( A(7) => X_Logic0_port, A(6)
                           => X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(7) => n9, B(6) => n9, B(5) => n9, 
                           B(4) => n9, B(3) => n9, B(2) => n9, B(1) => n9, B(0)
                           => n9, SEL => AnL, Y(7) => shr_new_block_7_port, 
                           Y(6) => shr_new_block_6_port, Y(5) => 
                           shr_new_block_5_port, Y(4) => shr_new_block_4_port, 
                           Y(3) => shr_new_block_3_port, Y(2) => 
                           shr_new_block_2_port, Y(1) => shr_new_block_1_port, 
                           Y(0) => shr_new_block_0_port);
   MUX_mask0_LSB_0_0 : MUX21_GENERIC_NBIT8_16 port map( A(7) => R1(7), A(6) => 
                           R1(6), A(5) => R1(5), A(4) => R1(4), A(3) => R1(3), 
                           A(2) => R1(2), A(1) => R1(1), A(0) => R1(0), B(7) =>
                           X_Logic0_port, B(6) => X_Logic0_port, B(5) => 
                           X_Logic0_port, B(4) => X_Logic0_port, B(3) => 
                           X_Logic0_port, B(2) => X_Logic0_port, B(1) => 
                           X_Logic0_port, B(0) => X_Logic0_port, SEL => n3, 
                           Y(7) => mask0_7_port, Y(6) => mask0_6_port, Y(5) => 
                           mask0_5_port, Y(4) => mask0_4_port, Y(3) => 
                           mask0_3_port, Y(2) => mask0_2_port, Y(1) => 
                           mask0_1_port, Y(0) => mask0_0_port);
   MUX_mask0_0_1 : MUX21_GENERIC_NBIT8_15 port map( A(7) => R1(15), A(6) => 
                           R1(14), A(5) => R1(13), A(4) => R1(12), A(3) => 
                           R1(11), A(2) => R1(10), A(1) => R1(9), A(0) => R1(8)
                           , B(7) => R1(7), B(6) => R1(6), B(5) => R1(5), B(4) 
                           => R1(4), B(3) => R1(3), B(2) => R1(2), B(1) => 
                           R1(1), B(0) => R1(0), SEL => n8, Y(7) => 
                           mask0_15_port, Y(6) => mask0_14_port, Y(5) => 
                           mask0_13_port, Y(4) => mask0_12_port, Y(3) => 
                           mask0_11_port, Y(2) => mask0_10_port, Y(1) => 
                           mask0_9_port, Y(0) => mask0_8_port);
   MUX_mask0_0_2 : MUX21_GENERIC_NBIT8_14 port map( A(7) => R1(23), A(6) => 
                           R1(22), A(5) => R1(21), A(4) => R1(20), A(3) => 
                           R1(19), A(2) => R1(18), A(1) => R1(17), A(0) => 
                           R1(16), B(7) => R1(15), B(6) => R1(14), B(5) => 
                           R1(13), B(4) => R1(12), B(3) => R1(11), B(2) => 
                           R1(10), B(1) => R1(9), B(0) => R1(8), SEL => n8, 
                           Y(7) => mask0_23_port, Y(6) => mask0_22_port, Y(5) 
                           => mask0_21_port, Y(4) => mask0_20_port, Y(3) => 
                           mask0_19_port, Y(2) => mask0_18_port, Y(1) => 
                           mask0_17_port, Y(0) => mask0_16_port);
   MUX_mask0_0_3 : MUX21_GENERIC_NBIT8_13 port map( A(7) => n9, A(6) => R1(30),
                           A(5) => R1(29), A(4) => R1(28), A(3) => R1(27), A(2)
                           => R1(26), A(1) => R1(25), A(0) => R1(24), B(7) => 
                           R1(23), B(6) => R1(22), B(5) => R1(21), B(4) => 
                           R1(20), B(3) => R1(19), B(2) => R1(18), B(1) => 
                           R1(17), B(0) => R1(16), SEL => n7, Y(7) => 
                           mask0_31_port, Y(6) => mask0_30_port, Y(5) => 
                           mask0_29_port, Y(4) => mask0_28_port, Y(3) => 
                           mask0_27_port, Y(2) => mask0_26_port, Y(1) => 
                           mask0_25_port, Y(0) => mask0_24_port);
   MUX_mask_MSB_0_4 : MUX41_GENERIC_NBIT8_0 port map( A(7) => 
                           shr_new_block_7_port, A(6) => shr_new_block_6_port, 
                           A(5) => shr_new_block_5_port, A(4) => 
                           shr_new_block_4_port, A(3) => shr_new_block_3_port, 
                           A(2) => shr_new_block_2_port, A(1) => 
                           shr_new_block_1_port, A(0) => shr_new_block_0_port, 
                           B(7) => R1(7), B(6) => R1(6), B(5) => R1(5), B(4) =>
                           R1(4), B(3) => R1(3), B(2) => R1(2), B(1) => R1(1), 
                           B(0) => R1(0), C(7) => n9, C(6) => R1(30), C(5) => 
                           R1(29), C(4) => R1(28), C(3) => R1(27), C(2) => 
                           R1(26), C(1) => R1(25), C(0) => R1(24), D(7) => n9, 
                           D(6) => R1(30), D(5) => R1(29), D(4) => R1(28), D(3)
                           => R1(27), D(2) => R1(26), D(1) => R1(25), D(0) => 
                           R1(24), SEL(1) => n3, SEL(0) => n1, Y(7) => 
                           mask0_39_port, Y(6) => mask0_38_port, Y(5) => 
                           mask0_37_port, Y(4) => mask0_36_port, Y(3) => 
                           mask0_35_port, Y(2) => mask0_34_port, Y(1) => 
                           mask0_33_port, Y(0) => mask0_32_port);
   MUX_mask_LSB_1_0 : MUX21_GENERIC_NBIT8_12 port map( A(7) => mask0_15_port, 
                           A(6) => mask0_14_port, A(5) => mask0_13_port, A(4) 
                           => mask0_12_port, A(3) => mask0_11_port, A(2) => 
                           mask0_10_port, A(1) => mask0_9_port, A(0) => 
                           mask0_8_port, B(7) => X_Logic0_port, B(6) => 
                           X_Logic0_port, B(5) => X_Logic0_port, B(4) => 
                           X_Logic0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           X_Logic0_port, SEL => n7, Y(7) => mask8_7_port, Y(6)
                           => mask8_6_port, Y(5) => mask8_5_port, Y(4) => 
                           mask8_4_port, Y(3) => mask8_3_port, Y(2) => 
                           mask8_2_port, Y(1) => mask8_1_port, Y(0) => 
                           mask8_0_port);
   MUX_mask_1_1 : MUX21_GENERIC_NBIT8_11 port map( A(7) => mask0_23_port, A(6) 
                           => mask0_22_port, A(5) => mask0_21_port, A(4) => 
                           mask0_20_port, A(3) => mask0_19_port, A(2) => 
                           mask0_18_port, A(1) => mask0_17_port, A(0) => 
                           mask0_16_port, B(7) => mask0_7_port, B(6) => 
                           mask0_6_port, B(5) => mask0_5_port, B(4) => 
                           mask0_4_port, B(3) => mask0_3_port, B(2) => 
                           mask0_2_port, B(1) => mask0_1_port, B(0) => 
                           mask0_0_port, SEL => n7, Y(7) => mask8_15_port, Y(6)
                           => mask8_14_port, Y(5) => mask8_13_port, Y(4) => 
                           mask8_12_port, Y(3) => mask8_11_port, Y(2) => 
                           mask8_10_port, Y(1) => mask8_9_port, Y(0) => 
                           mask8_8_port);
   MUX_mask_1_2 : MUX21_GENERIC_NBIT8_10 port map( A(7) => mask0_31_port, A(6) 
                           => mask0_30_port, A(5) => mask0_29_port, A(4) => 
                           mask0_28_port, A(3) => mask0_27_port, A(2) => 
                           mask0_26_port, A(1) => mask0_25_port, A(0) => 
                           mask0_24_port, B(7) => mask0_15_port, B(6) => 
                           mask0_14_port, B(5) => mask0_13_port, B(4) => 
                           mask0_12_port, B(3) => mask0_11_port, B(2) => 
                           mask0_10_port, B(1) => mask0_9_port, B(0) => 
                           mask0_8_port, SEL => n6, Y(7) => mask8_23_port, Y(6)
                           => mask8_22_port, Y(5) => mask8_21_port, Y(4) => 
                           mask8_20_port, Y(3) => mask8_19_port, Y(2) => 
                           mask8_18_port, Y(1) => mask8_17_port, Y(0) => 
                           mask8_16_port);
   MUX_mask_1_3 : MUX21_GENERIC_NBIT8_9 port map( A(7) => mask0_39_port, A(6) 
                           => mask0_38_port, A(5) => mask0_37_port, A(4) => 
                           mask0_36_port, A(3) => mask0_35_port, A(2) => 
                           mask0_34_port, A(1) => mask0_33_port, A(0) => 
                           mask0_32_port, B(7) => mask0_23_port, B(6) => 
                           mask0_22_port, B(5) => mask0_21_port, B(4) => 
                           mask0_20_port, B(3) => mask0_19_port, B(2) => 
                           mask0_18_port, B(1) => mask0_17_port, B(0) => 
                           mask0_16_port, SEL => n6, Y(7) => mask8_31_port, 
                           Y(6) => mask8_30_port, Y(5) => mask8_29_port, Y(4) 
                           => mask8_28_port, Y(3) => mask8_27_port, Y(2) => 
                           mask8_26_port, Y(1) => mask8_25_port, Y(0) => 
                           mask8_24_port);
   MUX_mask_MSB_1_4 : MUX41_GENERIC_NBIT8_3 port map( A(7) => 
                           shr_new_block_7_port, A(6) => shr_new_block_6_port, 
                           A(5) => shr_new_block_5_port, A(4) => 
                           shr_new_block_4_port, A(3) => shr_new_block_3_port, 
                           A(2) => shr_new_block_2_port, A(1) => 
                           shr_new_block_1_port, A(0) => shr_new_block_0_port, 
                           B(7) => mask0_15_port, B(6) => mask0_14_port, B(5) 
                           => mask0_13_port, B(4) => mask0_12_port, B(3) => 
                           mask0_11_port, B(2) => mask0_10_port, B(1) => 
                           mask0_9_port, B(0) => mask0_8_port, C(7) => 
                           mask0_31_port, C(6) => mask0_30_port, C(5) => 
                           mask0_29_port, C(4) => mask0_28_port, C(3) => 
                           mask0_27_port, C(2) => mask0_26_port, C(1) => 
                           mask0_25_port, C(0) => mask0_24_port, D(7) => 
                           mask0_31_port, D(6) => mask0_30_port, D(5) => 
                           mask0_29_port, D(4) => mask0_28_port, D(3) => 
                           mask0_27_port, D(2) => mask0_26_port, D(1) => 
                           mask0_25_port, D(0) => mask0_24_port, SEL(1) => n2, 
                           SEL(0) => n1, Y(7) => mask8_39_port, Y(6) => 
                           mask8_38_port, Y(5) => mask8_37_port, Y(4) => 
                           mask8_36_port, Y(3) => mask8_35_port, Y(2) => 
                           mask8_34_port, Y(1) => mask8_33_port, Y(0) => 
                           mask8_32_port);
   MUX_mask_LSB_2_0 : MUX21_GENERIC_NBIT8_8 port map( A(7) => mask8_15_port, 
                           A(6) => mask8_14_port, A(5) => mask8_13_port, A(4) 
                           => mask8_12_port, A(3) => mask8_11_port, A(2) => 
                           mask8_10_port, A(1) => mask8_9_port, A(0) => 
                           mask8_8_port, B(7) => X_Logic0_port, B(6) => 
                           X_Logic0_port, B(5) => X_Logic0_port, B(4) => 
                           X_Logic0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           X_Logic0_port, SEL => n6, Y(7) => mask16_7_port, 
                           Y(6) => mask16_6_port, Y(5) => mask16_5_port, Y(4) 
                           => mask16_4_port, Y(3) => mask16_3_port, Y(2) => 
                           mask16_2_port, Y(1) => mask16_1_port, Y(0) => 
                           mask16_0_port);
   MUX_mask_2_1 : MUX21_GENERIC_NBIT8_7 port map( A(7) => mask8_23_port, A(6) 
                           => mask8_22_port, A(5) => mask8_21_port, A(4) => 
                           mask8_20_port, A(3) => mask8_19_port, A(2) => 
                           mask8_18_port, A(1) => mask8_17_port, A(0) => 
                           mask8_16_port, B(7) => mask8_7_port, B(6) => 
                           mask8_6_port, B(5) => mask8_5_port, B(4) => 
                           mask8_4_port, B(3) => mask8_3_port, B(2) => 
                           mask8_2_port, B(1) => mask8_1_port, B(0) => 
                           mask8_0_port, SEL => n5, Y(7) => mask16_15_port, 
                           Y(6) => mask16_14_port, Y(5) => mask16_13_port, Y(4)
                           => mask16_12_port, Y(3) => mask16_11_port, Y(2) => 
                           mask16_10_port, Y(1) => mask16_9_port, Y(0) => 
                           mask16_8_port);
   MUX_mask_2_2 : MUX21_GENERIC_NBIT8_6 port map( A(7) => mask8_31_port, A(6) 
                           => mask8_30_port, A(5) => mask8_29_port, A(4) => 
                           mask8_28_port, A(3) => mask8_27_port, A(2) => 
                           mask8_26_port, A(1) => mask8_25_port, A(0) => 
                           mask8_24_port, B(7) => mask8_15_port, B(6) => 
                           mask8_14_port, B(5) => mask8_13_port, B(4) => 
                           mask8_12_port, B(3) => mask8_11_port, B(2) => 
                           mask8_10_port, B(1) => mask8_9_port, B(0) => 
                           mask8_8_port, SEL => n5, Y(7) => mask16_23_port, 
                           Y(6) => mask16_22_port, Y(5) => mask16_21_port, Y(4)
                           => mask16_20_port, Y(3) => mask16_19_port, Y(2) => 
                           mask16_18_port, Y(1) => mask16_17_port, Y(0) => 
                           mask16_16_port);
   MUX_mask_2_3 : MUX21_GENERIC_NBIT8_5 port map( A(7) => mask8_39_port, A(6) 
                           => mask8_38_port, A(5) => mask8_37_port, A(4) => 
                           mask8_36_port, A(3) => mask8_35_port, A(2) => 
                           mask8_34_port, A(1) => mask8_33_port, A(0) => 
                           mask8_32_port, B(7) => mask8_23_port, B(6) => 
                           mask8_22_port, B(5) => mask8_21_port, B(4) => 
                           mask8_20_port, B(3) => mask8_19_port, B(2) => 
                           mask8_18_port, B(1) => mask8_17_port, B(0) => 
                           mask8_16_port, SEL => n4, Y(7) => mask16_31_port, 
                           Y(6) => mask16_30_port, Y(5) => mask16_29_port, Y(4)
                           => mask16_28_port, Y(3) => mask16_27_port, Y(2) => 
                           mask16_26_port, Y(1) => mask16_25_port, Y(0) => 
                           mask16_24_port);
   MUX_mask_MSB_2_4 : MUX41_GENERIC_NBIT8_2 port map( A(7) => 
                           shr_new_block_7_port, A(6) => shr_new_block_6_port, 
                           A(5) => shr_new_block_5_port, A(4) => 
                           shr_new_block_4_port, A(3) => shr_new_block_3_port, 
                           A(2) => shr_new_block_2_port, A(1) => 
                           shr_new_block_1_port, A(0) => shr_new_block_0_port, 
                           B(7) => mask8_15_port, B(6) => mask8_14_port, B(5) 
                           => mask8_13_port, B(4) => mask8_12_port, B(3) => 
                           mask8_11_port, B(2) => mask8_10_port, B(1) => 
                           mask8_9_port, B(0) => mask8_8_port, C(7) => 
                           mask8_31_port, C(6) => mask8_30_port, C(5) => 
                           mask8_29_port, C(4) => mask8_28_port, C(3) => 
                           mask8_27_port, C(2) => mask8_26_port, C(1) => 
                           mask8_25_port, C(0) => mask8_24_port, D(7) => 
                           mask8_31_port, D(6) => mask8_30_port, D(5) => 
                           mask8_29_port, D(4) => mask8_28_port, D(3) => 
                           mask8_27_port, D(2) => mask8_26_port, D(1) => 
                           mask8_25_port, D(0) => mask8_24_port, SEL(1) => n2, 
                           SEL(0) => n1, Y(7) => mask16_39_port, Y(6) => 
                           mask16_38_port, Y(5) => mask16_37_port, Y(4) => 
                           mask16_36_port, Y(3) => mask16_35_port, Y(2) => 
                           mask16_34_port, Y(1) => mask16_33_port, Y(0) => 
                           mask16_32_port);
   MUX_mask_LSB_3_0 : MUX21_GENERIC_NBIT8_4 port map( A(7) => mask16_15_port, 
                           A(6) => mask16_14_port, A(5) => mask16_13_port, A(4)
                           => mask16_12_port, A(3) => mask16_11_port, A(2) => 
                           mask16_10_port, A(1) => mask16_9_port, A(0) => 
                           mask16_8_port, B(7) => X_Logic0_port, B(6) => 
                           X_Logic0_port, B(5) => X_Logic0_port, B(4) => 
                           X_Logic0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           X_Logic0_port, SEL => n5, Y(7) => mask24(7), Y(6) =>
                           mask24(6), Y(5) => mask24(5), Y(4) => mask24(4), 
                           Y(3) => mask24(3), Y(2) => mask24(2), Y(1) => 
                           mask24(1), Y(0) => mask24(0));
   MUX_mask_3_1 : MUX21_GENERIC_NBIT8_3 port map( A(7) => mask16_23_port, A(6) 
                           => mask16_22_port, A(5) => mask16_21_port, A(4) => 
                           mask16_20_port, A(3) => mask16_19_port, A(2) => 
                           mask16_18_port, A(1) => mask16_17_port, A(0) => 
                           mask16_16_port, B(7) => mask16_7_port, B(6) => 
                           mask16_6_port, B(5) => mask16_5_port, B(4) => 
                           mask16_4_port, B(3) => mask16_3_port, B(2) => 
                           mask16_2_port, B(1) => mask16_1_port, B(0) => 
                           mask16_0_port, SEL => n4, Y(7) => mask24(15), Y(6) 
                           => mask24(14), Y(5) => mask24(13), Y(4) => 
                           mask24(12), Y(3) => mask24(11), Y(2) => mask24(10), 
                           Y(1) => mask24(9), Y(0) => mask24(8));
   MUX_mask_3_2 : MUX21_GENERIC_NBIT8_2 port map( A(7) => mask16_31_port, A(6) 
                           => mask16_30_port, A(5) => mask16_29_port, A(4) => 
                           mask16_28_port, A(3) => mask16_27_port, A(2) => 
                           mask16_26_port, A(1) => mask16_25_port, A(0) => 
                           mask16_24_port, B(7) => mask16_15_port, B(6) => 
                           mask16_14_port, B(5) => mask16_13_port, B(4) => 
                           mask16_12_port, B(3) => mask16_11_port, B(2) => 
                           mask16_10_port, B(1) => mask16_9_port, B(0) => 
                           mask16_8_port, SEL => n4, Y(7) => mask24(23), Y(6) 
                           => mask24(22), Y(5) => mask24(21), Y(4) => 
                           mask24(20), Y(3) => mask24(19), Y(2) => mask24(18), 
                           Y(1) => mask24(17), Y(0) => mask24(16));
   MUX_mask_3_3 : MUX21_GENERIC_NBIT8_1 port map( A(7) => mask16_39_port, A(6) 
                           => mask16_38_port, A(5) => mask16_37_port, A(4) => 
                           mask16_36_port, A(3) => mask16_35_port, A(2) => 
                           mask16_34_port, A(1) => mask16_33_port, A(0) => 
                           mask16_32_port, B(7) => mask16_23_port, B(6) => 
                           mask16_22_port, B(5) => mask16_21_port, B(4) => 
                           mask16_20_port, B(3) => mask16_19_port, B(2) => 
                           mask16_18_port, B(1) => mask16_17_port, B(0) => 
                           mask16_16_port, SEL => n3, Y(7) => mask24(31), Y(6) 
                           => mask24(30), Y(5) => mask24(29), Y(4) => 
                           mask24(28), Y(3) => mask24(27), Y(2) => mask24(26), 
                           Y(1) => mask24(25), Y(0) => mask24(24));
   MUX_mask_MSB_3_4 : MUX41_GENERIC_NBIT8_1 port map( A(7) => 
                           shr_new_block_7_port, A(6) => shr_new_block_6_port, 
                           A(5) => shr_new_block_5_port, A(4) => 
                           shr_new_block_4_port, A(3) => shr_new_block_3_port, 
                           A(2) => shr_new_block_2_port, A(1) => 
                           shr_new_block_1_port, A(0) => shr_new_block_0_port, 
                           B(7) => mask16_15_port, B(6) => mask16_14_port, B(5)
                           => mask16_13_port, B(4) => mask16_12_port, B(3) => 
                           mask16_11_port, B(2) => mask16_10_port, B(1) => 
                           mask16_9_port, B(0) => mask16_8_port, C(7) => 
                           mask16_31_port, C(6) => mask16_30_port, C(5) => 
                           mask16_29_port, C(4) => mask16_28_port, C(3) => 
                           mask16_27_port, C(2) => mask16_26_port, C(1) => 
                           mask16_25_port, C(0) => mask16_24_port, D(7) => 
                           mask16_31_port, D(6) => mask16_30_port, D(5) => 
                           mask16_29_port, D(4) => mask16_28_port, D(3) => 
                           mask16_27_port, D(2) => mask16_26_port, D(1) => 
                           mask16_25_port, D(0) => mask16_24_port, SEL(1) => n2
                           , SEL(0) => n1, Y(7) => mask24(39), Y(6) => 
                           mask24(38), Y(5) => mask24(37), Y(4) => mask24(36), 
                           Y(3) => mask24(35), Y(2) => mask24(34), Y(1) => 
                           mask24(33), Y(0) => mask24(32));
   U2 : BUF_X2 port map( A => LnR, Z => n2);
   U3 : BUF_X2 port map( A => LnR, Z => n4);
   U4 : BUF_X2 port map( A => LnR, Z => n6);
   U5 : BUF_X2 port map( A => LnR, Z => n5);
   U6 : BUF_X2 port map( A => LnR, Z => n7);
   U7 : BUF_X2 port map( A => LnR, Z => n3);
   U8 : BUF_X1 port map( A => R1(31), Z => n9);
   U9 : BUF_X2 port map( A => LnR, Z => n8);
   U10 : BUF_X2 port map( A => RnS, Z => n1);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT4_0 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end MUX21_GENERIC_NBIT4_0;

architecture SYN_structural of MUX21_GENERIC_NBIT4_0 is

   component MUX21_389
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_390
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_391
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_392
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_392 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_391 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_390 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_389 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity RCA_GEN_NBIT4_0 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_0;

architecture SYN_STRUCTURAL of RCA_GEN_NBIT4_0 is

   component FA_509
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_510
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_511
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_0
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_0 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_511 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_510 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_509 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity P4_ADDER_NBIT64_0 is

   port( A, B : in std_logic_vector (63 downto 0);  Cin : in std_logic;  S : 
         out std_logic_vector (63 downto 0);  Cout, ovf : out std_logic);

end P4_ADDER_NBIT64_0;

architecture SYN_STRUCTURAL of P4_ADDER_NBIT64_0 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component sum_generator_n_bit64_n_CSB16_0
      port( A, B : in std_logic_vector (63 downto 0);  C_in : in 
            std_logic_vector (15 downto 0);  S : out std_logic_vector (63 
            downto 0));
   end component;
   
   component CARRY_GENERATOR_NBIT64_NBIT_PER_BLOCK4_0
      port( A, B : in std_logic_vector (63 downto 0);  Cin : in std_logic;  Co 
            : out std_logic_vector (15 downto 0));
   end component;
   
   component my_xor_129
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_130
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_131
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_132
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_133
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_134
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_135
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_136
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_137
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_138
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_139
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_140
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_141
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_142
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_143
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_144
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_145
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_146
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_147
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_148
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_149
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_150
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_151
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_152
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_153
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_154
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_155
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_156
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_157
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_158
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_159
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_160
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_161
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_162
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_163
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_164
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_165
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_166
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_167
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_168
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_169
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_170
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_171
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_172
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_173
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_174
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_175
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_176
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_177
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_178
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_179
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_180
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_181
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_182
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_183
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_184
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_185
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_186
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_187
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_188
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_189
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_190
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_191
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_192
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal S_63_port, S_62_port, S_61_port, S_60_port, S_59_port, S_58_port, 
      S_57_port, S_56_port, S_55_port, S_54_port, S_53_port, S_52_port, 
      S_51_port, S_50_port, S_49_port, S_48_port, S_47_port, S_46_port, 
      S_45_port, S_44_port, S_43_port, S_42_port, S_41_port, S_40_port, 
      S_39_port, S_38_port, S_37_port, S_36_port, S_35_port, S_34_port, 
      S_33_port, S_32_port, S_31_port, S_30_port, S_29_port, S_28_port, 
      S_27_port, S_26_port, S_25_port, S_24_port, S_23_port, S_22_port, 
      S_21_port, S_20_port, S_19_port, S_18_port, S_17_port, S_16_port, 
      S_15_port, S_14_port, S_13_port, S_12_port, S_11_port, S_10_port, 
      S_9_port, S_8_port, S_7_port, S_6_port, S_5_port, S_4_port, S_3_port, 
      S_2_port, S_1_port, S_0_port, xor_b_63_port, xor_b_62_port, xor_b_61_port
      , xor_b_60_port, xor_b_59_port, xor_b_58_port, xor_b_57_port, 
      xor_b_56_port, xor_b_55_port, xor_b_54_port, xor_b_53_port, xor_b_52_port
      , xor_b_51_port, xor_b_50_port, xor_b_49_port, xor_b_48_port, 
      xor_b_47_port, xor_b_46_port, xor_b_45_port, xor_b_44_port, xor_b_43_port
      , xor_b_42_port, xor_b_41_port, xor_b_40_port, xor_b_39_port, 
      xor_b_38_port, xor_b_37_port, xor_b_36_port, xor_b_35_port, xor_b_34_port
      , xor_b_33_port, xor_b_32_port, xor_b_31_port, xor_b_30_port, 
      xor_b_29_port, xor_b_28_port, xor_b_27_port, xor_b_26_port, xor_b_25_port
      , xor_b_24_port, xor_b_23_port, xor_b_22_port, xor_b_21_port, 
      xor_b_20_port, xor_b_19_port, xor_b_18_port, xor_b_17_port, xor_b_16_port
      , xor_b_15_port, xor_b_14_port, xor_b_13_port, xor_b_12_port, 
      xor_b_11_port, xor_b_10_port, xor_b_9_port, xor_b_8_port, xor_b_7_port, 
      xor_b_6_port, xor_b_5_port, xor_b_4_port, xor_b_3_port, xor_b_2_port, 
      xor_b_1_port, xor_b_0_port, carry_14_port, carry_13_port, carry_12_port, 
      carry_11_port, carry_10_port, carry_9_port, carry_8_port, carry_7_port, 
      carry_6_port, carry_5_port, carry_4_port, carry_3_port, carry_2_port, 
      carry_1_port, carry_0_port, n1, n2 : std_logic;

begin
   S <= ( S_63_port, S_62_port, S_61_port, S_60_port, S_59_port, S_58_port, 
      S_57_port, S_56_port, S_55_port, S_54_port, S_53_port, S_52_port, 
      S_51_port, S_50_port, S_49_port, S_48_port, S_47_port, S_46_port, 
      S_45_port, S_44_port, S_43_port, S_42_port, S_41_port, S_40_port, 
      S_39_port, S_38_port, S_37_port, S_36_port, S_35_port, S_34_port, 
      S_33_port, S_32_port, S_31_port, S_30_port, S_29_port, S_28_port, 
      S_27_port, S_26_port, S_25_port, S_24_port, S_23_port, S_22_port, 
      S_21_port, S_20_port, S_19_port, S_18_port, S_17_port, S_16_port, 
      S_15_port, S_14_port, S_13_port, S_12_port, S_11_port, S_10_port, 
      S_9_port, S_8_port, S_7_port, S_6_port, S_5_port, S_4_port, S_3_port, 
      S_2_port, S_1_port, S_0_port );
   
   U3 : XOR2_X1 port map( A => xor_b_63_port, B => A(63), Z => n2);
   bc_xor_63 : my_xor_192 port map( A => B(63), B => Cin, xor_out => 
                           xor_b_63_port);
   bc_xor_62 : my_xor_191 port map( A => B(62), B => Cin, xor_out => 
                           xor_b_62_port);
   bc_xor_61 : my_xor_190 port map( A => B(61), B => Cin, xor_out => 
                           xor_b_61_port);
   bc_xor_60 : my_xor_189 port map( A => B(60), B => Cin, xor_out => 
                           xor_b_60_port);
   bc_xor_59 : my_xor_188 port map( A => B(59), B => Cin, xor_out => 
                           xor_b_59_port);
   bc_xor_58 : my_xor_187 port map( A => B(58), B => Cin, xor_out => 
                           xor_b_58_port);
   bc_xor_57 : my_xor_186 port map( A => B(57), B => Cin, xor_out => 
                           xor_b_57_port);
   bc_xor_56 : my_xor_185 port map( A => B(56), B => Cin, xor_out => 
                           xor_b_56_port);
   bc_xor_55 : my_xor_184 port map( A => B(55), B => Cin, xor_out => 
                           xor_b_55_port);
   bc_xor_54 : my_xor_183 port map( A => B(54), B => Cin, xor_out => 
                           xor_b_54_port);
   bc_xor_53 : my_xor_182 port map( A => B(53), B => Cin, xor_out => 
                           xor_b_53_port);
   bc_xor_52 : my_xor_181 port map( A => B(52), B => Cin, xor_out => 
                           xor_b_52_port);
   bc_xor_51 : my_xor_180 port map( A => B(51), B => Cin, xor_out => 
                           xor_b_51_port);
   bc_xor_50 : my_xor_179 port map( A => B(50), B => Cin, xor_out => 
                           xor_b_50_port);
   bc_xor_49 : my_xor_178 port map( A => B(49), B => Cin, xor_out => 
                           xor_b_49_port);
   bc_xor_48 : my_xor_177 port map( A => B(48), B => Cin, xor_out => 
                           xor_b_48_port);
   bc_xor_47 : my_xor_176 port map( A => B(47), B => Cin, xor_out => 
                           xor_b_47_port);
   bc_xor_46 : my_xor_175 port map( A => B(46), B => Cin, xor_out => 
                           xor_b_46_port);
   bc_xor_45 : my_xor_174 port map( A => B(45), B => Cin, xor_out => 
                           xor_b_45_port);
   bc_xor_44 : my_xor_173 port map( A => B(44), B => Cin, xor_out => 
                           xor_b_44_port);
   bc_xor_43 : my_xor_172 port map( A => B(43), B => Cin, xor_out => 
                           xor_b_43_port);
   bc_xor_42 : my_xor_171 port map( A => B(42), B => Cin, xor_out => 
                           xor_b_42_port);
   bc_xor_41 : my_xor_170 port map( A => B(41), B => Cin, xor_out => 
                           xor_b_41_port);
   bc_xor_40 : my_xor_169 port map( A => B(40), B => Cin, xor_out => 
                           xor_b_40_port);
   bc_xor_39 : my_xor_168 port map( A => B(39), B => Cin, xor_out => 
                           xor_b_39_port);
   bc_xor_38 : my_xor_167 port map( A => B(38), B => Cin, xor_out => 
                           xor_b_38_port);
   bc_xor_37 : my_xor_166 port map( A => B(37), B => Cin, xor_out => 
                           xor_b_37_port);
   bc_xor_36 : my_xor_165 port map( A => B(36), B => Cin, xor_out => 
                           xor_b_36_port);
   bc_xor_35 : my_xor_164 port map( A => B(35), B => Cin, xor_out => 
                           xor_b_35_port);
   bc_xor_34 : my_xor_163 port map( A => B(34), B => Cin, xor_out => 
                           xor_b_34_port);
   bc_xor_33 : my_xor_162 port map( A => B(33), B => Cin, xor_out => 
                           xor_b_33_port);
   bc_xor_32 : my_xor_161 port map( A => B(32), B => Cin, xor_out => 
                           xor_b_32_port);
   bc_xor_31 : my_xor_160 port map( A => B(31), B => Cin, xor_out => 
                           xor_b_31_port);
   bc_xor_30 : my_xor_159 port map( A => B(30), B => Cin, xor_out => 
                           xor_b_30_port);
   bc_xor_29 : my_xor_158 port map( A => B(29), B => Cin, xor_out => 
                           xor_b_29_port);
   bc_xor_28 : my_xor_157 port map( A => B(28), B => Cin, xor_out => 
                           xor_b_28_port);
   bc_xor_27 : my_xor_156 port map( A => B(27), B => Cin, xor_out => 
                           xor_b_27_port);
   bc_xor_26 : my_xor_155 port map( A => B(26), B => Cin, xor_out => 
                           xor_b_26_port);
   bc_xor_25 : my_xor_154 port map( A => B(25), B => Cin, xor_out => 
                           xor_b_25_port);
   bc_xor_24 : my_xor_153 port map( A => B(24), B => Cin, xor_out => 
                           xor_b_24_port);
   bc_xor_23 : my_xor_152 port map( A => B(23), B => Cin, xor_out => 
                           xor_b_23_port);
   bc_xor_22 : my_xor_151 port map( A => B(22), B => Cin, xor_out => 
                           xor_b_22_port);
   bc_xor_21 : my_xor_150 port map( A => B(21), B => Cin, xor_out => 
                           xor_b_21_port);
   bc_xor_20 : my_xor_149 port map( A => B(20), B => Cin, xor_out => 
                           xor_b_20_port);
   bc_xor_19 : my_xor_148 port map( A => B(19), B => Cin, xor_out => 
                           xor_b_19_port);
   bc_xor_18 : my_xor_147 port map( A => B(18), B => Cin, xor_out => 
                           xor_b_18_port);
   bc_xor_17 : my_xor_146 port map( A => B(17), B => Cin, xor_out => 
                           xor_b_17_port);
   bc_xor_16 : my_xor_145 port map( A => B(16), B => Cin, xor_out => 
                           xor_b_16_port);
   bc_xor_15 : my_xor_144 port map( A => B(15), B => Cin, xor_out => 
                           xor_b_15_port);
   bc_xor_14 : my_xor_143 port map( A => B(14), B => Cin, xor_out => 
                           xor_b_14_port);
   bc_xor_13 : my_xor_142 port map( A => B(13), B => Cin, xor_out => 
                           xor_b_13_port);
   bc_xor_12 : my_xor_141 port map( A => B(12), B => Cin, xor_out => 
                           xor_b_12_port);
   bc_xor_11 : my_xor_140 port map( A => B(11), B => Cin, xor_out => 
                           xor_b_11_port);
   bc_xor_10 : my_xor_139 port map( A => B(10), B => Cin, xor_out => 
                           xor_b_10_port);
   bc_xor_9 : my_xor_138 port map( A => B(9), B => Cin, xor_out => xor_b_9_port
                           );
   bc_xor_8 : my_xor_137 port map( A => B(8), B => Cin, xor_out => xor_b_8_port
                           );
   bc_xor_7 : my_xor_136 port map( A => B(7), B => Cin, xor_out => xor_b_7_port
                           );
   bc_xor_6 : my_xor_135 port map( A => B(6), B => Cin, xor_out => xor_b_6_port
                           );
   bc_xor_5 : my_xor_134 port map( A => B(5), B => Cin, xor_out => xor_b_5_port
                           );
   bc_xor_4 : my_xor_133 port map( A => B(4), B => Cin, xor_out => xor_b_4_port
                           );
   bc_xor_3 : my_xor_132 port map( A => B(3), B => Cin, xor_out => xor_b_3_port
                           );
   bc_xor_2 : my_xor_131 port map( A => B(2), B => Cin, xor_out => xor_b_2_port
                           );
   bc_xor_1 : my_xor_130 port map( A => B(1), B => Cin, xor_out => xor_b_1_port
                           );
   bc_xor_0 : my_xor_129 port map( A => B(0), B => Cin, xor_out => xor_b_0_port
                           );
   CG : CARRY_GENERATOR_NBIT64_NBIT_PER_BLOCK4_0 port map( A(63) => A(63), 
                           A(62) => A(62), A(61) => A(61), A(60) => A(60), 
                           A(59) => A(59), A(58) => A(58), A(57) => A(57), 
                           A(56) => A(56), A(55) => A(55), A(54) => A(54), 
                           A(53) => A(53), A(52) => A(52), A(51) => A(51), 
                           A(50) => A(50), A(49) => A(49), A(48) => A(48), 
                           A(47) => A(47), A(46) => A(46), A(45) => A(45), 
                           A(44) => A(44), A(43) => A(43), A(42) => A(42), 
                           A(41) => A(41), A(40) => A(40), A(39) => A(39), 
                           A(38) => A(38), A(37) => A(37), A(36) => A(36), 
                           A(35) => A(35), A(34) => A(34), A(33) => A(33), 
                           A(32) => A(32), A(31) => A(31), A(30) => A(30), 
                           A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(63) => xor_b_63_port, B(62) =>
                           xor_b_62_port, B(61) => xor_b_61_port, B(60) => 
                           xor_b_60_port, B(59) => xor_b_59_port, B(58) => 
                           xor_b_58_port, B(57) => xor_b_57_port, B(56) => 
                           xor_b_56_port, B(55) => xor_b_55_port, B(54) => 
                           xor_b_54_port, B(53) => xor_b_53_port, B(52) => 
                           xor_b_52_port, B(51) => xor_b_51_port, B(50) => 
                           xor_b_50_port, B(49) => xor_b_49_port, B(48) => 
                           xor_b_48_port, B(47) => xor_b_47_port, B(46) => 
                           xor_b_46_port, B(45) => xor_b_45_port, B(44) => 
                           xor_b_44_port, B(43) => xor_b_43_port, B(42) => 
                           xor_b_42_port, B(41) => xor_b_41_port, B(40) => 
                           xor_b_40_port, B(39) => xor_b_39_port, B(38) => 
                           xor_b_38_port, B(37) => xor_b_37_port, B(36) => 
                           xor_b_36_port, B(35) => xor_b_35_port, B(34) => 
                           xor_b_34_port, B(33) => xor_b_33_port, B(32) => 
                           xor_b_32_port, B(31) => xor_b_31_port, B(30) => 
                           xor_b_30_port, B(29) => xor_b_29_port, B(28) => 
                           xor_b_28_port, B(27) => xor_b_27_port, B(26) => 
                           xor_b_26_port, B(25) => xor_b_25_port, B(24) => 
                           xor_b_24_port, B(23) => xor_b_23_port, B(22) => 
                           xor_b_22_port, B(21) => xor_b_21_port, B(20) => 
                           xor_b_20_port, B(19) => xor_b_19_port, B(18) => 
                           xor_b_18_port, B(17) => xor_b_17_port, B(16) => 
                           xor_b_16_port, B(15) => xor_b_15_port, B(14) => 
                           xor_b_14_port, B(13) => xor_b_13_port, B(12) => 
                           xor_b_12_port, B(11) => xor_b_11_port, B(10) => 
                           xor_b_10_port, B(9) => xor_b_9_port, B(8) => 
                           xor_b_8_port, B(7) => xor_b_7_port, B(6) => 
                           xor_b_6_port, B(5) => xor_b_5_port, B(4) => 
                           xor_b_4_port, B(3) => xor_b_3_port, B(2) => 
                           xor_b_2_port, B(1) => xor_b_1_port, B(0) => 
                           xor_b_0_port, Cin => Cin, Co(15) => Cout, Co(14) => 
                           carry_14_port, Co(13) => carry_13_port, Co(12) => 
                           carry_12_port, Co(11) => carry_11_port, Co(10) => 
                           carry_10_port, Co(9) => carry_9_port, Co(8) => 
                           carry_8_port, Co(7) => carry_7_port, Co(6) => 
                           carry_6_port, Co(5) => carry_5_port, Co(4) => 
                           carry_4_port, Co(3) => carry_3_port, Co(2) => 
                           carry_2_port, Co(1) => carry_1_port, Co(0) => 
                           carry_0_port);
   SG : sum_generator_n_bit64_n_CSB16_0 port map( A(63) => A(63), A(62) => 
                           A(62), A(61) => A(61), A(60) => A(60), A(59) => 
                           A(59), A(58) => A(58), A(57) => A(57), A(56) => 
                           A(56), A(55) => A(55), A(54) => A(54), A(53) => 
                           A(53), A(52) => A(52), A(51) => A(51), A(50) => 
                           A(50), A(49) => A(49), A(48) => A(48), A(47) => 
                           A(47), A(46) => A(46), A(45) => A(45), A(44) => 
                           A(44), A(43) => A(43), A(42) => A(42), A(41) => 
                           A(41), A(40) => A(40), A(39) => A(39), A(38) => 
                           A(38), A(37) => A(37), A(36) => A(36), A(35) => 
                           A(35), A(34) => A(34), A(33) => A(33), A(32) => 
                           A(32), A(31) => A(31), A(30) => A(30), A(29) => 
                           A(29), A(28) => A(28), A(27) => A(27), A(26) => 
                           A(26), A(25) => A(25), A(24) => A(24), A(23) => 
                           A(23), A(22) => A(22), A(21) => A(21), A(20) => 
                           A(20), A(19) => A(19), A(18) => A(18), A(17) => 
                           A(17), A(16) => A(16), A(15) => A(15), A(14) => 
                           A(14), A(13) => A(13), A(12) => A(12), A(11) => 
                           A(11), A(10) => A(10), A(9) => A(9), A(8) => A(8), 
                           A(7) => A(7), A(6) => A(6), A(5) => A(5), A(4) => 
                           A(4), A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), B(63) => xor_b_63_port, B(62) => 
                           xor_b_62_port, B(61) => xor_b_61_port, B(60) => 
                           xor_b_60_port, B(59) => xor_b_59_port, B(58) => 
                           xor_b_58_port, B(57) => xor_b_57_port, B(56) => 
                           xor_b_56_port, B(55) => xor_b_55_port, B(54) => 
                           xor_b_54_port, B(53) => xor_b_53_port, B(52) => 
                           xor_b_52_port, B(51) => xor_b_51_port, B(50) => 
                           xor_b_50_port, B(49) => xor_b_49_port, B(48) => 
                           xor_b_48_port, B(47) => xor_b_47_port, B(46) => 
                           xor_b_46_port, B(45) => xor_b_45_port, B(44) => 
                           xor_b_44_port, B(43) => xor_b_43_port, B(42) => 
                           xor_b_42_port, B(41) => xor_b_41_port, B(40) => 
                           xor_b_40_port, B(39) => xor_b_39_port, B(38) => 
                           xor_b_38_port, B(37) => xor_b_37_port, B(36) => 
                           xor_b_36_port, B(35) => xor_b_35_port, B(34) => 
                           xor_b_34_port, B(33) => xor_b_33_port, B(32) => 
                           xor_b_32_port, B(31) => xor_b_31_port, B(30) => 
                           xor_b_30_port, B(29) => xor_b_29_port, B(28) => 
                           xor_b_28_port, B(27) => xor_b_27_port, B(26) => 
                           xor_b_26_port, B(25) => xor_b_25_port, B(24) => 
                           xor_b_24_port, B(23) => xor_b_23_port, B(22) => 
                           xor_b_22_port, B(21) => xor_b_21_port, B(20) => 
                           xor_b_20_port, B(19) => xor_b_19_port, B(18) => 
                           xor_b_18_port, B(17) => xor_b_17_port, B(16) => 
                           xor_b_16_port, B(15) => xor_b_15_port, B(14) => 
                           xor_b_14_port, B(13) => xor_b_13_port, B(12) => 
                           xor_b_12_port, B(11) => xor_b_11_port, B(10) => 
                           xor_b_10_port, B(9) => xor_b_9_port, B(8) => 
                           xor_b_8_port, B(7) => xor_b_7_port, B(6) => 
                           xor_b_6_port, B(5) => xor_b_5_port, B(4) => 
                           xor_b_4_port, B(3) => xor_b_3_port, B(2) => 
                           xor_b_2_port, B(1) => xor_b_1_port, B(0) => 
                           xor_b_0_port, C_in(15) => carry_14_port, C_in(14) =>
                           carry_13_port, C_in(13) => carry_12_port, C_in(12) 
                           => carry_11_port, C_in(11) => carry_10_port, 
                           C_in(10) => carry_9_port, C_in(9) => carry_8_port, 
                           C_in(8) => carry_7_port, C_in(7) => carry_6_port, 
                           C_in(6) => carry_5_port, C_in(5) => carry_4_port, 
                           C_in(4) => carry_3_port, C_in(3) => carry_2_port, 
                           C_in(2) => carry_1_port, C_in(1) => carry_0_port, 
                           C_in(0) => Cin, S(63) => S_63_port, S(62) => 
                           S_62_port, S(61) => S_61_port, S(60) => S_60_port, 
                           S(59) => S_59_port, S(58) => S_58_port, S(57) => 
                           S_57_port, S(56) => S_56_port, S(55) => S_55_port, 
                           S(54) => S_54_port, S(53) => S_53_port, S(52) => 
                           S_52_port, S(51) => S_51_port, S(50) => S_50_port, 
                           S(49) => S_49_port, S(48) => S_48_port, S(47) => 
                           S_47_port, S(46) => S_46_port, S(45) => S_45_port, 
                           S(44) => S_44_port, S(43) => S_43_port, S(42) => 
                           S_42_port, S(41) => S_41_port, S(40) => S_40_port, 
                           S(39) => S_39_port, S(38) => S_38_port, S(37) => 
                           S_37_port, S(36) => S_36_port, S(35) => S_35_port, 
                           S(34) => S_34_port, S(33) => S_33_port, S(32) => 
                           S_32_port, S(31) => S_31_port, S(30) => S_30_port, 
                           S(29) => S_29_port, S(28) => S_28_port, S(27) => 
                           S_27_port, S(26) => S_26_port, S(25) => S_25_port, 
                           S(24) => S_24_port, S(23) => S_23_port, S(22) => 
                           S_22_port, S(21) => S_21_port, S(20) => S_20_port, 
                           S(19) => S_19_port, S(18) => S_18_port, S(17) => 
                           S_17_port, S(16) => S_16_port, S(15) => S_15_port, 
                           S(14) => S_14_port, S(13) => S_13_port, S(12) => 
                           S_12_port, S(11) => S_11_port, S(10) => S_10_port, 
                           S(9) => S_9_port, S(8) => S_8_port, S(7) => S_7_port
                           , S(6) => S_6_port, S(5) => S_5_port, S(4) => 
                           S_4_port, S(3) => S_3_port, S(2) => S_2_port, S(1) 
                           => S_1_port, S(0) => S_0_port);
   U1 : XNOR2_X1 port map( A => A(63), B => S_63_port, ZN => n1);
   U2 : NOR2_X1 port map( A1 => n1, A2 => n2, ZN => ovf);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity mux51_gen_NBIT32_0 is

   port( A0, A1, A2, A3, A4 : in std_logic_vector (31 downto 0);  SEL : in 
         std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end mux51_gen_NBIT32_0;

architecture SYN_data_fl of mux51_gen_NBIT32_0 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, 
      n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32
      , n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, 
      n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61
      , n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n1, n2, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86 : std_logic;

begin
   
   U2 : BUF_X1 port map( A => n8, Z => n73);
   U3 : BUF_X1 port map( A => n8, Z => n74);
   U4 : BUF_X1 port map( A => n9, Z => n1);
   U5 : BUF_X1 port map( A => n5, Z => n82);
   U6 : BUF_X1 port map( A => n5, Z => n83);
   U7 : BUF_X1 port map( A => n5, Z => n84);
   U8 : BUF_X1 port map( A => n6, Z => n79);
   U9 : BUF_X1 port map( A => n6, Z => n80);
   U10 : BUF_X1 port map( A => n7, Z => n76);
   U11 : BUF_X1 port map( A => n7, Z => n77);
   U12 : BUF_X1 port map( A => n8, Z => n75);
   U13 : BUF_X1 port map( A => n6, Z => n81);
   U14 : BUF_X1 port map( A => n7, Z => n78);
   U15 : INV_X1 port map( A => SEL(1), ZN => n85);
   U16 : BUF_X1 port map( A => n9, Z => n2);
   U17 : BUF_X1 port map( A => n9, Z => n72);
   U18 : NOR3_X1 port map( A1 => SEL(0), A2 => SEL(2), A3 => n85, ZN => n5);
   U19 : NOR3_X1 port map( A1 => SEL(0), A2 => SEL(1), A3 => n1, ZN => n8);
   U20 : NOR3_X1 port map( A1 => SEL(1), A2 => SEL(2), A3 => SEL(0), ZN => n9);
   U21 : AND3_X1 port map( A1 => SEL(0), A2 => n86, A3 => SEL(1), ZN => n7);
   U22 : AND3_X1 port map( A1 => n85, A2 => n86, A3 => SEL(0), ZN => n6);
   U23 : INV_X1 port map( A => SEL(2), ZN => n86);
   U24 : NAND2_X1 port map( A1 => n28, A2 => n29, ZN => Y(29));
   U25 : AOI22_X1 port map( A1 => A4(29), A2 => n74, B1 => A0(29), B2 => n2, ZN
                           => n28);
   U26 : AOI222_X1 port map( A1 => A2(29), A2 => n83, B1 => A1(29), B2 => n80, 
                           C1 => A3(29), C2 => n77, ZN => n29);
   U27 : NAND2_X1 port map( A1 => n24, A2 => n25, ZN => Y(30));
   U28 : AOI22_X1 port map( A1 => A4(30), A2 => n74, B1 => A0(30), B2 => n72, 
                           ZN => n24);
   U29 : AOI222_X1 port map( A1 => A2(30), A2 => n84, B1 => A1(30), B2 => n80, 
                           C1 => A3(30), C2 => n77, ZN => n25);
   U30 : NAND2_X1 port map( A1 => n36, A2 => n37, ZN => Y(25));
   U31 : AOI22_X1 port map( A1 => A4(25), A2 => n74, B1 => A0(25), B2 => n2, ZN
                           => n36);
   U32 : AOI222_X1 port map( A1 => A2(25), A2 => n83, B1 => A1(25), B2 => n80, 
                           C1 => A3(25), C2 => n77, ZN => n37);
   U33 : NAND2_X1 port map( A1 => n34, A2 => n35, ZN => Y(26));
   U34 : AOI22_X1 port map( A1 => A4(26), A2 => n74, B1 => A0(26), B2 => n2, ZN
                           => n34);
   U35 : AOI222_X1 port map( A1 => A2(26), A2 => n83, B1 => A1(26), B2 => n80, 
                           C1 => A3(26), C2 => n77, ZN => n35);
   U36 : NAND2_X1 port map( A1 => n32, A2 => n33, ZN => Y(27));
   U37 : AOI22_X1 port map( A1 => A4(27), A2 => n74, B1 => A0(27), B2 => n2, ZN
                           => n32);
   U38 : AOI222_X1 port map( A1 => A2(27), A2 => n83, B1 => A1(27), B2 => n80, 
                           C1 => A3(27), C2 => n77, ZN => n33);
   U39 : NAND2_X1 port map( A1 => n30, A2 => n31, ZN => Y(28));
   U40 : AOI22_X1 port map( A1 => A4(28), A2 => n74, B1 => A0(28), B2 => n2, ZN
                           => n30);
   U41 : AOI222_X1 port map( A1 => A2(28), A2 => n83, B1 => A1(28), B2 => n80, 
                           C1 => A3(28), C2 => n77, ZN => n31);
   U42 : NAND2_X1 port map( A1 => n40, A2 => n41, ZN => Y(23));
   U43 : AOI22_X1 port map( A1 => A4(23), A2 => n74, B1 => A0(23), B2 => n2, ZN
                           => n40);
   U44 : AOI222_X1 port map( A1 => A2(23), A2 => n83, B1 => A1(23), B2 => n80, 
                           C1 => A3(23), C2 => n77, ZN => n41);
   U45 : NAND2_X1 port map( A1 => n38, A2 => n39, ZN => Y(24));
   U46 : AOI22_X1 port map( A1 => A4(24), A2 => n74, B1 => A0(24), B2 => n2, ZN
                           => n38);
   U47 : AOI222_X1 port map( A1 => A2(24), A2 => n83, B1 => A1(24), B2 => n80, 
                           C1 => A3(24), C2 => n77, ZN => n39);
   U48 : NAND2_X1 port map( A1 => n22, A2 => n23, ZN => Y(31));
   U49 : AOI22_X1 port map( A1 => A4(31), A2 => n75, B1 => A0(31), B2 => n72, 
                           ZN => n22);
   U50 : AOI222_X1 port map( A1 => A2(31), A2 => n84, B1 => A1(31), B2 => n81, 
                           C1 => A3(31), C2 => n78, ZN => n23);
   U51 : NAND2_X1 port map( A1 => n64, A2 => n65, ZN => Y(12));
   U52 : AOI22_X1 port map( A1 => A4(12), A2 => n73, B1 => A0(12), B2 => n1, ZN
                           => n64);
   U53 : AOI222_X1 port map( A1 => A2(12), A2 => n82, B1 => A1(12), B2 => n79, 
                           C1 => A3(12), C2 => n76, ZN => n65);
   U54 : NAND2_X1 port map( A1 => n62, A2 => n63, ZN => Y(13));
   U55 : AOI22_X1 port map( A1 => A4(13), A2 => n73, B1 => A0(13), B2 => n1, ZN
                           => n62);
   U56 : AOI222_X1 port map( A1 => A2(13), A2 => n82, B1 => A1(13), B2 => n79, 
                           C1 => A3(13), C2 => n76, ZN => n63);
   U57 : NAND2_X1 port map( A1 => n60, A2 => n61, ZN => Y(14));
   U58 : AOI22_X1 port map( A1 => A4(14), A2 => n73, B1 => A0(14), B2 => n1, ZN
                           => n60);
   U59 : AOI222_X1 port map( A1 => A2(14), A2 => n82, B1 => A1(14), B2 => n79, 
                           C1 => A3(14), C2 => n76, ZN => n61);
   U60 : NAND2_X1 port map( A1 => n58, A2 => n59, ZN => Y(15));
   U61 : AOI22_X1 port map( A1 => A4(15), A2 => n73, B1 => A0(15), B2 => n1, ZN
                           => n58);
   U62 : AOI222_X1 port map( A1 => A2(15), A2 => n82, B1 => A1(15), B2 => n79, 
                           C1 => A3(15), C2 => n76, ZN => n59);
   U63 : NAND2_X1 port map( A1 => n56, A2 => n57, ZN => Y(16));
   U64 : AOI22_X1 port map( A1 => A4(16), A2 => n73, B1 => A0(16), B2 => n1, ZN
                           => n56);
   U65 : AOI222_X1 port map( A1 => A2(16), A2 => n82, B1 => A1(16), B2 => n79, 
                           C1 => A3(16), C2 => n76, ZN => n57);
   U66 : NAND2_X1 port map( A1 => n54, A2 => n55, ZN => Y(17));
   U67 : AOI22_X1 port map( A1 => A4(17), A2 => n73, B1 => A0(17), B2 => n1, ZN
                           => n54);
   U68 : AOI222_X1 port map( A1 => A2(17), A2 => n82, B1 => A1(17), B2 => n79, 
                           C1 => A3(17), C2 => n76, ZN => n55);
   U69 : NAND2_X1 port map( A1 => n52, A2 => n53, ZN => Y(18));
   U70 : AOI22_X1 port map( A1 => A4(18), A2 => n73, B1 => A0(18), B2 => n1, ZN
                           => n52);
   U71 : AOI222_X1 port map( A1 => A2(18), A2 => n82, B1 => A1(18), B2 => n79, 
                           C1 => A3(18), C2 => n76, ZN => n53);
   U72 : NAND2_X1 port map( A1 => n50, A2 => n51, ZN => Y(19));
   U73 : AOI22_X1 port map( A1 => A4(19), A2 => n73, B1 => A0(19), B2 => n1, ZN
                           => n50);
   U74 : AOI222_X1 port map( A1 => A2(19), A2 => n82, B1 => A1(19), B2 => n79, 
                           C1 => A3(19), C2 => n76, ZN => n51);
   U75 : NAND2_X1 port map( A1 => n46, A2 => n47, ZN => Y(20));
   U76 : AOI22_X1 port map( A1 => A4(20), A2 => n74, B1 => A0(20), B2 => n2, ZN
                           => n46);
   U77 : AOI222_X1 port map( A1 => A2(20), A2 => n83, B1 => A1(20), B2 => n80, 
                           C1 => A3(20), C2 => n77, ZN => n47);
   U78 : NAND2_X1 port map( A1 => n44, A2 => n45, ZN => Y(21));
   U79 : AOI22_X1 port map( A1 => A4(21), A2 => n74, B1 => A0(21), B2 => n2, ZN
                           => n44);
   U80 : AOI222_X1 port map( A1 => A2(21), A2 => n83, B1 => A1(21), B2 => n80, 
                           C1 => A3(21), C2 => n77, ZN => n45);
   U81 : NAND2_X1 port map( A1 => n42, A2 => n43, ZN => Y(22));
   U82 : AOI22_X1 port map( A1 => A4(22), A2 => n74, B1 => A0(22), B2 => n2, ZN
                           => n42);
   U83 : AOI222_X1 port map( A1 => A2(22), A2 => n83, B1 => A1(22), B2 => n80, 
                           C1 => A3(22), C2 => n77, ZN => n43);
   U84 : NAND2_X1 port map( A1 => n10, A2 => n11, ZN => Y(8));
   U85 : AOI22_X1 port map( A1 => A4(8), A2 => n75, B1 => A0(8), B2 => n72, ZN 
                           => n10);
   U86 : AOI222_X1 port map( A1 => A2(8), A2 => n84, B1 => A1(8), B2 => n81, C1
                           => A3(8), C2 => n78, ZN => n11);
   U87 : NAND2_X1 port map( A1 => n3, A2 => n4, ZN => Y(9));
   U88 : AOI22_X1 port map( A1 => A4(9), A2 => n75, B1 => A0(9), B2 => n72, ZN 
                           => n3);
   U89 : AOI222_X1 port map( A1 => A2(9), A2 => n84, B1 => A1(9), B2 => n81, C1
                           => A3(9), C2 => n78, ZN => n4);
   U90 : NAND2_X1 port map( A1 => n68, A2 => n69, ZN => Y(10));
   U91 : AOI22_X1 port map( A1 => A4(10), A2 => n73, B1 => A0(10), B2 => n1, ZN
                           => n68);
   U92 : AOI222_X1 port map( A1 => A2(10), A2 => n82, B1 => A1(10), B2 => n79, 
                           C1 => A3(10), C2 => n76, ZN => n69);
   U93 : NAND2_X1 port map( A1 => n66, A2 => n67, ZN => Y(11));
   U94 : AOI22_X1 port map( A1 => A4(11), A2 => n73, B1 => A0(11), B2 => n1, ZN
                           => n66);
   U95 : AOI222_X1 port map( A1 => A2(11), A2 => n82, B1 => A1(11), B2 => n79, 
                           C1 => A3(11), C2 => n76, ZN => n67);
   U96 : NAND2_X1 port map( A1 => n48, A2 => n49, ZN => Y(1));
   U97 : AOI222_X1 port map( A1 => A2(1), A2 => n83, B1 => A1(1), B2 => n79, C1
                           => A3(1), C2 => n76, ZN => n49);
   U98 : AOI22_X1 port map( A1 => A4(1), A2 => n73, B1 => A0(1), B2 => n2, ZN 
                           => n48);
   U99 : NAND2_X1 port map( A1 => n26, A2 => n27, ZN => Y(2));
   U100 : AOI222_X1 port map( A1 => A2(2), A2 => n84, B1 => A1(2), B2 => n80, 
                           C1 => A3(2), C2 => n77, ZN => n27);
   U101 : AOI22_X1 port map( A1 => A4(2), A2 => n74, B1 => A0(2), B2 => n2, ZN 
                           => n26);
   U102 : NAND2_X1 port map( A1 => n20, A2 => n21, ZN => Y(3));
   U103 : AOI222_X1 port map( A1 => A2(3), A2 => n84, B1 => A1(3), B2 => n81, 
                           C1 => A3(3), C2 => n78, ZN => n21);
   U104 : AOI22_X1 port map( A1 => A4(3), A2 => n75, B1 => A0(3), B2 => n72, ZN
                           => n20);
   U105 : NAND2_X1 port map( A1 => n18, A2 => n19, ZN => Y(4));
   U106 : AOI222_X1 port map( A1 => A2(4), A2 => n84, B1 => A1(4), B2 => n81, 
                           C1 => A3(4), C2 => n78, ZN => n19);
   U107 : AOI22_X1 port map( A1 => A4(4), A2 => n75, B1 => A0(4), B2 => n72, ZN
                           => n18);
   U108 : NAND2_X1 port map( A1 => n16, A2 => n17, ZN => Y(5));
   U109 : AOI22_X1 port map( A1 => A4(5), A2 => n75, B1 => A0(5), B2 => n72, ZN
                           => n16);
   U110 : AOI222_X1 port map( A1 => A2(5), A2 => n84, B1 => A1(5), B2 => n81, 
                           C1 => A3(5), C2 => n78, ZN => n17);
   U111 : NAND2_X1 port map( A1 => n14, A2 => n15, ZN => Y(6));
   U112 : AOI22_X1 port map( A1 => A4(6), A2 => n75, B1 => A0(6), B2 => n72, ZN
                           => n14);
   U113 : AOI222_X1 port map( A1 => A2(6), A2 => n84, B1 => A1(6), B2 => n81, 
                           C1 => A3(6), C2 => n78, ZN => n15);
   U114 : NAND2_X1 port map( A1 => n12, A2 => n13, ZN => Y(7));
   U115 : AOI22_X1 port map( A1 => A4(7), A2 => n75, B1 => A0(7), B2 => n72, ZN
                           => n12);
   U116 : AOI222_X1 port map( A1 => A2(7), A2 => n84, B1 => A1(7), B2 => n81, 
                           C1 => A3(7), C2 => n78, ZN => n13);
   U117 : NAND2_X1 port map( A1 => n70, A2 => n71, ZN => Y(0));
   U118 : AOI22_X1 port map( A1 => A4(0), A2 => n73, B1 => A0(0), B2 => n1, ZN 
                           => n70);
   U119 : AOI222_X1 port map( A1 => A2(0), A2 => n82, B1 => A1(0), B2 => n79, 
                           C1 => A3(0), C2 => n76, ZN => n71);

end SYN_data_fl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity negate_NBIT32_0 is

   port( A : in std_logic_vector (31 downto 0);  Y : out std_logic_vector (31 
         downto 0));

end negate_NBIT32_0;

architecture SYN_data_fl of negate_NBIT32_0 is

   component negate_NBIT32_0_DW01_sub_0
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  DIFF
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   signal n1, n2, n_1572 : std_logic;

begin
   
   n1 <= '0';
   n2 <= '0';
   sub_add_14_b0 : negate_NBIT32_0_DW01_sub_0 port map( A(31) => n1, A(30) => 
                           n1, A(29) => n1, A(28) => n1, A(27) => n1, A(26) => 
                           n1, A(25) => n1, A(24) => n1, A(23) => n1, A(22) => 
                           n1, A(21) => n1, A(20) => n1, A(19) => n1, A(18) => 
                           n1, A(17) => n1, A(16) => n1, A(15) => n1, A(14) => 
                           n1, A(13) => n1, A(12) => n1, A(11) => n1, A(10) => 
                           n1, A(9) => n1, A(8) => n1, A(7) => n1, A(6) => n1, 
                           A(5) => n1, A(4) => n1, A(3) => n1, A(2) => n1, A(1)
                           => n1, A(0) => n1, B(31) => A(31), B(30) => A(30), 
                           B(29) => A(29), B(28) => A(28), B(27) => A(27), 
                           B(26) => A(26), B(25) => A(25), B(24) => A(24), 
                           B(23) => A(23), B(22) => A(22), B(21) => A(21), 
                           B(20) => A(20), B(19) => A(19), B(18) => A(18), 
                           B(17) => A(17), B(16) => A(16), B(15) => A(15), 
                           B(14) => A(14), B(13) => A(13), B(12) => A(12), 
                           B(11) => A(11), B(10) => A(10), B(9) => A(9), B(8) 
                           => A(8), B(7) => A(7), B(6) => A(6), B(5) => A(5), 
                           B(4) => A(4), B(3) => A(3), B(2) => A(2), B(1) => 
                           A(1), B(0) => A(0), CI => n2, DIFF(31) => Y(31), 
                           DIFF(30) => Y(30), DIFF(29) => Y(29), DIFF(28) => 
                           Y(28), DIFF(27) => Y(27), DIFF(26) => Y(26), 
                           DIFF(25) => Y(25), DIFF(24) => Y(24), DIFF(23) => 
                           Y(23), DIFF(22) => Y(22), DIFF(21) => Y(21), 
                           DIFF(20) => Y(20), DIFF(19) => Y(19), DIFF(18) => 
                           Y(18), DIFF(17) => Y(17), DIFF(16) => Y(16), 
                           DIFF(15) => Y(15), DIFF(14) => Y(14), DIFF(13) => 
                           Y(13), DIFF(12) => Y(12), DIFF(11) => Y(11), 
                           DIFF(10) => Y(10), DIFF(9) => Y(9), DIFF(8) => Y(8),
                           DIFF(7) => Y(7), DIFF(6) => Y(6), DIFF(5) => Y(5), 
                           DIFF(4) => Y(4), DIFF(3) => Y(3), DIFF(2) => Y(2), 
                           DIFF(1) => Y(1), DIFF(0) => Y(0), CO => n_1572);

end SYN_data_fl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity shl3_NBIT32 is

   port( A : in std_logic_vector (31 downto 0);  Y : out std_logic_vector (31 
         downto 0));

end shl3_NBIT32;

architecture SYN_behavioral of shl3_NBIT32 is

signal X_Logic0_port : std_logic;

begin
   Y <= ( A(28), A(27), A(26), A(25), A(24), A(23), A(22), A(21), A(20), A(19),
      A(18), A(17), A(16), A(15), A(14), A(13), A(12), A(11), A(10), A(9), A(8)
      , A(7), A(6), A(5), A(4), A(3), A(2), A(1), A(0), X_Logic0_port, 
      X_Logic0_port, X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity shl2_NBIT32_0 is

   port( A : in std_logic_vector (31 downto 0);  Y : out std_logic_vector (31 
         downto 0));

end shl2_NBIT32_0;

architecture SYN_behavioral of shl2_NBIT32_0 is

signal X_Logic0_port : std_logic;

begin
   Y <= ( A(29), A(28), A(27), A(26), A(25), A(24), A(23), A(22), A(21), A(20),
      A(19), A(18), A(17), A(16), A(15), A(14), A(13), A(12), A(11), A(10), 
      A(9), A(8), A(7), A(6), A(5), A(4), A(3), A(2), A(1), A(0), X_Logic0_port
      , X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity shl1_NBIT32_0 is

   port( A : in std_logic_vector (31 downto 0);  Y : out std_logic_vector (31 
         downto 0));

end shl1_NBIT32_0;

architecture SYN_datafl of shl1_NBIT32_0 is

signal X_Logic0_port : std_logic;

begin
   Y <= ( A(30), A(29), A(28), A(27), A(26), A(25), A(24), A(23), A(22), A(21),
      A(20), A(19), A(18), A(17), A(16), A(15), A(14), A(13), A(12), A(11), 
      A(10), A(9), A(8), A(7), A(6), A(5), A(4), A(3), A(2), A(1), A(0), 
      X_Logic0_port );
   
   X_Logic0_port <= '0';

end SYN_datafl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity enc33_0 is

   port( A : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (2 
         downto 0));

end enc33_0;

architecture SYN_behavioral of enc33_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n1, n2 : std_logic;

begin
   
   U8 : XOR2_X1 port map( A => A(0), B => A(1), Z => n4);
   U1 : OAI21_X1 port map( B1 => n2, B2 => n1, A => n5, ZN => Y(1));
   U2 : NOR3_X1 port map( A1 => n1, A2 => n3, A3 => n4, ZN => Y(2));
   U3 : OAI21_X1 port map( B1 => A(2), B2 => n2, A => n5, ZN => Y(0));
   U4 : INV_X1 port map( A => n4, ZN => n2);
   U5 : NAND2_X1 port map( A1 => n3, A2 => n1, ZN => n5);
   U6 : AND2_X1 port map( A1 => A(1), A2 => A(0), ZN => n3);
   U7 : INV_X1 port map( A => A(2), ZN => n1);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity comparator is

   port( Z, cout : in std_logic;  eq, neq, gt, lt, ge, le : out std_logic);

end comparator;

architecture SYN_Structural of comparator is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal le_port, neq_port : std_logic;

begin
   eq <= Z;
   neq <= neq_port;
   ge <= cout;
   le <= le_port;
   
   U1 : INV_X1 port map( A => le_port, ZN => gt);
   U2 : INV_X1 port map( A => cout, ZN => lt);
   U3 : NAND2_X1 port map( A1 => cout, A2 => neq_port, ZN => le_port);
   U4 : INV_X1 port map( A => Z, ZN => neq_port);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity nor_generic_NBITS32 is

   port( input : in std_logic_vector (31 downto 0);  result : out std_logic);

end nor_generic_NBITS32;

architecture SYN_Behavioral of nor_generic_NBITS32 is

   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10 : std_logic;

begin
   
   U1 : NOR4_X1 port map( A1 => input(1), A2 => input(19), A3 => input(18), A4 
                           => input(17), ZN => n5);
   U2 : NOR4_X1 port map( A1 => input(9), A2 => input(8), A3 => input(7), A4 =>
                           input(6), ZN => n10);
   U3 : NOR4_X1 port map( A1 => input(23), A2 => input(22), A3 => input(21), A4
                           => input(20), ZN => n6);
   U4 : NOR4_X1 port map( A1 => input(5), A2 => input(4), A3 => input(3), A4 =>
                           input(31), ZN => n9);
   U5 : NOR4_X1 port map( A1 => input(30), A2 => input(2), A3 => input(29), A4 
                           => input(28), ZN => n8);
   U6 : NOR4_X1 port map( A1 => input(16), A2 => input(15), A3 => input(14), A4
                           => input(13), ZN => n4);
   U7 : NOR4_X1 port map( A1 => input(27), A2 => input(26), A3 => input(25), A4
                           => input(24), ZN => n7);
   U8 : NOR2_X1 port map( A1 => n1, A2 => n2, ZN => result);
   U9 : NAND4_X1 port map( A1 => n3, A2 => n4, A3 => n5, A4 => n6, ZN => n2);
   U10 : NAND4_X1 port map( A1 => n7, A2 => n8, A3 => n9, A4 => n10, ZN => n1);
   U11 : NOR4_X1 port map( A1 => input(12), A2 => input(11), A3 => input(10), 
                           A4 => input(0), ZN => n3);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity logicals_nbit32 is

   port( func : in std_logic_vector (3 downto 0);  SN : in std_logic;  in1, in2
         : in std_logic_vector (31 downto 0);  o : out std_logic_vector (31 
         downto 0));

end logicals_nbit32;

architecture SYN_behavioral of logicals_nbit32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component nand41_1
      port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);
   end component;
   
   component nand41_2
      port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);
   end component;
   
   component nand41_3
      port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);
   end component;
   
   component nand41_4
      port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);
   end component;
   
   component nand41_5
      port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);
   end component;
   
   component nand41_6
      port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);
   end component;
   
   component nand41_7
      port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);
   end component;
   
   component nand41_8
      port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);
   end component;
   
   component nand41_9
      port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);
   end component;
   
   component nand41_10
      port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);
   end component;
   
   component nand41_11
      port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);
   end component;
   
   component nand41_12
      port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);
   end component;
   
   component nand41_13
      port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);
   end component;
   
   component nand41_14
      port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);
   end component;
   
   component nand41_15
      port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);
   end component;
   
   component nand41_16
      port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);
   end component;
   
   component nand41_17
      port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);
   end component;
   
   component nand41_18
      port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);
   end component;
   
   component nand41_19
      port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);
   end component;
   
   component nand41_20
      port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);
   end component;
   
   component nand41_21
      port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);
   end component;
   
   component nand41_22
      port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);
   end component;
   
   component nand41_23
      port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);
   end component;
   
   component nand41_24
      port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);
   end component;
   
   component nand41_25
      port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);
   end component;
   
   component nand41_26
      port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);
   end component;
   
   component nand41_27
      port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);
   end component;
   
   component nand41_28
      port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);
   end component;
   
   component nand41_29
      port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);
   end component;
   
   component nand41_30
      port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);
   end component;
   
   component nand41_31
      port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);
   end component;
   
   component nand41_0
      port( in1, in2, in3, in4 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_1
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_2
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_3
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_4
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_5
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_6
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_7
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_8
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_9
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_10
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_11
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_12
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_13
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_14
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_15
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_16
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_17
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_18
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_19
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_20
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_21
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_22
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_23
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_24
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_25
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_26
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_27
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_28
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_29
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_30
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_31
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_32
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_33
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_34
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_35
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_36
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_37
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_38
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_39
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_40
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_41
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_42
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_43
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_44
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_45
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_46
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_47
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_48
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_49
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_50
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_51
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_52
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_53
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_54
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_55
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_56
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_57
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_58
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_59
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_60
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_61
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_62
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_63
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_64
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_65
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_66
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_67
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_68
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_69
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_70
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_71
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_72
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_73
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_74
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_75
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_76
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_77
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_78
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_79
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_80
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_81
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_82
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_83
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_84
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_85
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_86
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_87
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_88
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_89
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_90
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_91
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_92
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_93
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_94
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_95
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_96
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_97
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_98
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_99
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_100
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_101
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_102
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_103
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_104
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_105
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_106
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_107
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_108
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_109
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_110
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_111
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_112
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_113
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_114
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_115
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_116
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_117
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_118
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_119
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_120
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_121
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_122
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_123
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_124
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_125
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_126
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_127
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component nand31_0
      port( in1, in2, in3 : in std_logic;  o : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal l0_31_port, l0_30_port, l0_29_port, l0_28_port, l0_27_port, 
      l0_26_port, l0_25_port, l0_24_port, l0_23_port, l0_22_port, l0_21_port, 
      l0_20_port, l0_19_port, l0_18_port, l0_17_port, l0_16_port, l0_15_port, 
      l0_14_port, l0_13_port, l0_12_port, l0_11_port, l0_10_port, l0_9_port, 
      l0_8_port, l0_7_port, l0_6_port, l0_5_port, l0_4_port, l0_3_port, 
      l0_2_port, l0_1_port, l0_0_port, s0_9_port, l1_31_port, l1_30_port, 
      l1_29_port, l1_28_port, l1_27_port, l1_26_port, l1_25_port, l1_24_port, 
      l1_23_port, l1_22_port, l1_21_port, l1_20_port, l1_19_port, l1_18_port, 
      l1_17_port, l1_16_port, l1_15_port, l1_14_port, l1_13_port, l1_12_port, 
      l1_11_port, l1_10_port, l1_9_port, l1_8_port, l1_7_port, l1_6_port, 
      l1_5_port, l1_4_port, l1_3_port, l1_2_port, l1_1_port, l1_0_port, 
      l2_31_port, l2_30_port, l2_29_port, l2_28_port, l2_27_port, l2_26_port, 
      l2_25_port, l2_24_port, l2_23_port, l2_22_port, l2_21_port, l2_20_port, 
      l2_19_port, l2_18_port, l2_17_port, l2_16_port, l2_15_port, l2_14_port, 
      l2_13_port, l2_12_port, l2_11_port, l2_10_port, l2_9_port, l2_8_port, 
      l2_7_port, l2_6_port, l2_5_port, l2_4_port, l2_3_port, l2_2_port, 
      l2_1_port, l2_0_port, s2_9_port, l3_31_port, l3_30_port, l3_29_port, 
      l3_28_port, l3_27_port, l3_26_port, l3_25_port, l3_24_port, l3_23_port, 
      l3_22_port, l3_21_port, l3_20_port, l3_19_port, l3_18_port, l3_17_port, 
      l3_16_port, l3_15_port, l3_14_port, l3_13_port, l3_12_port, l3_11_port, 
      l3_10_port, l3_9_port, l3_8_port, l3_7_port, l3_6_port, l3_5_port, 
      l3_4_port, l3_3_port, l3_2_port, l3_1_port, l3_0_port, s3_9_port, n69, 
      n70, n71, n72, n73, n74, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, 
      n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26
      , n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, 
      n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55
      , n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n75, 
      n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86 : std_logic;

begin
   
   U77 : NAND3_X1 port map( A1 => n69, A2 => n71, A3 => n72, ZN => s2_9_port);
   U78 : NAND3_X1 port map( A1 => n73, A2 => n86, A3 => func(0), ZN => n72);
   U79 : NAND3_X1 port map( A1 => n73, A2 => n21, A3 => SN, ZN => n71);
   g1_a_31 : nand31_0 port map( in1 => n12, in2 => n18, in3 => n85, o => 
                           l0_31_port);
   g1_b_31 : nand31_127 port map( in1 => n4, in2 => n18, in3 => in2(31), o => 
                           l1_31_port);
   g1_c_31 : nand31_126 port map( in1 => n4, in2 => in1(31), in3 => n85, o => 
                           l2_31_port);
   g1_d_31 : nand31_125 port map( in1 => n3, in2 => in1(31), in3 => in2(31), o 
                           => l3_31_port);
   g1_a_30 : nand31_124 port map( in1 => n10, in2 => n51, in3 => n84, o => 
                           l0_30_port);
   g1_b_30 : nand31_123 port map( in1 => n4, in2 => n51, in3 => in2(30), o => 
                           l1_30_port);
   g1_c_30 : nand31_122 port map( in1 => n4, in2 => in1(30), in3 => n84, o => 
                           l2_30_port);
   g1_d_30 : nand31_121 port map( in1 => n3, in2 => in1(30), in3 => in2(30), o 
                           => l3_30_port);
   g1_a_29 : nand31_120 port map( in1 => n10, in2 => n50, in3 => n83, o => 
                           l0_29_port);
   g1_b_29 : nand31_119 port map( in1 => n4, in2 => n50, in3 => in2(29), o => 
                           l1_29_port);
   g1_c_29 : nand31_118 port map( in1 => n4, in2 => in1(29), in3 => n83, o => 
                           l2_29_port);
   g1_d_29 : nand31_117 port map( in1 => n3, in2 => in1(29), in3 => in2(29), o 
                           => l3_29_port);
   g1_a_28 : nand31_116 port map( in1 => n10, in2 => n49, in3 => n82, o => 
                           l0_28_port);
   g1_b_28 : nand31_115 port map( in1 => n4, in2 => n49, in3 => in2(28), o => 
                           l1_28_port);
   g1_c_28 : nand31_114 port map( in1 => n4, in2 => in1(28), in3 => n82, o => 
                           l2_28_port);
   g1_d_28 : nand31_113 port map( in1 => n3, in2 => in1(28), in3 => in2(28), o 
                           => l3_28_port);
   g1_a_27 : nand31_112 port map( in1 => n10, in2 => n48, in3 => n81, o => 
                           l0_27_port);
   g1_b_27 : nand31_111 port map( in1 => n4, in2 => n48, in3 => in2(27), o => 
                           l1_27_port);
   g1_c_27 : nand31_110 port map( in1 => n4, in2 => in1(27), in3 => n81, o => 
                           l2_27_port);
   g1_d_27 : nand31_109 port map( in1 => n3, in2 => in1(27), in3 => in2(27), o 
                           => l3_27_port);
   g1_a_26 : nand31_108 port map( in1 => n10, in2 => n47, in3 => n80, o => 
                           l0_26_port);
   g1_b_26 : nand31_107 port map( in1 => n4, in2 => n47, in3 => in2(26), o => 
                           l1_26_port);
   g1_c_26 : nand31_106 port map( in1 => n5, in2 => in1(26), in3 => n80, o => 
                           l2_26_port);
   g1_d_26 : nand31_105 port map( in1 => n3, in2 => in1(26), in3 => in2(26), o 
                           => l3_26_port);
   g1_a_25 : nand31_104 port map( in1 => n10, in2 => n46, in3 => n79, o => 
                           l0_25_port);
   g1_b_25 : nand31_103 port map( in1 => n5, in2 => n46, in3 => in2(25), o => 
                           l1_25_port);
   g1_c_25 : nand31_102 port map( in1 => n5, in2 => in1(25), in3 => n79, o => 
                           l2_25_port);
   g1_d_25 : nand31_101 port map( in1 => n3, in2 => in1(25), in3 => in2(25), o 
                           => l3_25_port);
   g1_a_24 : nand31_100 port map( in1 => n10, in2 => n45, in3 => n78, o => 
                           l0_24_port);
   g1_b_24 : nand31_99 port map( in1 => n5, in2 => n45, in3 => in2(24), o => 
                           l1_24_port);
   g1_c_24 : nand31_98 port map( in1 => n5, in2 => in1(24), in3 => n78, o => 
                           l2_24_port);
   g1_d_24 : nand31_97 port map( in1 => n3, in2 => in1(24), in3 => in2(24), o 
                           => l3_24_port);
   g1_a_23 : nand31_96 port map( in1 => n10, in2 => n44, in3 => n77, o => 
                           l0_23_port);
   g1_b_23 : nand31_95 port map( in1 => n5, in2 => n44, in3 => in2(23), o => 
                           l1_23_port);
   g1_c_23 : nand31_94 port map( in1 => n5, in2 => in1(23), in3 => n77, o => 
                           l2_23_port);
   g1_d_23 : nand31_93 port map( in1 => n3, in2 => in1(23), in3 => in2(23), o 
                           => l3_23_port);
   g1_a_22 : nand31_92 port map( in1 => n10, in2 => n43, in3 => n76, o => 
                           l0_22_port);
   g1_b_22 : nand31_91 port map( in1 => n5, in2 => n43, in3 => in2(22), o => 
                           l1_22_port);
   g1_c_22 : nand31_90 port map( in1 => n5, in2 => in1(22), in3 => n76, o => 
                           l2_22_port);
   g1_d_22 : nand31_89 port map( in1 => n3, in2 => in1(22), in3 => in2(22), o 
                           => l3_22_port);
   g1_a_21 : nand31_88 port map( in1 => n10, in2 => n42, in3 => n75, o => 
                           l0_21_port);
   g1_b_21 : nand31_87 port map( in1 => n5, in2 => n42, in3 => in2(21), o => 
                           l1_21_port);
   g1_c_21 : nand31_86 port map( in1 => n5, in2 => in1(21), in3 => n75, o => 
                           l2_21_port);
   g1_d_21 : nand31_85 port map( in1 => n2, in2 => in1(21), in3 => in2(21), o 
                           => l3_21_port);
   g1_a_20 : nand31_84 port map( in1 => n10, in2 => n41, in3 => n68, o => 
                           l0_20_port);
   g1_b_20 : nand31_83 port map( in1 => n6, in2 => n41, in3 => in2(20), o => 
                           l1_20_port);
   g1_c_20 : nand31_82 port map( in1 => n6, in2 => in1(20), in3 => n68, o => 
                           l2_20_port);
   g1_d_20 : nand31_81 port map( in1 => n2, in2 => in1(20), in3 => in2(20), o 
                           => l3_20_port);
   g1_a_19 : nand31_80 port map( in1 => n11, in2 => n40, in3 => n67, o => 
                           l0_19_port);
   g1_b_19 : nand31_79 port map( in1 => n6, in2 => n40, in3 => in2(19), o => 
                           l1_19_port);
   g1_c_19 : nand31_78 port map( in1 => n6, in2 => in1(19), in3 => n67, o => 
                           l2_19_port);
   g1_d_19 : nand31_77 port map( in1 => n2, in2 => in1(19), in3 => in2(19), o 
                           => l3_19_port);
   g1_a_18 : nand31_76 port map( in1 => n11, in2 => n39, in3 => n66, o => 
                           l0_18_port);
   g1_b_18 : nand31_75 port map( in1 => n6, in2 => n39, in3 => in2(18), o => 
                           l1_18_port);
   g1_c_18 : nand31_74 port map( in1 => n6, in2 => in1(18), in3 => n66, o => 
                           l2_18_port);
   g1_d_18 : nand31_73 port map( in1 => n2, in2 => in1(18), in3 => in2(18), o 
                           => l3_18_port);
   g1_a_17 : nand31_72 port map( in1 => n11, in2 => n38, in3 => n65, o => 
                           l0_17_port);
   g1_b_17 : nand31_71 port map( in1 => n6, in2 => n38, in3 => in2(17), o => 
                           l1_17_port);
   g1_c_17 : nand31_70 port map( in1 => n6, in2 => in1(17), in3 => n65, o => 
                           l2_17_port);
   g1_d_17 : nand31_69 port map( in1 => n2, in2 => in1(17), in3 => in2(17), o 
                           => l3_17_port);
   g1_a_16 : nand31_68 port map( in1 => n11, in2 => n37, in3 => n64, o => 
                           l0_16_port);
   g1_b_16 : nand31_67 port map( in1 => n6, in2 => n37, in3 => in2(16), o => 
                           l1_16_port);
   g1_c_16 : nand31_66 port map( in1 => n6, in2 => in1(16), in3 => n64, o => 
                           l2_16_port);
   g1_d_16 : nand31_65 port map( in1 => n2, in2 => in1(16), in3 => in2(16), o 
                           => l3_16_port);
   g1_a_15 : nand31_64 port map( in1 => n11, in2 => n36, in3 => n63, o => 
                           l0_15_port);
   g1_b_15 : nand31_63 port map( in1 => n6, in2 => n36, in3 => in2(15), o => 
                           l1_15_port);
   g1_c_15 : nand31_62 port map( in1 => n7, in2 => in1(15), in3 => n63, o => 
                           l2_15_port);
   g1_d_15 : nand31_61 port map( in1 => n2, in2 => in1(15), in3 => in2(15), o 
                           => l3_15_port);
   g1_a_14 : nand31_60 port map( in1 => n11, in2 => n35, in3 => n62, o => 
                           l0_14_port);
   g1_b_14 : nand31_59 port map( in1 => n7, in2 => n35, in3 => in2(14), o => 
                           l1_14_port);
   g1_c_14 : nand31_58 port map( in1 => n7, in2 => in1(14), in3 => n62, o => 
                           l2_14_port);
   g1_d_14 : nand31_57 port map( in1 => n2, in2 => in1(14), in3 => in2(14), o 
                           => l3_14_port);
   g1_a_13 : nand31_56 port map( in1 => n11, in2 => n34, in3 => n61, o => 
                           l0_13_port);
   g1_b_13 : nand31_55 port map( in1 => n7, in2 => n34, in3 => in2(13), o => 
                           l1_13_port);
   g1_c_13 : nand31_54 port map( in1 => n7, in2 => in1(13), in3 => n61, o => 
                           l2_13_port);
   g1_d_13 : nand31_53 port map( in1 => n2, in2 => in1(13), in3 => in2(13), o 
                           => l3_13_port);
   g1_a_12 : nand31_52 port map( in1 => n11, in2 => n33, in3 => n60, o => 
                           l0_12_port);
   g1_b_12 : nand31_51 port map( in1 => n7, in2 => n33, in3 => in2(12), o => 
                           l1_12_port);
   g1_c_12 : nand31_50 port map( in1 => n7, in2 => in1(12), in3 => n60, o => 
                           l2_12_port);
   g1_d_12 : nand31_49 port map( in1 => n2, in2 => in1(12), in3 => in2(12), o 
                           => l3_12_port);
   g1_a_11 : nand31_48 port map( in1 => n11, in2 => n32, in3 => n59, o => 
                           l0_11_port);
   g1_b_11 : nand31_47 port map( in1 => n7, in2 => n32, in3 => in2(11), o => 
                           l1_11_port);
   g1_c_11 : nand31_46 port map( in1 => n7, in2 => in1(11), in3 => n59, o => 
                           l2_11_port);
   g1_d_11 : nand31_45 port map( in1 => n2, in2 => in1(11), in3 => in2(11), o 
                           => l3_11_port);
   g1_a_10 : nand31_44 port map( in1 => n11, in2 => n31, in3 => n58, o => 
                           l0_10_port);
   g1_b_10 : nand31_43 port map( in1 => n7, in2 => n31, in3 => in2(10), o => 
                           l1_10_port);
   g1_c_10 : nand31_42 port map( in1 => n7, in2 => in1(10), in3 => n58, o => 
                           l2_10_port);
   g1_d_10 : nand31_41 port map( in1 => n1, in2 => in1(10), in3 => in2(10), o 
                           => l3_10_port);
   g1_a_9 : nand31_40 port map( in1 => n11, in2 => n30, in3 => n57, o => 
                           l0_9_port);
   g1_b_9 : nand31_39 port map( in1 => n8, in2 => n30, in3 => in2(9), o => 
                           l1_9_port);
   g1_c_9 : nand31_38 port map( in1 => n8, in2 => in1(9), in3 => n57, o => 
                           l2_9_port);
   g1_d_9 : nand31_37 port map( in1 => n1, in2 => in1(9), in3 => in2(9), o => 
                           l3_9_port);
   g1_a_8 : nand31_36 port map( in1 => n12, in2 => n29, in3 => n56, o => 
                           l0_8_port);
   g1_b_8 : nand31_35 port map( in1 => n8, in2 => n29, in3 => in2(8), o => 
                           l1_8_port);
   g1_c_8 : nand31_34 port map( in1 => n8, in2 => in1(8), in3 => n56, o => 
                           l2_8_port);
   g1_d_8 : nand31_33 port map( in1 => n1, in2 => in1(8), in3 => in2(8), o => 
                           l3_8_port);
   g1_a_7 : nand31_32 port map( in1 => n12, in2 => n28, in3 => n55, o => 
                           l0_7_port);
   g1_b_7 : nand31_31 port map( in1 => n8, in2 => n28, in3 => in2(7), o => 
                           l1_7_port);
   g1_c_7 : nand31_30 port map( in1 => n8, in2 => in1(7), in3 => n55, o => 
                           l2_7_port);
   g1_d_7 : nand31_29 port map( in1 => n1, in2 => in1(7), in3 => in2(7), o => 
                           l3_7_port);
   g1_a_6 : nand31_28 port map( in1 => n12, in2 => n27, in3 => n54, o => 
                           l0_6_port);
   g1_b_6 : nand31_27 port map( in1 => n8, in2 => n27, in3 => in2(6), o => 
                           l1_6_port);
   g1_c_6 : nand31_26 port map( in1 => n8, in2 => in1(6), in3 => n54, o => 
                           l2_6_port);
   g1_d_6 : nand31_25 port map( in1 => n1, in2 => in1(6), in3 => in2(6), o => 
                           l3_6_port);
   g1_a_5 : nand31_24 port map( in1 => n12, in2 => n26, in3 => n53, o => 
                           l0_5_port);
   g1_b_5 : nand31_23 port map( in1 => n8, in2 => n26, in3 => in2(5), o => 
                           l1_5_port);
   g1_c_5 : nand31_22 port map( in1 => n8, in2 => in1(5), in3 => n53, o => 
                           l2_5_port);
   g1_d_5 : nand31_21 port map( in1 => n1, in2 => in1(5), in3 => in2(5), o => 
                           l3_5_port);
   g1_a_4 : nand31_20 port map( in1 => n12, in2 => n25, in3 => n17, o => 
                           l0_4_port);
   g1_b_4 : nand31_19 port map( in1 => n8, in2 => n25, in3 => in2(4), o => 
                           l1_4_port);
   g1_c_4 : nand31_18 port map( in1 => n9, in2 => in1(4), in3 => n17, o => 
                           l2_4_port);
   g1_d_4 : nand31_17 port map( in1 => n1, in2 => in1(4), in3 => in2(4), o => 
                           l3_4_port);
   g1_a_3 : nand31_16 port map( in1 => n12, in2 => n24, in3 => n16, o => 
                           l0_3_port);
   g1_b_3 : nand31_15 port map( in1 => n9, in2 => n24, in3 => in2(3), o => 
                           l1_3_port);
   g1_c_3 : nand31_14 port map( in1 => n9, in2 => in1(3), in3 => n16, o => 
                           l2_3_port);
   g1_d_3 : nand31_13 port map( in1 => n1, in2 => in1(3), in3 => in2(3), o => 
                           l3_3_port);
   g1_a_2 : nand31_12 port map( in1 => n12, in2 => n23, in3 => n15, o => 
                           l0_2_port);
   g1_b_2 : nand31_11 port map( in1 => n9, in2 => n23, in3 => in2(2), o => 
                           l1_2_port);
   g1_c_2 : nand31_10 port map( in1 => n9, in2 => in1(2), in3 => n15, o => 
                           l2_2_port);
   g1_d_2 : nand31_9 port map( in1 => n1, in2 => in1(2), in3 => in2(2), o => 
                           l3_2_port);
   g1_a_1 : nand31_8 port map( in1 => n12, in2 => n22, in3 => n14, o => 
                           l0_1_port);
   g1_b_1 : nand31_7 port map( in1 => n9, in2 => n22, in3 => in2(1), o => 
                           l1_1_port);
   g1_c_1 : nand31_6 port map( in1 => n9, in2 => in1(1), in3 => n14, o => 
                           l2_1_port);
   g1_d_1 : nand31_5 port map( in1 => n1, in2 => in1(1), in3 => in2(1), o => 
                           l3_1_port);
   g1_a_0 : nand31_4 port map( in1 => n12, in2 => n52, in3 => n13, o => 
                           l0_0_port);
   g1_b_0 : nand31_3 port map( in1 => n9, in2 => n52, in3 => in2(0), o => 
                           l1_0_port);
   g1_c_0 : nand31_2 port map( in1 => n9, in2 => in1(0), in3 => n13, o => 
                           l2_0_port);
   g1_d_0 : nand31_1 port map( in1 => n1, in2 => in1(0), in3 => in2(0), o => 
                           l3_0_port);
   g2_a_31 : nand41_0 port map( in1 => l0_31_port, in2 => l1_31_port, in3 => 
                           l2_31_port, in4 => l3_31_port, o => o(31));
   g2_a_30 : nand41_31 port map( in1 => l0_30_port, in2 => l1_30_port, in3 => 
                           l2_30_port, in4 => l3_30_port, o => o(30));
   g2_a_29 : nand41_30 port map( in1 => l0_29_port, in2 => l1_29_port, in3 => 
                           l2_29_port, in4 => l3_29_port, o => o(29));
   g2_a_28 : nand41_29 port map( in1 => l0_28_port, in2 => l1_28_port, in3 => 
                           l2_28_port, in4 => l3_28_port, o => o(28));
   g2_a_27 : nand41_28 port map( in1 => l0_27_port, in2 => l1_27_port, in3 => 
                           l2_27_port, in4 => l3_27_port, o => o(27));
   g2_a_26 : nand41_27 port map( in1 => l0_26_port, in2 => l1_26_port, in3 => 
                           l2_26_port, in4 => l3_26_port, o => o(26));
   g2_a_25 : nand41_26 port map( in1 => l0_25_port, in2 => l1_25_port, in3 => 
                           l2_25_port, in4 => l3_25_port, o => o(25));
   g2_a_24 : nand41_25 port map( in1 => l0_24_port, in2 => l1_24_port, in3 => 
                           l2_24_port, in4 => l3_24_port, o => o(24));
   g2_a_23 : nand41_24 port map( in1 => l0_23_port, in2 => l1_23_port, in3 => 
                           l2_23_port, in4 => l3_23_port, o => o(23));
   g2_a_22 : nand41_23 port map( in1 => l0_22_port, in2 => l1_22_port, in3 => 
                           l2_22_port, in4 => l3_22_port, o => o(22));
   g2_a_21 : nand41_22 port map( in1 => l0_21_port, in2 => l1_21_port, in3 => 
                           l2_21_port, in4 => l3_21_port, o => o(21));
   g2_a_20 : nand41_21 port map( in1 => l0_20_port, in2 => l1_20_port, in3 => 
                           l2_20_port, in4 => l3_20_port, o => o(20));
   g2_a_19 : nand41_20 port map( in1 => l0_19_port, in2 => l1_19_port, in3 => 
                           l2_19_port, in4 => l3_19_port, o => o(19));
   g2_a_18 : nand41_19 port map( in1 => l0_18_port, in2 => l1_18_port, in3 => 
                           l2_18_port, in4 => l3_18_port, o => o(18));
   g2_a_17 : nand41_18 port map( in1 => l0_17_port, in2 => l1_17_port, in3 => 
                           l2_17_port, in4 => l3_17_port, o => o(17));
   g2_a_16 : nand41_17 port map( in1 => l0_16_port, in2 => l1_16_port, in3 => 
                           l2_16_port, in4 => l3_16_port, o => o(16));
   g2_a_15 : nand41_16 port map( in1 => l0_15_port, in2 => l1_15_port, in3 => 
                           l2_15_port, in4 => l3_15_port, o => o(15));
   g2_a_14 : nand41_15 port map( in1 => l0_14_port, in2 => l1_14_port, in3 => 
                           l2_14_port, in4 => l3_14_port, o => o(14));
   g2_a_13 : nand41_14 port map( in1 => l0_13_port, in2 => l1_13_port, in3 => 
                           l2_13_port, in4 => l3_13_port, o => o(13));
   g2_a_12 : nand41_13 port map( in1 => l0_12_port, in2 => l1_12_port, in3 => 
                           l2_12_port, in4 => l3_12_port, o => o(12));
   g2_a_11 : nand41_12 port map( in1 => l0_11_port, in2 => l1_11_port, in3 => 
                           l2_11_port, in4 => l3_11_port, o => o(11));
   g2_a_10 : nand41_11 port map( in1 => l0_10_port, in2 => l1_10_port, in3 => 
                           l2_10_port, in4 => l3_10_port, o => o(10));
   g2_a_9 : nand41_10 port map( in1 => l0_9_port, in2 => l1_9_port, in3 => 
                           l2_9_port, in4 => l3_9_port, o => o(9));
   g2_a_8 : nand41_9 port map( in1 => l0_8_port, in2 => l1_8_port, in3 => 
                           l2_8_port, in4 => l3_8_port, o => o(8));
   g2_a_7 : nand41_8 port map( in1 => l0_7_port, in2 => l1_7_port, in3 => 
                           l2_7_port, in4 => l3_7_port, o => o(7));
   g2_a_6 : nand41_7 port map( in1 => l0_6_port, in2 => l1_6_port, in3 => 
                           l2_6_port, in4 => l3_6_port, o => o(6));
   g2_a_5 : nand41_6 port map( in1 => l0_5_port, in2 => l1_5_port, in3 => 
                           l2_5_port, in4 => l3_5_port, o => o(5));
   g2_a_4 : nand41_5 port map( in1 => l0_4_port, in2 => l1_4_port, in3 => 
                           l2_4_port, in4 => l3_4_port, o => o(4));
   g2_a_3 : nand41_4 port map( in1 => l0_3_port, in2 => l1_3_port, in3 => 
                           l2_3_port, in4 => l3_3_port, o => o(3));
   g2_a_2 : nand41_3 port map( in1 => l0_2_port, in2 => l1_2_port, in3 => 
                           l2_2_port, in4 => l3_2_port, o => o(2));
   g2_a_1 : nand41_2 port map( in1 => l0_1_port, in2 => l1_1_port, in3 => 
                           l2_1_port, in4 => l3_1_port, o => o(1));
   g2_a_0 : nand41_1 port map( in1 => l0_0_port, in2 => l1_0_port, in3 => 
                           l2_0_port, in4 => l3_0_port, o => o(0));
   U3 : BUF_X1 port map( A => s0_9_port, Z => n10);
   U4 : BUF_X1 port map( A => s0_9_port, Z => n11);
   U5 : BUF_X1 port map( A => s3_9_port, Z => n2);
   U6 : BUF_X1 port map( A => s3_9_port, Z => n1);
   U7 : BUF_X1 port map( A => s0_9_port, Z => n12);
   U8 : BUF_X1 port map( A => s3_9_port, Z => n3);
   U9 : INV_X1 port map( A => in1(0), ZN => n52);
   U10 : INV_X1 port map( A => in1(28), ZN => n49);
   U11 : INV_X1 port map( A => in1(27), ZN => n48);
   U12 : INV_X1 port map( A => in1(26), ZN => n47);
   U13 : INV_X1 port map( A => in1(25), ZN => n46);
   U14 : INV_X1 port map( A => in1(24), ZN => n45);
   U15 : INV_X1 port map( A => in1(7), ZN => n28);
   U16 : INV_X1 port map( A => in1(6), ZN => n27);
   U17 : INV_X1 port map( A => in1(5), ZN => n26);
   U18 : INV_X1 port map( A => in1(4), ZN => n25);
   U19 : INV_X1 port map( A => in1(3), ZN => n24);
   U20 : INV_X1 port map( A => in1(2), ZN => n23);
   U21 : INV_X1 port map( A => in1(1), ZN => n22);
   U22 : INV_X1 port map( A => in1(23), ZN => n44);
   U23 : INV_X1 port map( A => in1(22), ZN => n43);
   U24 : INV_X1 port map( A => in1(21), ZN => n42);
   U25 : INV_X1 port map( A => in1(20), ZN => n41);
   U26 : INV_X1 port map( A => in1(19), ZN => n40);
   U27 : INV_X1 port map( A => in1(18), ZN => n39);
   U28 : INV_X1 port map( A => in1(17), ZN => n38);
   U29 : INV_X1 port map( A => in1(16), ZN => n37);
   U30 : INV_X1 port map( A => in1(15), ZN => n36);
   U31 : INV_X1 port map( A => in1(14), ZN => n35);
   U32 : INV_X1 port map( A => in1(13), ZN => n34);
   U33 : INV_X1 port map( A => in1(12), ZN => n33);
   U34 : INV_X1 port map( A => in1(11), ZN => n32);
   U35 : INV_X1 port map( A => in1(10), ZN => n31);
   U36 : INV_X1 port map( A => in1(9), ZN => n30);
   U37 : INV_X1 port map( A => in1(8), ZN => n29);
   U38 : INV_X1 port map( A => in1(29), ZN => n50);
   U39 : INV_X1 port map( A => in1(30), ZN => n51);
   U40 : INV_X1 port map( A => in2(5), ZN => n53);
   U41 : BUF_X1 port map( A => s2_9_port, Z => n4);
   U42 : BUF_X1 port map( A => s2_9_port, Z => n5);
   U43 : BUF_X1 port map( A => s2_9_port, Z => n6);
   U44 : BUF_X1 port map( A => s2_9_port, Z => n7);
   U45 : BUF_X1 port map( A => s2_9_port, Z => n8);
   U46 : BUF_X1 port map( A => s2_9_port, Z => n9);
   U47 : OAI21_X1 port map( B1 => n86, B2 => n74, A => n70, ZN => s0_9_port);
   U48 : INV_X1 port map( A => in2(7), ZN => n55);
   U49 : INV_X1 port map( A => in2(6), ZN => n54);
   U50 : INV_X1 port map( A => in2(31), ZN => n85);
   U51 : INV_X1 port map( A => in2(8), ZN => n56);
   U52 : INV_X1 port map( A => in2(30), ZN => n84);
   U53 : INV_X1 port map( A => in2(29), ZN => n83);
   U54 : INV_X1 port map( A => in2(28), ZN => n82);
   U55 : INV_X1 port map( A => in2(27), ZN => n81);
   U56 : INV_X1 port map( A => in2(26), ZN => n80);
   U57 : INV_X1 port map( A => in2(25), ZN => n79);
   U58 : INV_X1 port map( A => in2(24), ZN => n78);
   U59 : INV_X1 port map( A => in2(23), ZN => n77);
   U60 : INV_X1 port map( A => in2(22), ZN => n76);
   U61 : INV_X1 port map( A => in2(21), ZN => n75);
   U62 : INV_X1 port map( A => in2(20), ZN => n68);
   U63 : INV_X1 port map( A => in2(19), ZN => n67);
   U64 : INV_X1 port map( A => in2(18), ZN => n66);
   U65 : INV_X1 port map( A => in2(17), ZN => n65);
   U66 : INV_X1 port map( A => in2(16), ZN => n64);
   U67 : INV_X1 port map( A => in2(15), ZN => n63);
   U68 : INV_X1 port map( A => in2(14), ZN => n62);
   U69 : INV_X1 port map( A => in2(13), ZN => n61);
   U70 : INV_X1 port map( A => in2(12), ZN => n60);
   U71 : INV_X1 port map( A => in2(11), ZN => n59);
   U72 : INV_X1 port map( A => in2(10), ZN => n58);
   U73 : INV_X1 port map( A => in2(9), ZN => n57);
   U74 : AND2_X1 port map( A1 => n69, A2 => n70, ZN => s3_9_port);
   U75 : NAND2_X1 port map( A1 => SN, A2 => n73, ZN => n70);
   U76 : INV_X1 port map( A => SN, ZN => n86);
   U80 : OR2_X1 port map( A1 => n74, A2 => SN, ZN => n69);
   U81 : NOR3_X1 port map( A1 => func(2), A2 => func(3), A3 => n20, ZN => n73);
   U82 : NAND4_X1 port map( A1 => func(2), A2 => n21, A3 => n20, A4 => n19, ZN 
                           => n74);
   U83 : INV_X1 port map( A => func(3), ZN => n19);
   U84 : INV_X1 port map( A => func(1), ZN => n20);
   U85 : INV_X1 port map( A => func(0), ZN => n21);
   U86 : INV_X1 port map( A => in2(0), ZN => n13);
   U87 : INV_X1 port map( A => in2(1), ZN => n14);
   U88 : INV_X1 port map( A => in2(2), ZN => n15);
   U89 : INV_X1 port map( A => in2(3), ZN => n16);
   U90 : INV_X1 port map( A => in2(4), ZN => n17);
   U91 : INV_X1 port map( A => in1(31), ZN => n18);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity shifter_NBITS32 is

   port( R1, R2 : in std_logic_vector (31 downto 0);  LnR, AnL, RnS : in 
         std_logic;  Rout : out std_logic_vector (31 downto 0));

end shifter_NBITS32;

architecture SYN_structural of shifter_NBITS32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX81_GENERIC_NBIT32
      port( A, B, C, D, E, F, G, H : in std_logic_vector (31 downto 0);  SEL : 
            in std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 
            downto 0));
   end component;
   
   component mask_shifter_NBITS40
      port( R1 : in std_logic_vector (39 downto 0);  LnR : in std_logic;  
            mask_sh0, mask_sh1, mask_sh2, mask_sh3, mask_sh4, mask_sh5, 
            mask_sh6, mask_sh7 : out std_logic_vector (31 downto 0));
   end component;
   
   component MUX41_GENERIC_NBIT40
      port( A, B, C, D : in std_logic_vector (39 downto 0);  SEL : in 
            std_logic_vector (1 downto 0);  Y : out std_logic_vector (39 downto
            0));
   end component;
   
   component mask_generator_NBITS32
      port( R1, R2 : in std_logic_vector (31 downto 0);  LnR, AnL, RnS : in 
            std_logic;  mask0, mask8, mask16, mask24 : out std_logic_vector (39
            downto 0));
   end component;
   
   signal s_RnS, s_mask0_39_port, s_mask0_38_port, s_mask0_37_port, 
      s_mask0_36_port, s_mask0_35_port, s_mask0_34_port, s_mask0_33_port, 
      s_mask0_32_port, s_mask0_31_port, s_mask0_30_port, s_mask0_29_port, 
      s_mask0_28_port, s_mask0_27_port, s_mask0_26_port, s_mask0_25_port, 
      s_mask0_24_port, s_mask0_23_port, s_mask0_22_port, s_mask0_21_port, 
      s_mask0_20_port, s_mask0_19_port, s_mask0_18_port, s_mask0_17_port, 
      s_mask0_16_port, s_mask0_15_port, s_mask0_14_port, s_mask0_13_port, 
      s_mask0_12_port, s_mask0_11_port, s_mask0_10_port, s_mask0_9_port, 
      s_mask0_8_port, s_mask0_7_port, s_mask0_6_port, s_mask0_5_port, 
      s_mask0_4_port, s_mask0_3_port, s_mask0_2_port, s_mask0_1_port, 
      s_mask0_0_port, s_mask8_39_port, s_mask8_38_port, s_mask8_37_port, 
      s_mask8_36_port, s_mask8_35_port, s_mask8_34_port, s_mask8_33_port, 
      s_mask8_32_port, s_mask8_31_port, s_mask8_30_port, s_mask8_29_port, 
      s_mask8_28_port, s_mask8_27_port, s_mask8_26_port, s_mask8_25_port, 
      s_mask8_24_port, s_mask8_23_port, s_mask8_22_port, s_mask8_21_port, 
      s_mask8_20_port, s_mask8_19_port, s_mask8_18_port, s_mask8_17_port, 
      s_mask8_16_port, s_mask8_15_port, s_mask8_14_port, s_mask8_13_port, 
      s_mask8_12_port, s_mask8_11_port, s_mask8_10_port, s_mask8_9_port, 
      s_mask8_8_port, s_mask8_7_port, s_mask8_6_port, s_mask8_5_port, 
      s_mask8_4_port, s_mask8_3_port, s_mask8_2_port, s_mask8_1_port, 
      s_mask8_0_port, s_mask16_39_port, s_mask16_38_port, s_mask16_37_port, 
      s_mask16_36_port, s_mask16_35_port, s_mask16_34_port, s_mask16_33_port, 
      s_mask16_32_port, s_mask16_31_port, s_mask16_30_port, s_mask16_29_port, 
      s_mask16_28_port, s_mask16_27_port, s_mask16_26_port, s_mask16_25_port, 
      s_mask16_24_port, s_mask16_23_port, s_mask16_22_port, s_mask16_21_port, 
      s_mask16_20_port, s_mask16_19_port, s_mask16_18_port, s_mask16_17_port, 
      s_mask16_16_port, s_mask16_15_port, s_mask16_14_port, s_mask16_13_port, 
      s_mask16_12_port, s_mask16_11_port, s_mask16_10_port, s_mask16_9_port, 
      s_mask16_8_port, s_mask16_7_port, s_mask16_6_port, s_mask16_5_port, 
      s_mask16_4_port, s_mask16_3_port, s_mask16_2_port, s_mask16_1_port, 
      s_mask16_0_port, s_mask24_39_port, s_mask24_38_port, s_mask24_37_port, 
      s_mask24_36_port, s_mask24_35_port, s_mask24_34_port, s_mask24_33_port, 
      s_mask24_32_port, s_mask24_31_port, s_mask24_30_port, s_mask24_29_port, 
      s_mask24_28_port, s_mask24_27_port, s_mask24_26_port, s_mask24_25_port, 
      s_mask24_24_port, s_mask24_23_port, s_mask24_22_port, s_mask24_21_port, 
      s_mask24_20_port, s_mask24_19_port, s_mask24_18_port, s_mask24_17_port, 
      s_mask24_16_port, s_mask24_15_port, s_mask24_14_port, s_mask24_13_port, 
      s_mask24_12_port, s_mask24_11_port, s_mask24_10_port, s_mask24_9_port, 
      s_mask24_8_port, s_mask24_7_port, s_mask24_6_port, s_mask24_5_port, 
      s_mask24_4_port, s_mask24_3_port, s_mask24_2_port, s_mask24_1_port, 
      s_mask24_0_port, s_selected_mask_39_port, s_selected_mask_38_port, 
      s_selected_mask_37_port, s_selected_mask_36_port, s_selected_mask_35_port
      , s_selected_mask_34_port, s_selected_mask_33_port, 
      s_selected_mask_32_port, s_selected_mask_31_port, s_selected_mask_30_port
      , s_selected_mask_29_port, s_selected_mask_28_port, 
      s_selected_mask_27_port, s_selected_mask_26_port, s_selected_mask_25_port
      , s_selected_mask_24_port, s_selected_mask_23_port, 
      s_selected_mask_22_port, s_selected_mask_21_port, s_selected_mask_20_port
      , s_selected_mask_19_port, s_selected_mask_18_port, 
      s_selected_mask_17_port, s_selected_mask_16_port, s_selected_mask_15_port
      , s_selected_mask_14_port, s_selected_mask_13_port, 
      s_selected_mask_12_port, s_selected_mask_11_port, s_selected_mask_10_port
      , s_selected_mask_9_port, s_selected_mask_8_port, s_selected_mask_7_port,
      s_selected_mask_6_port, s_selected_mask_5_port, s_selected_mask_4_port, 
      s_selected_mask_3_port, s_selected_mask_2_port, s_selected_mask_1_port, 
      s_selected_mask_0_port, s_sh0_31_port, s_sh0_30_port, s_sh0_29_port, 
      s_sh0_28_port, s_sh0_27_port, s_sh0_26_port, s_sh0_25_port, s_sh0_24_port
      , s_sh0_23_port, s_sh0_22_port, s_sh0_21_port, s_sh0_20_port, 
      s_sh0_19_port, s_sh0_18_port, s_sh0_17_port, s_sh0_16_port, s_sh0_15_port
      , s_sh0_14_port, s_sh0_13_port, s_sh0_12_port, s_sh0_11_port, 
      s_sh0_10_port, s_sh0_9_port, s_sh0_8_port, s_sh0_7_port, s_sh0_6_port, 
      s_sh0_5_port, s_sh0_4_port, s_sh0_3_port, s_sh0_2_port, s_sh0_1_port, 
      s_sh0_0_port, s_sh1_31_port, s_sh1_30_port, s_sh1_29_port, s_sh1_28_port,
      s_sh1_27_port, s_sh1_26_port, s_sh1_25_port, s_sh1_24_port, s_sh1_23_port
      , s_sh1_22_port, s_sh1_21_port, s_sh1_20_port, s_sh1_19_port, 
      s_sh1_18_port, s_sh1_17_port, s_sh1_16_port, s_sh1_15_port, s_sh1_14_port
      , s_sh1_13_port, s_sh1_12_port, s_sh1_11_port, s_sh1_10_port, 
      s_sh1_9_port, s_sh1_8_port, s_sh1_7_port, s_sh1_6_port, s_sh1_5_port, 
      s_sh1_4_port, s_sh1_3_port, s_sh1_2_port, s_sh1_1_port, s_sh1_0_port, 
      s_sh2_31_port, s_sh2_30_port, s_sh2_29_port, s_sh2_28_port, s_sh2_27_port
      , s_sh2_26_port, s_sh2_25_port, s_sh2_24_port, s_sh2_23_port, 
      s_sh2_22_port, s_sh2_21_port, s_sh2_20_port, s_sh2_19_port, s_sh2_18_port
      , s_sh2_17_port, s_sh2_16_port, s_sh2_15_port, s_sh2_14_port, 
      s_sh2_13_port, s_sh2_12_port, s_sh2_11_port, s_sh2_10_port, s_sh2_9_port,
      s_sh2_8_port, s_sh2_7_port, s_sh2_6_port, s_sh2_5_port, s_sh2_4_port, 
      s_sh2_3_port, s_sh2_2_port, s_sh2_1_port, s_sh2_0_port, s_sh3_31_port, 
      s_sh3_30_port, s_sh3_29_port, s_sh3_28_port, s_sh3_27_port, s_sh3_26_port
      , s_sh3_25_port, s_sh3_24_port, s_sh3_23_port, s_sh3_22_port, 
      s_sh3_21_port, s_sh3_20_port, s_sh3_19_port, s_sh3_18_port, s_sh3_17_port
      , s_sh3_16_port, s_sh3_15_port, s_sh3_14_port, s_sh3_13_port, 
      s_sh3_12_port, s_sh3_11_port, s_sh3_10_port, s_sh3_9_port, s_sh3_8_port, 
      s_sh3_7_port, s_sh3_6_port, s_sh3_5_port, s_sh3_4_port, s_sh3_3_port, 
      s_sh3_2_port, s_sh3_1_port, s_sh3_0_port, s_sh4_31_port, s_sh4_30_port, 
      s_sh4_29_port, s_sh4_28_port, s_sh4_27_port, s_sh4_26_port, s_sh4_25_port
      , s_sh4_24_port, s_sh4_23_port, s_sh4_22_port, s_sh4_21_port, 
      s_sh4_20_port, s_sh4_19_port, s_sh4_18_port, s_sh4_17_port, s_sh4_16_port
      , s_sh4_15_port, s_sh4_14_port, s_sh4_13_port, s_sh4_12_port, 
      s_sh4_11_port, s_sh4_10_port, s_sh4_9_port, s_sh4_8_port, s_sh4_7_port, 
      s_sh4_6_port, s_sh4_5_port, s_sh4_4_port, s_sh4_3_port, s_sh4_2_port, 
      s_sh4_1_port, s_sh4_0_port, s_sh5_31_port, s_sh5_30_port, s_sh5_29_port, 
      s_sh5_28_port, s_sh5_27_port, s_sh5_26_port, s_sh5_25_port, s_sh5_24_port
      , s_sh5_23_port, s_sh5_22_port, s_sh5_21_port, s_sh5_20_port, 
      s_sh5_19_port, s_sh5_18_port, s_sh5_17_port, s_sh5_16_port, s_sh5_15_port
      , s_sh5_14_port, s_sh5_13_port, s_sh5_12_port, s_sh5_11_port, 
      s_sh5_10_port, s_sh5_9_port, s_sh5_8_port, s_sh5_7_port, s_sh5_6_port, 
      s_sh5_5_port, s_sh5_4_port, s_sh5_3_port, s_sh5_2_port, s_sh5_1_port, 
      s_sh5_0_port, s_sh6_31_port, s_sh6_30_port, s_sh6_29_port, s_sh6_28_port,
      s_sh6_27_port, s_sh6_26_port, s_sh6_25_port, s_sh6_24_port, s_sh6_23_port
      , s_sh6_22_port, s_sh6_21_port, s_sh6_20_port, s_sh6_19_port, 
      s_sh6_18_port, s_sh6_17_port, s_sh6_16_port, s_sh6_15_port, s_sh6_14_port
      , s_sh6_13_port, s_sh6_12_port, s_sh6_11_port, s_sh6_10_port, 
      s_sh6_9_port, s_sh6_8_port, s_sh6_7_port, s_sh6_6_port, s_sh6_5_port, 
      s_sh6_4_port, s_sh6_3_port, s_sh6_2_port, s_sh6_1_port, s_sh6_0_port, 
      s_sh7_31_port, s_sh7_30_port, s_sh7_29_port, s_sh7_28_port, s_sh7_27_port
      , s_sh7_26_port, s_sh7_25_port, s_sh7_24_port, s_sh7_23_port, 
      s_sh7_22_port, s_sh7_21_port, s_sh7_20_port, s_sh7_19_port, s_sh7_18_port
      , s_sh7_17_port, s_sh7_16_port, s_sh7_15_port, s_sh7_14_port, 
      s_sh7_13_port, s_sh7_12_port, s_sh7_11_port, s_sh7_10_port, s_sh7_9_port,
      s_sh7_8_port, s_sh7_7_port, s_sh7_6_port, s_sh7_5_port, s_sh7_4_port, 
      s_sh7_3_port, s_sh7_2_port, s_sh7_1_port, s_sh7_0_port, n1 : std_logic;

begin
   
   mask_gen : mask_generator_NBITS32 port map( R1(31) => R1(31), R1(30) => 
                           R1(30), R1(29) => R1(29), R1(28) => R1(28), R1(27) 
                           => R1(27), R1(26) => R1(26), R1(25) => R1(25), 
                           R1(24) => R1(24), R1(23) => R1(23), R1(22) => R1(22)
                           , R1(21) => R1(21), R1(20) => R1(20), R1(19) => 
                           R1(19), R1(18) => R1(18), R1(17) => R1(17), R1(16) 
                           => R1(16), R1(15) => R1(15), R1(14) => R1(14), 
                           R1(13) => R1(13), R1(12) => R1(12), R1(11) => R1(11)
                           , R1(10) => R1(10), R1(9) => R1(9), R1(8) => R1(8), 
                           R1(7) => R1(7), R1(6) => R1(6), R1(5) => R1(5), 
                           R1(4) => R1(4), R1(3) => R1(3), R1(2) => R1(2), 
                           R1(1) => R1(1), R1(0) => R1(0), R2(31) => R2(31), 
                           R2(30) => R2(30), R2(29) => R2(29), R2(28) => R2(28)
                           , R2(27) => R2(27), R2(26) => R2(26), R2(25) => 
                           R2(25), R2(24) => R2(24), R2(23) => R2(23), R2(22) 
                           => R2(22), R2(21) => R2(21), R2(20) => R2(20), 
                           R2(19) => R2(19), R2(18) => R2(18), R2(17) => R2(17)
                           , R2(16) => R2(16), R2(15) => R2(15), R2(14) => 
                           R2(14), R2(13) => R2(13), R2(12) => R2(12), R2(11) 
                           => R2(11), R2(10) => R2(10), R2(9) => R2(9), R2(8) 
                           => R2(8), R2(7) => R2(7), R2(6) => R2(6), R2(5) => 
                           R2(5), R2(4) => R2(4), R2(3) => R2(3), R2(2) => 
                           R2(2), R2(1) => R2(1), R2(0) => R2(0), LnR => LnR, 
                           AnL => AnL, RnS => s_RnS, mask0(39) => 
                           s_mask0_39_port, mask0(38) => s_mask0_38_port, 
                           mask0(37) => s_mask0_37_port, mask0(36) => 
                           s_mask0_36_port, mask0(35) => s_mask0_35_port, 
                           mask0(34) => s_mask0_34_port, mask0(33) => 
                           s_mask0_33_port, mask0(32) => s_mask0_32_port, 
                           mask0(31) => s_mask0_31_port, mask0(30) => 
                           s_mask0_30_port, mask0(29) => s_mask0_29_port, 
                           mask0(28) => s_mask0_28_port, mask0(27) => 
                           s_mask0_27_port, mask0(26) => s_mask0_26_port, 
                           mask0(25) => s_mask0_25_port, mask0(24) => 
                           s_mask0_24_port, mask0(23) => s_mask0_23_port, 
                           mask0(22) => s_mask0_22_port, mask0(21) => 
                           s_mask0_21_port, mask0(20) => s_mask0_20_port, 
                           mask0(19) => s_mask0_19_port, mask0(18) => 
                           s_mask0_18_port, mask0(17) => s_mask0_17_port, 
                           mask0(16) => s_mask0_16_port, mask0(15) => 
                           s_mask0_15_port, mask0(14) => s_mask0_14_port, 
                           mask0(13) => s_mask0_13_port, mask0(12) => 
                           s_mask0_12_port, mask0(11) => s_mask0_11_port, 
                           mask0(10) => s_mask0_10_port, mask0(9) => 
                           s_mask0_9_port, mask0(8) => s_mask0_8_port, mask0(7)
                           => s_mask0_7_port, mask0(6) => s_mask0_6_port, 
                           mask0(5) => s_mask0_5_port, mask0(4) => 
                           s_mask0_4_port, mask0(3) => s_mask0_3_port, mask0(2)
                           => s_mask0_2_port, mask0(1) => s_mask0_1_port, 
                           mask0(0) => s_mask0_0_port, mask8(39) => 
                           s_mask8_39_port, mask8(38) => s_mask8_38_port, 
                           mask8(37) => s_mask8_37_port, mask8(36) => 
                           s_mask8_36_port, mask8(35) => s_mask8_35_port, 
                           mask8(34) => s_mask8_34_port, mask8(33) => 
                           s_mask8_33_port, mask8(32) => s_mask8_32_port, 
                           mask8(31) => s_mask8_31_port, mask8(30) => 
                           s_mask8_30_port, mask8(29) => s_mask8_29_port, 
                           mask8(28) => s_mask8_28_port, mask8(27) => 
                           s_mask8_27_port, mask8(26) => s_mask8_26_port, 
                           mask8(25) => s_mask8_25_port, mask8(24) => 
                           s_mask8_24_port, mask8(23) => s_mask8_23_port, 
                           mask8(22) => s_mask8_22_port, mask8(21) => 
                           s_mask8_21_port, mask8(20) => s_mask8_20_port, 
                           mask8(19) => s_mask8_19_port, mask8(18) => 
                           s_mask8_18_port, mask8(17) => s_mask8_17_port, 
                           mask8(16) => s_mask8_16_port, mask8(15) => 
                           s_mask8_15_port, mask8(14) => s_mask8_14_port, 
                           mask8(13) => s_mask8_13_port, mask8(12) => 
                           s_mask8_12_port, mask8(11) => s_mask8_11_port, 
                           mask8(10) => s_mask8_10_port, mask8(9) => 
                           s_mask8_9_port, mask8(8) => s_mask8_8_port, mask8(7)
                           => s_mask8_7_port, mask8(6) => s_mask8_6_port, 
                           mask8(5) => s_mask8_5_port, mask8(4) => 
                           s_mask8_4_port, mask8(3) => s_mask8_3_port, mask8(2)
                           => s_mask8_2_port, mask8(1) => s_mask8_1_port, 
                           mask8(0) => s_mask8_0_port, mask16(39) => 
                           s_mask16_39_port, mask16(38) => s_mask16_38_port, 
                           mask16(37) => s_mask16_37_port, mask16(36) => 
                           s_mask16_36_port, mask16(35) => s_mask16_35_port, 
                           mask16(34) => s_mask16_34_port, mask16(33) => 
                           s_mask16_33_port, mask16(32) => s_mask16_32_port, 
                           mask16(31) => s_mask16_31_port, mask16(30) => 
                           s_mask16_30_port, mask16(29) => s_mask16_29_port, 
                           mask16(28) => s_mask16_28_port, mask16(27) => 
                           s_mask16_27_port, mask16(26) => s_mask16_26_port, 
                           mask16(25) => s_mask16_25_port, mask16(24) => 
                           s_mask16_24_port, mask16(23) => s_mask16_23_port, 
                           mask16(22) => s_mask16_22_port, mask16(21) => 
                           s_mask16_21_port, mask16(20) => s_mask16_20_port, 
                           mask16(19) => s_mask16_19_port, mask16(18) => 
                           s_mask16_18_port, mask16(17) => s_mask16_17_port, 
                           mask16(16) => s_mask16_16_port, mask16(15) => 
                           s_mask16_15_port, mask16(14) => s_mask16_14_port, 
                           mask16(13) => s_mask16_13_port, mask16(12) => 
                           s_mask16_12_port, mask16(11) => s_mask16_11_port, 
                           mask16(10) => s_mask16_10_port, mask16(9) => 
                           s_mask16_9_port, mask16(8) => s_mask16_8_port, 
                           mask16(7) => s_mask16_7_port, mask16(6) => 
                           s_mask16_6_port, mask16(5) => s_mask16_5_port, 
                           mask16(4) => s_mask16_4_port, mask16(3) => 
                           s_mask16_3_port, mask16(2) => s_mask16_2_port, 
                           mask16(1) => s_mask16_1_port, mask16(0) => 
                           s_mask16_0_port, mask24(39) => s_mask24_39_port, 
                           mask24(38) => s_mask24_38_port, mask24(37) => 
                           s_mask24_37_port, mask24(36) => s_mask24_36_port, 
                           mask24(35) => s_mask24_35_port, mask24(34) => 
                           s_mask24_34_port, mask24(33) => s_mask24_33_port, 
                           mask24(32) => s_mask24_32_port, mask24(31) => 
                           s_mask24_31_port, mask24(30) => s_mask24_30_port, 
                           mask24(29) => s_mask24_29_port, mask24(28) => 
                           s_mask24_28_port, mask24(27) => s_mask24_27_port, 
                           mask24(26) => s_mask24_26_port, mask24(25) => 
                           s_mask24_25_port, mask24(24) => s_mask24_24_port, 
                           mask24(23) => s_mask24_23_port, mask24(22) => 
                           s_mask24_22_port, mask24(21) => s_mask24_21_port, 
                           mask24(20) => s_mask24_20_port, mask24(19) => 
                           s_mask24_19_port, mask24(18) => s_mask24_18_port, 
                           mask24(17) => s_mask24_17_port, mask24(16) => 
                           s_mask24_16_port, mask24(15) => s_mask24_15_port, 
                           mask24(14) => s_mask24_14_port, mask24(13) => 
                           s_mask24_13_port, mask24(12) => s_mask24_12_port, 
                           mask24(11) => s_mask24_11_port, mask24(10) => 
                           s_mask24_10_port, mask24(9) => s_mask24_9_port, 
                           mask24(8) => s_mask24_8_port, mask24(7) => 
                           s_mask24_7_port, mask24(6) => s_mask24_6_port, 
                           mask24(5) => s_mask24_5_port, mask24(4) => 
                           s_mask24_4_port, mask24(3) => s_mask24_3_port, 
                           mask24(2) => s_mask24_2_port, mask24(1) => 
                           s_mask24_1_port, mask24(0) => s_mask24_0_port);
   MUX_mask_select : MUX41_GENERIC_NBIT40 port map( A(39) => s_mask0_39_port, 
                           A(38) => s_mask0_38_port, A(37) => s_mask0_37_port, 
                           A(36) => s_mask0_36_port, A(35) => s_mask0_35_port, 
                           A(34) => s_mask0_34_port, A(33) => s_mask0_33_port, 
                           A(32) => s_mask0_32_port, A(31) => s_mask0_31_port, 
                           A(30) => s_mask0_30_port, A(29) => s_mask0_29_port, 
                           A(28) => s_mask0_28_port, A(27) => s_mask0_27_port, 
                           A(26) => s_mask0_26_port, A(25) => s_mask0_25_port, 
                           A(24) => s_mask0_24_port, A(23) => s_mask0_23_port, 
                           A(22) => s_mask0_22_port, A(21) => s_mask0_21_port, 
                           A(20) => s_mask0_20_port, A(19) => s_mask0_19_port, 
                           A(18) => s_mask0_18_port, A(17) => s_mask0_17_port, 
                           A(16) => s_mask0_16_port, A(15) => s_mask0_15_port, 
                           A(14) => s_mask0_14_port, A(13) => s_mask0_13_port, 
                           A(12) => s_mask0_12_port, A(11) => s_mask0_11_port, 
                           A(10) => s_mask0_10_port, A(9) => s_mask0_9_port, 
                           A(8) => s_mask0_8_port, A(7) => s_mask0_7_port, A(6)
                           => s_mask0_6_port, A(5) => s_mask0_5_port, A(4) => 
                           s_mask0_4_port, A(3) => s_mask0_3_port, A(2) => 
                           s_mask0_2_port, A(1) => s_mask0_1_port, A(0) => 
                           s_mask0_0_port, B(39) => s_mask8_39_port, B(38) => 
                           s_mask8_38_port, B(37) => s_mask8_37_port, B(36) => 
                           s_mask8_36_port, B(35) => s_mask8_35_port, B(34) => 
                           s_mask8_34_port, B(33) => s_mask8_33_port, B(32) => 
                           s_mask8_32_port, B(31) => s_mask8_31_port, B(30) => 
                           s_mask8_30_port, B(29) => s_mask8_29_port, B(28) => 
                           s_mask8_28_port, B(27) => s_mask8_27_port, B(26) => 
                           s_mask8_26_port, B(25) => s_mask8_25_port, B(24) => 
                           s_mask8_24_port, B(23) => s_mask8_23_port, B(22) => 
                           s_mask8_22_port, B(21) => s_mask8_21_port, B(20) => 
                           s_mask8_20_port, B(19) => s_mask8_19_port, B(18) => 
                           s_mask8_18_port, B(17) => s_mask8_17_port, B(16) => 
                           s_mask8_16_port, B(15) => s_mask8_15_port, B(14) => 
                           s_mask8_14_port, B(13) => s_mask8_13_port, B(12) => 
                           s_mask8_12_port, B(11) => s_mask8_11_port, B(10) => 
                           s_mask8_10_port, B(9) => s_mask8_9_port, B(8) => 
                           s_mask8_8_port, B(7) => s_mask8_7_port, B(6) => 
                           s_mask8_6_port, B(5) => s_mask8_5_port, B(4) => 
                           s_mask8_4_port, B(3) => s_mask8_3_port, B(2) => 
                           s_mask8_2_port, B(1) => s_mask8_1_port, B(0) => 
                           s_mask8_0_port, C(39) => s_mask16_39_port, C(38) => 
                           s_mask16_38_port, C(37) => s_mask16_37_port, C(36) 
                           => s_mask16_36_port, C(35) => s_mask16_35_port, 
                           C(34) => s_mask16_34_port, C(33) => s_mask16_33_port
                           , C(32) => s_mask16_32_port, C(31) => 
                           s_mask16_31_port, C(30) => s_mask16_30_port, C(29) 
                           => s_mask16_29_port, C(28) => s_mask16_28_port, 
                           C(27) => s_mask16_27_port, C(26) => s_mask16_26_port
                           , C(25) => s_mask16_25_port, C(24) => 
                           s_mask16_24_port, C(23) => s_mask16_23_port, C(22) 
                           => s_mask16_22_port, C(21) => s_mask16_21_port, 
                           C(20) => s_mask16_20_port, C(19) => s_mask16_19_port
                           , C(18) => s_mask16_18_port, C(17) => 
                           s_mask16_17_port, C(16) => s_mask16_16_port, C(15) 
                           => s_mask16_15_port, C(14) => s_mask16_14_port, 
                           C(13) => s_mask16_13_port, C(12) => s_mask16_12_port
                           , C(11) => s_mask16_11_port, C(10) => 
                           s_mask16_10_port, C(9) => s_mask16_9_port, C(8) => 
                           s_mask16_8_port, C(7) => s_mask16_7_port, C(6) => 
                           s_mask16_6_port, C(5) => s_mask16_5_port, C(4) => 
                           s_mask16_4_port, C(3) => s_mask16_3_port, C(2) => 
                           s_mask16_2_port, C(1) => s_mask16_1_port, C(0) => 
                           s_mask16_0_port, D(39) => s_mask24_39_port, D(38) =>
                           s_mask24_38_port, D(37) => s_mask24_37_port, D(36) 
                           => s_mask24_36_port, D(35) => s_mask24_35_port, 
                           D(34) => s_mask24_34_port, D(33) => s_mask24_33_port
                           , D(32) => s_mask24_32_port, D(31) => 
                           s_mask24_31_port, D(30) => s_mask24_30_port, D(29) 
                           => s_mask24_29_port, D(28) => s_mask24_28_port, 
                           D(27) => s_mask24_27_port, D(26) => s_mask24_26_port
                           , D(25) => s_mask24_25_port, D(24) => 
                           s_mask24_24_port, D(23) => s_mask24_23_port, D(22) 
                           => s_mask24_22_port, D(21) => s_mask24_21_port, 
                           D(20) => s_mask24_20_port, D(19) => s_mask24_19_port
                           , D(18) => s_mask24_18_port, D(17) => 
                           s_mask24_17_port, D(16) => s_mask24_16_port, D(15) 
                           => s_mask24_15_port, D(14) => s_mask24_14_port, 
                           D(13) => s_mask24_13_port, D(12) => s_mask24_12_port
                           , D(11) => s_mask24_11_port, D(10) => 
                           s_mask24_10_port, D(9) => s_mask24_9_port, D(8) => 
                           s_mask24_8_port, D(7) => s_mask24_7_port, D(6) => 
                           s_mask24_6_port, D(5) => s_mask24_5_port, D(4) => 
                           s_mask24_4_port, D(3) => s_mask24_3_port, D(2) => 
                           s_mask24_2_port, D(1) => s_mask24_1_port, D(0) => 
                           s_mask24_0_port, SEL(1) => R2(4), SEL(0) => R2(3), 
                           Y(39) => s_selected_mask_39_port, Y(38) => 
                           s_selected_mask_38_port, Y(37) => 
                           s_selected_mask_37_port, Y(36) => 
                           s_selected_mask_36_port, Y(35) => 
                           s_selected_mask_35_port, Y(34) => 
                           s_selected_mask_34_port, Y(33) => 
                           s_selected_mask_33_port, Y(32) => 
                           s_selected_mask_32_port, Y(31) => 
                           s_selected_mask_31_port, Y(30) => 
                           s_selected_mask_30_port, Y(29) => 
                           s_selected_mask_29_port, Y(28) => 
                           s_selected_mask_28_port, Y(27) => 
                           s_selected_mask_27_port, Y(26) => 
                           s_selected_mask_26_port, Y(25) => 
                           s_selected_mask_25_port, Y(24) => 
                           s_selected_mask_24_port, Y(23) => 
                           s_selected_mask_23_port, Y(22) => 
                           s_selected_mask_22_port, Y(21) => 
                           s_selected_mask_21_port, Y(20) => 
                           s_selected_mask_20_port, Y(19) => 
                           s_selected_mask_19_port, Y(18) => 
                           s_selected_mask_18_port, Y(17) => 
                           s_selected_mask_17_port, Y(16) => 
                           s_selected_mask_16_port, Y(15) => 
                           s_selected_mask_15_port, Y(14) => 
                           s_selected_mask_14_port, Y(13) => 
                           s_selected_mask_13_port, Y(12) => 
                           s_selected_mask_12_port, Y(11) => 
                           s_selected_mask_11_port, Y(10) => 
                           s_selected_mask_10_port, Y(9) => 
                           s_selected_mask_9_port, Y(8) => 
                           s_selected_mask_8_port, Y(7) => 
                           s_selected_mask_7_port, Y(6) => 
                           s_selected_mask_6_port, Y(5) => 
                           s_selected_mask_5_port, Y(4) => 
                           s_selected_mask_4_port, Y(3) => 
                           s_selected_mask_3_port, Y(2) => 
                           s_selected_mask_2_port, Y(1) => 
                           s_selected_mask_1_port, Y(0) => 
                           s_selected_mask_0_port);
   mask_shift : mask_shifter_NBITS40 port map( R1(39) => 
                           s_selected_mask_39_port, R1(38) => 
                           s_selected_mask_38_port, R1(37) => 
                           s_selected_mask_37_port, R1(36) => 
                           s_selected_mask_36_port, R1(35) => 
                           s_selected_mask_35_port, R1(34) => 
                           s_selected_mask_34_port, R1(33) => 
                           s_selected_mask_33_port, R1(32) => 
                           s_selected_mask_32_port, R1(31) => 
                           s_selected_mask_31_port, R1(30) => 
                           s_selected_mask_30_port, R1(29) => 
                           s_selected_mask_29_port, R1(28) => 
                           s_selected_mask_28_port, R1(27) => 
                           s_selected_mask_27_port, R1(26) => 
                           s_selected_mask_26_port, R1(25) => 
                           s_selected_mask_25_port, R1(24) => 
                           s_selected_mask_24_port, R1(23) => 
                           s_selected_mask_23_port, R1(22) => 
                           s_selected_mask_22_port, R1(21) => 
                           s_selected_mask_21_port, R1(20) => 
                           s_selected_mask_20_port, R1(19) => 
                           s_selected_mask_19_port, R1(18) => 
                           s_selected_mask_18_port, R1(17) => 
                           s_selected_mask_17_port, R1(16) => 
                           s_selected_mask_16_port, R1(15) => 
                           s_selected_mask_15_port, R1(14) => 
                           s_selected_mask_14_port, R1(13) => 
                           s_selected_mask_13_port, R1(12) => 
                           s_selected_mask_12_port, R1(11) => 
                           s_selected_mask_11_port, R1(10) => 
                           s_selected_mask_10_port, R1(9) => 
                           s_selected_mask_9_port, R1(8) => 
                           s_selected_mask_8_port, R1(7) => 
                           s_selected_mask_7_port, R1(6) => 
                           s_selected_mask_6_port, R1(5) => 
                           s_selected_mask_5_port, R1(4) => 
                           s_selected_mask_4_port, R1(3) => 
                           s_selected_mask_3_port, R1(2) => 
                           s_selected_mask_2_port, R1(1) => 
                           s_selected_mask_1_port, R1(0) => 
                           s_selected_mask_0_port, LnR => LnR, mask_sh0(31) => 
                           s_sh0_31_port, mask_sh0(30) => s_sh0_30_port, 
                           mask_sh0(29) => s_sh0_29_port, mask_sh0(28) => 
                           s_sh0_28_port, mask_sh0(27) => s_sh0_27_port, 
                           mask_sh0(26) => s_sh0_26_port, mask_sh0(25) => 
                           s_sh0_25_port, mask_sh0(24) => s_sh0_24_port, 
                           mask_sh0(23) => s_sh0_23_port, mask_sh0(22) => 
                           s_sh0_22_port, mask_sh0(21) => s_sh0_21_port, 
                           mask_sh0(20) => s_sh0_20_port, mask_sh0(19) => 
                           s_sh0_19_port, mask_sh0(18) => s_sh0_18_port, 
                           mask_sh0(17) => s_sh0_17_port, mask_sh0(16) => 
                           s_sh0_16_port, mask_sh0(15) => s_sh0_15_port, 
                           mask_sh0(14) => s_sh0_14_port, mask_sh0(13) => 
                           s_sh0_13_port, mask_sh0(12) => s_sh0_12_port, 
                           mask_sh0(11) => s_sh0_11_port, mask_sh0(10) => 
                           s_sh0_10_port, mask_sh0(9) => s_sh0_9_port, 
                           mask_sh0(8) => s_sh0_8_port, mask_sh0(7) => 
                           s_sh0_7_port, mask_sh0(6) => s_sh0_6_port, 
                           mask_sh0(5) => s_sh0_5_port, mask_sh0(4) => 
                           s_sh0_4_port, mask_sh0(3) => s_sh0_3_port, 
                           mask_sh0(2) => s_sh0_2_port, mask_sh0(1) => 
                           s_sh0_1_port, mask_sh0(0) => s_sh0_0_port, 
                           mask_sh1(31) => s_sh1_31_port, mask_sh1(30) => 
                           s_sh1_30_port, mask_sh1(29) => s_sh1_29_port, 
                           mask_sh1(28) => s_sh1_28_port, mask_sh1(27) => 
                           s_sh1_27_port, mask_sh1(26) => s_sh1_26_port, 
                           mask_sh1(25) => s_sh1_25_port, mask_sh1(24) => 
                           s_sh1_24_port, mask_sh1(23) => s_sh1_23_port, 
                           mask_sh1(22) => s_sh1_22_port, mask_sh1(21) => 
                           s_sh1_21_port, mask_sh1(20) => s_sh1_20_port, 
                           mask_sh1(19) => s_sh1_19_port, mask_sh1(18) => 
                           s_sh1_18_port, mask_sh1(17) => s_sh1_17_port, 
                           mask_sh1(16) => s_sh1_16_port, mask_sh1(15) => 
                           s_sh1_15_port, mask_sh1(14) => s_sh1_14_port, 
                           mask_sh1(13) => s_sh1_13_port, mask_sh1(12) => 
                           s_sh1_12_port, mask_sh1(11) => s_sh1_11_port, 
                           mask_sh1(10) => s_sh1_10_port, mask_sh1(9) => 
                           s_sh1_9_port, mask_sh1(8) => s_sh1_8_port, 
                           mask_sh1(7) => s_sh1_7_port, mask_sh1(6) => 
                           s_sh1_6_port, mask_sh1(5) => s_sh1_5_port, 
                           mask_sh1(4) => s_sh1_4_port, mask_sh1(3) => 
                           s_sh1_3_port, mask_sh1(2) => s_sh1_2_port, 
                           mask_sh1(1) => s_sh1_1_port, mask_sh1(0) => 
                           s_sh1_0_port, mask_sh2(31) => s_sh2_31_port, 
                           mask_sh2(30) => s_sh2_30_port, mask_sh2(29) => 
                           s_sh2_29_port, mask_sh2(28) => s_sh2_28_port, 
                           mask_sh2(27) => s_sh2_27_port, mask_sh2(26) => 
                           s_sh2_26_port, mask_sh2(25) => s_sh2_25_port, 
                           mask_sh2(24) => s_sh2_24_port, mask_sh2(23) => 
                           s_sh2_23_port, mask_sh2(22) => s_sh2_22_port, 
                           mask_sh2(21) => s_sh2_21_port, mask_sh2(20) => 
                           s_sh2_20_port, mask_sh2(19) => s_sh2_19_port, 
                           mask_sh2(18) => s_sh2_18_port, mask_sh2(17) => 
                           s_sh2_17_port, mask_sh2(16) => s_sh2_16_port, 
                           mask_sh2(15) => s_sh2_15_port, mask_sh2(14) => 
                           s_sh2_14_port, mask_sh2(13) => s_sh2_13_port, 
                           mask_sh2(12) => s_sh2_12_port, mask_sh2(11) => 
                           s_sh2_11_port, mask_sh2(10) => s_sh2_10_port, 
                           mask_sh2(9) => s_sh2_9_port, mask_sh2(8) => 
                           s_sh2_8_port, mask_sh2(7) => s_sh2_7_port, 
                           mask_sh2(6) => s_sh2_6_port, mask_sh2(5) => 
                           s_sh2_5_port, mask_sh2(4) => s_sh2_4_port, 
                           mask_sh2(3) => s_sh2_3_port, mask_sh2(2) => 
                           s_sh2_2_port, mask_sh2(1) => s_sh2_1_port, 
                           mask_sh2(0) => s_sh2_0_port, mask_sh3(31) => 
                           s_sh3_31_port, mask_sh3(30) => s_sh3_30_port, 
                           mask_sh3(29) => s_sh3_29_port, mask_sh3(28) => 
                           s_sh3_28_port, mask_sh3(27) => s_sh3_27_port, 
                           mask_sh3(26) => s_sh3_26_port, mask_sh3(25) => 
                           s_sh3_25_port, mask_sh3(24) => s_sh3_24_port, 
                           mask_sh3(23) => s_sh3_23_port, mask_sh3(22) => 
                           s_sh3_22_port, mask_sh3(21) => s_sh3_21_port, 
                           mask_sh3(20) => s_sh3_20_port, mask_sh3(19) => 
                           s_sh3_19_port, mask_sh3(18) => s_sh3_18_port, 
                           mask_sh3(17) => s_sh3_17_port, mask_sh3(16) => 
                           s_sh3_16_port, mask_sh3(15) => s_sh3_15_port, 
                           mask_sh3(14) => s_sh3_14_port, mask_sh3(13) => 
                           s_sh3_13_port, mask_sh3(12) => s_sh3_12_port, 
                           mask_sh3(11) => s_sh3_11_port, mask_sh3(10) => 
                           s_sh3_10_port, mask_sh3(9) => s_sh3_9_port, 
                           mask_sh3(8) => s_sh3_8_port, mask_sh3(7) => 
                           s_sh3_7_port, mask_sh3(6) => s_sh3_6_port, 
                           mask_sh3(5) => s_sh3_5_port, mask_sh3(4) => 
                           s_sh3_4_port, mask_sh3(3) => s_sh3_3_port, 
                           mask_sh3(2) => s_sh3_2_port, mask_sh3(1) => 
                           s_sh3_1_port, mask_sh3(0) => s_sh3_0_port, 
                           mask_sh4(31) => s_sh4_31_port, mask_sh4(30) => 
                           s_sh4_30_port, mask_sh4(29) => s_sh4_29_port, 
                           mask_sh4(28) => s_sh4_28_port, mask_sh4(27) => 
                           s_sh4_27_port, mask_sh4(26) => s_sh4_26_port, 
                           mask_sh4(25) => s_sh4_25_port, mask_sh4(24) => 
                           s_sh4_24_port, mask_sh4(23) => s_sh4_23_port, 
                           mask_sh4(22) => s_sh4_22_port, mask_sh4(21) => 
                           s_sh4_21_port, mask_sh4(20) => s_sh4_20_port, 
                           mask_sh4(19) => s_sh4_19_port, mask_sh4(18) => 
                           s_sh4_18_port, mask_sh4(17) => s_sh4_17_port, 
                           mask_sh4(16) => s_sh4_16_port, mask_sh4(15) => 
                           s_sh4_15_port, mask_sh4(14) => s_sh4_14_port, 
                           mask_sh4(13) => s_sh4_13_port, mask_sh4(12) => 
                           s_sh4_12_port, mask_sh4(11) => s_sh4_11_port, 
                           mask_sh4(10) => s_sh4_10_port, mask_sh4(9) => 
                           s_sh4_9_port, mask_sh4(8) => s_sh4_8_port, 
                           mask_sh4(7) => s_sh4_7_port, mask_sh4(6) => 
                           s_sh4_6_port, mask_sh4(5) => s_sh4_5_port, 
                           mask_sh4(4) => s_sh4_4_port, mask_sh4(3) => 
                           s_sh4_3_port, mask_sh4(2) => s_sh4_2_port, 
                           mask_sh4(1) => s_sh4_1_port, mask_sh4(0) => 
                           s_sh4_0_port, mask_sh5(31) => s_sh5_31_port, 
                           mask_sh5(30) => s_sh5_30_port, mask_sh5(29) => 
                           s_sh5_29_port, mask_sh5(28) => s_sh5_28_port, 
                           mask_sh5(27) => s_sh5_27_port, mask_sh5(26) => 
                           s_sh5_26_port, mask_sh5(25) => s_sh5_25_port, 
                           mask_sh5(24) => s_sh5_24_port, mask_sh5(23) => 
                           s_sh5_23_port, mask_sh5(22) => s_sh5_22_port, 
                           mask_sh5(21) => s_sh5_21_port, mask_sh5(20) => 
                           s_sh5_20_port, mask_sh5(19) => s_sh5_19_port, 
                           mask_sh5(18) => s_sh5_18_port, mask_sh5(17) => 
                           s_sh5_17_port, mask_sh5(16) => s_sh5_16_port, 
                           mask_sh5(15) => s_sh5_15_port, mask_sh5(14) => 
                           s_sh5_14_port, mask_sh5(13) => s_sh5_13_port, 
                           mask_sh5(12) => s_sh5_12_port, mask_sh5(11) => 
                           s_sh5_11_port, mask_sh5(10) => s_sh5_10_port, 
                           mask_sh5(9) => s_sh5_9_port, mask_sh5(8) => 
                           s_sh5_8_port, mask_sh5(7) => s_sh5_7_port, 
                           mask_sh5(6) => s_sh5_6_port, mask_sh5(5) => 
                           s_sh5_5_port, mask_sh5(4) => s_sh5_4_port, 
                           mask_sh5(3) => s_sh5_3_port, mask_sh5(2) => 
                           s_sh5_2_port, mask_sh5(1) => s_sh5_1_port, 
                           mask_sh5(0) => s_sh5_0_port, mask_sh6(31) => 
                           s_sh6_31_port, mask_sh6(30) => s_sh6_30_port, 
                           mask_sh6(29) => s_sh6_29_port, mask_sh6(28) => 
                           s_sh6_28_port, mask_sh6(27) => s_sh6_27_port, 
                           mask_sh6(26) => s_sh6_26_port, mask_sh6(25) => 
                           s_sh6_25_port, mask_sh6(24) => s_sh6_24_port, 
                           mask_sh6(23) => s_sh6_23_port, mask_sh6(22) => 
                           s_sh6_22_port, mask_sh6(21) => s_sh6_21_port, 
                           mask_sh6(20) => s_sh6_20_port, mask_sh6(19) => 
                           s_sh6_19_port, mask_sh6(18) => s_sh6_18_port, 
                           mask_sh6(17) => s_sh6_17_port, mask_sh6(16) => 
                           s_sh6_16_port, mask_sh6(15) => s_sh6_15_port, 
                           mask_sh6(14) => s_sh6_14_port, mask_sh6(13) => 
                           s_sh6_13_port, mask_sh6(12) => s_sh6_12_port, 
                           mask_sh6(11) => s_sh6_11_port, mask_sh6(10) => 
                           s_sh6_10_port, mask_sh6(9) => s_sh6_9_port, 
                           mask_sh6(8) => s_sh6_8_port, mask_sh6(7) => 
                           s_sh6_7_port, mask_sh6(6) => s_sh6_6_port, 
                           mask_sh6(5) => s_sh6_5_port, mask_sh6(4) => 
                           s_sh6_4_port, mask_sh6(3) => s_sh6_3_port, 
                           mask_sh6(2) => s_sh6_2_port, mask_sh6(1) => 
                           s_sh6_1_port, mask_sh6(0) => s_sh6_0_port, 
                           mask_sh7(31) => s_sh7_31_port, mask_sh7(30) => 
                           s_sh7_30_port, mask_sh7(29) => s_sh7_29_port, 
                           mask_sh7(28) => s_sh7_28_port, mask_sh7(27) => 
                           s_sh7_27_port, mask_sh7(26) => s_sh7_26_port, 
                           mask_sh7(25) => s_sh7_25_port, mask_sh7(24) => 
                           s_sh7_24_port, mask_sh7(23) => s_sh7_23_port, 
                           mask_sh7(22) => s_sh7_22_port, mask_sh7(21) => 
                           s_sh7_21_port, mask_sh7(20) => s_sh7_20_port, 
                           mask_sh7(19) => s_sh7_19_port, mask_sh7(18) => 
                           s_sh7_18_port, mask_sh7(17) => s_sh7_17_port, 
                           mask_sh7(16) => s_sh7_16_port, mask_sh7(15) => 
                           s_sh7_15_port, mask_sh7(14) => s_sh7_14_port, 
                           mask_sh7(13) => s_sh7_13_port, mask_sh7(12) => 
                           s_sh7_12_port, mask_sh7(11) => s_sh7_11_port, 
                           mask_sh7(10) => s_sh7_10_port, mask_sh7(9) => 
                           s_sh7_9_port, mask_sh7(8) => s_sh7_8_port, 
                           mask_sh7(7) => s_sh7_7_port, mask_sh7(6) => 
                           s_sh7_6_port, mask_sh7(5) => s_sh7_5_port, 
                           mask_sh7(4) => s_sh7_4_port, mask_sh7(3) => 
                           s_sh7_3_port, mask_sh7(2) => s_sh7_2_port, 
                           mask_sh7(1) => s_sh7_1_port, mask_sh7(0) => 
                           s_sh7_0_port);
   MUX_shift_select : MUX81_GENERIC_NBIT32 port map( A(31) => s_sh0_31_port, 
                           A(30) => s_sh0_30_port, A(29) => s_sh0_29_port, 
                           A(28) => s_sh0_28_port, A(27) => s_sh0_27_port, 
                           A(26) => s_sh0_26_port, A(25) => s_sh0_25_port, 
                           A(24) => s_sh0_24_port, A(23) => s_sh0_23_port, 
                           A(22) => s_sh0_22_port, A(21) => s_sh0_21_port, 
                           A(20) => s_sh0_20_port, A(19) => s_sh0_19_port, 
                           A(18) => s_sh0_18_port, A(17) => s_sh0_17_port, 
                           A(16) => s_sh0_16_port, A(15) => s_sh0_15_port, 
                           A(14) => s_sh0_14_port, A(13) => s_sh0_13_port, 
                           A(12) => s_sh0_12_port, A(11) => s_sh0_11_port, 
                           A(10) => s_sh0_10_port, A(9) => s_sh0_9_port, A(8) 
                           => s_sh0_8_port, A(7) => s_sh0_7_port, A(6) => 
                           s_sh0_6_port, A(5) => s_sh0_5_port, A(4) => 
                           s_sh0_4_port, A(3) => s_sh0_3_port, A(2) => 
                           s_sh0_2_port, A(1) => s_sh0_1_port, A(0) => 
                           s_sh0_0_port, B(31) => s_sh1_31_port, B(30) => 
                           s_sh1_30_port, B(29) => s_sh1_29_port, B(28) => 
                           s_sh1_28_port, B(27) => s_sh1_27_port, B(26) => 
                           s_sh1_26_port, B(25) => s_sh1_25_port, B(24) => 
                           s_sh1_24_port, B(23) => s_sh1_23_port, B(22) => 
                           s_sh1_22_port, B(21) => s_sh1_21_port, B(20) => 
                           s_sh1_20_port, B(19) => s_sh1_19_port, B(18) => 
                           s_sh1_18_port, B(17) => s_sh1_17_port, B(16) => 
                           s_sh1_16_port, B(15) => s_sh1_15_port, B(14) => 
                           s_sh1_14_port, B(13) => s_sh1_13_port, B(12) => 
                           s_sh1_12_port, B(11) => s_sh1_11_port, B(10) => 
                           s_sh1_10_port, B(9) => s_sh1_9_port, B(8) => 
                           s_sh1_8_port, B(7) => s_sh1_7_port, B(6) => 
                           s_sh1_6_port, B(5) => s_sh1_5_port, B(4) => 
                           s_sh1_4_port, B(3) => s_sh1_3_port, B(2) => 
                           s_sh1_2_port, B(1) => s_sh1_1_port, B(0) => 
                           s_sh1_0_port, C(31) => s_sh2_31_port, C(30) => 
                           s_sh2_30_port, C(29) => s_sh2_29_port, C(28) => 
                           s_sh2_28_port, C(27) => s_sh2_27_port, C(26) => 
                           s_sh2_26_port, C(25) => s_sh2_25_port, C(24) => 
                           s_sh2_24_port, C(23) => s_sh2_23_port, C(22) => 
                           s_sh2_22_port, C(21) => s_sh2_21_port, C(20) => 
                           s_sh2_20_port, C(19) => s_sh2_19_port, C(18) => 
                           s_sh2_18_port, C(17) => s_sh2_17_port, C(16) => 
                           s_sh2_16_port, C(15) => s_sh2_15_port, C(14) => 
                           s_sh2_14_port, C(13) => s_sh2_13_port, C(12) => 
                           s_sh2_12_port, C(11) => s_sh2_11_port, C(10) => 
                           s_sh2_10_port, C(9) => s_sh2_9_port, C(8) => 
                           s_sh2_8_port, C(7) => s_sh2_7_port, C(6) => 
                           s_sh2_6_port, C(5) => s_sh2_5_port, C(4) => 
                           s_sh2_4_port, C(3) => s_sh2_3_port, C(2) => 
                           s_sh2_2_port, C(1) => s_sh2_1_port, C(0) => 
                           s_sh2_0_port, D(31) => s_sh3_31_port, D(30) => 
                           s_sh3_30_port, D(29) => s_sh3_29_port, D(28) => 
                           s_sh3_28_port, D(27) => s_sh3_27_port, D(26) => 
                           s_sh3_26_port, D(25) => s_sh3_25_port, D(24) => 
                           s_sh3_24_port, D(23) => s_sh3_23_port, D(22) => 
                           s_sh3_22_port, D(21) => s_sh3_21_port, D(20) => 
                           s_sh3_20_port, D(19) => s_sh3_19_port, D(18) => 
                           s_sh3_18_port, D(17) => s_sh3_17_port, D(16) => 
                           s_sh3_16_port, D(15) => s_sh3_15_port, D(14) => 
                           s_sh3_14_port, D(13) => s_sh3_13_port, D(12) => 
                           s_sh3_12_port, D(11) => s_sh3_11_port, D(10) => 
                           s_sh3_10_port, D(9) => s_sh3_9_port, D(8) => 
                           s_sh3_8_port, D(7) => s_sh3_7_port, D(6) => 
                           s_sh3_6_port, D(5) => s_sh3_5_port, D(4) => 
                           s_sh3_4_port, D(3) => s_sh3_3_port, D(2) => 
                           s_sh3_2_port, D(1) => s_sh3_1_port, D(0) => 
                           s_sh3_0_port, E(31) => s_sh4_31_port, E(30) => 
                           s_sh4_30_port, E(29) => s_sh4_29_port, E(28) => 
                           s_sh4_28_port, E(27) => s_sh4_27_port, E(26) => 
                           s_sh4_26_port, E(25) => s_sh4_25_port, E(24) => 
                           s_sh4_24_port, E(23) => s_sh4_23_port, E(22) => 
                           s_sh4_22_port, E(21) => s_sh4_21_port, E(20) => 
                           s_sh4_20_port, E(19) => s_sh4_19_port, E(18) => 
                           s_sh4_18_port, E(17) => s_sh4_17_port, E(16) => 
                           s_sh4_16_port, E(15) => s_sh4_15_port, E(14) => 
                           s_sh4_14_port, E(13) => s_sh4_13_port, E(12) => 
                           s_sh4_12_port, E(11) => s_sh4_11_port, E(10) => 
                           s_sh4_10_port, E(9) => s_sh4_9_port, E(8) => 
                           s_sh4_8_port, E(7) => s_sh4_7_port, E(6) => 
                           s_sh4_6_port, E(5) => s_sh4_5_port, E(4) => 
                           s_sh4_4_port, E(3) => s_sh4_3_port, E(2) => 
                           s_sh4_2_port, E(1) => s_sh4_1_port, E(0) => 
                           s_sh4_0_port, F(31) => s_sh5_31_port, F(30) => 
                           s_sh5_30_port, F(29) => s_sh5_29_port, F(28) => 
                           s_sh5_28_port, F(27) => s_sh5_27_port, F(26) => 
                           s_sh5_26_port, F(25) => s_sh5_25_port, F(24) => 
                           s_sh5_24_port, F(23) => s_sh5_23_port, F(22) => 
                           s_sh5_22_port, F(21) => s_sh5_21_port, F(20) => 
                           s_sh5_20_port, F(19) => s_sh5_19_port, F(18) => 
                           s_sh5_18_port, F(17) => s_sh5_17_port, F(16) => 
                           s_sh5_16_port, F(15) => s_sh5_15_port, F(14) => 
                           s_sh5_14_port, F(13) => s_sh5_13_port, F(12) => 
                           s_sh5_12_port, F(11) => s_sh5_11_port, F(10) => 
                           s_sh5_10_port, F(9) => s_sh5_9_port, F(8) => 
                           s_sh5_8_port, F(7) => s_sh5_7_port, F(6) => 
                           s_sh5_6_port, F(5) => s_sh5_5_port, F(4) => 
                           s_sh5_4_port, F(3) => s_sh5_3_port, F(2) => 
                           s_sh5_2_port, F(1) => s_sh5_1_port, F(0) => 
                           s_sh5_0_port, G(31) => s_sh6_31_port, G(30) => 
                           s_sh6_30_port, G(29) => s_sh6_29_port, G(28) => 
                           s_sh6_28_port, G(27) => s_sh6_27_port, G(26) => 
                           s_sh6_26_port, G(25) => s_sh6_25_port, G(24) => 
                           s_sh6_24_port, G(23) => s_sh6_23_port, G(22) => 
                           s_sh6_22_port, G(21) => s_sh6_21_port, G(20) => 
                           s_sh6_20_port, G(19) => s_sh6_19_port, G(18) => 
                           s_sh6_18_port, G(17) => s_sh6_17_port, G(16) => 
                           s_sh6_16_port, G(15) => s_sh6_15_port, G(14) => 
                           s_sh6_14_port, G(13) => s_sh6_13_port, G(12) => 
                           s_sh6_12_port, G(11) => s_sh6_11_port, G(10) => 
                           s_sh6_10_port, G(9) => s_sh6_9_port, G(8) => 
                           s_sh6_8_port, G(7) => s_sh6_7_port, G(6) => 
                           s_sh6_6_port, G(5) => s_sh6_5_port, G(4) => 
                           s_sh6_4_port, G(3) => s_sh6_3_port, G(2) => 
                           s_sh6_2_port, G(1) => s_sh6_1_port, G(0) => 
                           s_sh6_0_port, H(31) => s_sh7_31_port, H(30) => 
                           s_sh7_30_port, H(29) => s_sh7_29_port, H(28) => 
                           s_sh7_28_port, H(27) => s_sh7_27_port, H(26) => 
                           s_sh7_26_port, H(25) => s_sh7_25_port, H(24) => 
                           s_sh7_24_port, H(23) => s_sh7_23_port, H(22) => 
                           s_sh7_22_port, H(21) => s_sh7_21_port, H(20) => 
                           s_sh7_20_port, H(19) => s_sh7_19_port, H(18) => 
                           s_sh7_18_port, H(17) => s_sh7_17_port, H(16) => 
                           s_sh7_16_port, H(15) => s_sh7_15_port, H(14) => 
                           s_sh7_14_port, H(13) => s_sh7_13_port, H(12) => 
                           s_sh7_12_port, H(11) => s_sh7_11_port, H(10) => 
                           s_sh7_10_port, H(9) => s_sh7_9_port, H(8) => 
                           s_sh7_8_port, H(7) => s_sh7_7_port, H(6) => 
                           s_sh7_6_port, H(5) => s_sh7_5_port, H(4) => 
                           s_sh7_4_port, H(3) => s_sh7_3_port, H(2) => 
                           s_sh7_2_port, H(1) => s_sh7_1_port, H(0) => 
                           s_sh7_0_port, SEL(2) => R2(2), SEL(1) => R2(1), 
                           SEL(0) => R2(0), Y(31) => Rout(31), Y(30) => 
                           Rout(30), Y(29) => Rout(29), Y(28) => Rout(28), 
                           Y(27) => Rout(27), Y(26) => Rout(26), Y(25) => 
                           Rout(25), Y(24) => Rout(24), Y(23) => Rout(23), 
                           Y(22) => Rout(22), Y(21) => Rout(21), Y(20) => 
                           Rout(20), Y(19) => Rout(19), Y(18) => Rout(18), 
                           Y(17) => Rout(17), Y(16) => Rout(16), Y(15) => 
                           Rout(15), Y(14) => Rout(14), Y(13) => Rout(13), 
                           Y(12) => Rout(12), Y(11) => Rout(11), Y(10) => 
                           Rout(10), Y(9) => Rout(9), Y(8) => Rout(8), Y(7) => 
                           Rout(7), Y(6) => Rout(6), Y(5) => Rout(5), Y(4) => 
                           Rout(4), Y(3) => Rout(3), Y(2) => Rout(2), Y(1) => 
                           Rout(1), Y(0) => Rout(0));
   U1 : NOR2_X1 port map( A1 => LnR, A2 => n1, ZN => s_RnS);
   U2 : INV_X1 port map( A => RnS, ZN => n1);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity carry_select_block_n4_0 is

   port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S : 
         out std_logic_vector (3 downto 0));

end carry_select_block_n4_0;

architecture SYN_STRUCTURAL of carry_select_block_n4_0 is

   component MUX21_GENERIC_NBIT4_0
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_127
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_0
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, n_1573, 
      n_1574 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : RCA_GEN_NBIT4_0 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           sum0_3_port, S(2) => sum0_2_port, S(1) => 
                           sum0_1_port, S(0) => sum0_0_port, Co => n_1573);
   RCA1 : RCA_GEN_NBIT4_127 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1),
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           sum1_3_port, S(2) => sum1_2_port, S(1) => 
                           sum1_1_port, S(0) => sum1_0_port, Co => n_1574);
   mux : MUX21_GENERIC_NBIT4_0 port map( A(3) => sum0_3_port, A(2) => 
                           sum0_2_port, A(1) => sum0_1_port, A(0) => 
                           sum0_0_port, B(3) => sum1_3_port, B(2) => 
                           sum1_2_port, B(1) => sum1_1_port, B(0) => 
                           sum1_0_port, SEL => C_sel, Y(3) => S(3), Y(2) => 
                           S(2), Y(1) => S(1), Y(0) => S(0));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity G_BLOCK_0 is

   port( p2, g2, g1 : in std_logic;  G : out std_logic);

end G_BLOCK_0;

architecture SYN_behavioral of G_BLOCK_0 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => G);
   U2 : AOI21_X1 port map( B1 => p2, B2 => g1, A => g2, ZN => n2);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity PG_BLOCK_0 is

   port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);

end PG_BLOCK_0;

architecture SYN_behavioral of PG_BLOCK_0 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => p2, A2 => p1, ZN => PG_P);
   U2 : INV_X1 port map( A => n2, ZN => PG_G);
   U3 : AOI21_X1 port map( B1 => g1, B2 => p2, A => g2, ZN => n2);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity pg_net_0 is

   port( a, b : in std_logic;  p, g : out std_logic);

end pg_net_0;

architecture SYN_behavioral of pg_net_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U2 : XOR2_X1 port map( A => b, B => a, Z => p);
   U1 : AND2_X1 port map( A1 => b, A2 => a, ZN => g);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX51_0 is

   port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0);  
         Y : out std_logic);

end MUX51_0;

architecture SYN_BEHAVIORAL of MUX51_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n7, n8, n1, n2, n3 : std_logic;

begin
   
   U1 : AOI22_X1 port map( A1 => C, A2 => n1, B1 => D, B2 => S(0), ZN => n7);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S(0), B2 => B, ZN => n8);
   U3 : INV_X1 port map( A => n5, ZN => Y);
   U4 : AOI22_X1 port map( A1 => n6, A2 => n3, B1 => S(2), B2 => E, ZN => n5);
   U5 : OAI22_X1 port map( A1 => n7, A2 => n2, B1 => S(1), B2 => n8, ZN => n6);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);
   U8 : INV_X1 port map( A => S(2), ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity boothmul_NBIT_in32 is

   port( A, B : in std_logic_vector (31 downto 0);  mulin_flag, CLK, RST : in 
         std_logic;  MULready : out std_logic;  P : out std_logic_vector (63 
         downto 0));

end boothmul_NBIT_in32;

architecture SYN_structural of boothmul_NBIT_in32 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component P4_ADDER_NBIT64_1
      port( A, B : in std_logic_vector (63 downto 0);  Cin : in std_logic;  S :
            out std_logic_vector (63 downto 0);  Cout, ovf : out std_logic);
   end component;
   
   component P4_ADDER_NBIT64_2
      port( A, B : in std_logic_vector (63 downto 0);  Cin : in std_logic;  S :
            out std_logic_vector (63 downto 0);  Cout, ovf : out std_logic);
   end component;
   
   component mux51_gen_NBIT32_1
      port( A0, A1, A2, A3, A4 : in std_logic_vector (31 downto 0);  SEL : in 
            std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component negate_NBIT32_1
      port( A : in std_logic_vector (31 downto 0);  Y : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component negate_NBIT32_2
      port( A : in std_logic_vector (31 downto 0);  Y : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component shl2_NBIT32_1
      port( A : in std_logic_vector (31 downto 0);  Y : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component shl1_NBIT32_1
      port( A : in std_logic_vector (31 downto 0);  Y : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component P4_ADDER_NBIT64_0
      port( A, B : in std_logic_vector (63 downto 0);  Cin : in std_logic;  S :
            out std_logic_vector (63 downto 0);  Cout, ovf : out std_logic);
   end component;
   
   component mux51_gen_NBIT32_2
      port( A0, A1, A2, A3, A4 : in std_logic_vector (31 downto 0);  SEL : in 
            std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component negate_NBIT32_3
      port( A : in std_logic_vector (31 downto 0);  Y : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component negate_NBIT32_4
      port( A : in std_logic_vector (31 downto 0);  Y : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component shl2_NBIT32_2
      port( A : in std_logic_vector (31 downto 0);  Y : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component shl1_NBIT32_2
      port( A : in std_logic_vector (31 downto 0);  Y : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component mux51_gen_NBIT32_3
      port( A0, A1, A2, A3, A4 : in std_logic_vector (31 downto 0);  SEL : in 
            std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component mux51_gen_NBIT32_0
      port( A0, A1, A2, A3, A4 : in std_logic_vector (31 downto 0);  SEL : in 
            std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component negate_NBIT32_5
      port( A : in std_logic_vector (31 downto 0);  Y : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component negate_NBIT32_6
      port( A : in std_logic_vector (31 downto 0);  Y : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component negate_NBIT32_7
      port( A : in std_logic_vector (31 downto 0);  Y : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component negate_NBIT32_0
      port( A : in std_logic_vector (31 downto 0);  Y : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component shl3_NBIT32
      port( A : in std_logic_vector (31 downto 0);  Y : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component shl2_NBIT32_0
      port( A : in std_logic_vector (31 downto 0);  Y : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component shl1_NBIT32_0
      port( A : in std_logic_vector (31 downto 0);  Y : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component enc33_1
      port( A : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (2 
            downto 0));
   end component;
   
   component enc33_2
      port( A : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (2 
            downto 0));
   end component;
   
   component enc33_3
      port( A : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (2 
            downto 0));
   end component;
   
   component enc33_0
      port( A : in std_logic_vector (2 downto 0);  Y : out std_logic_vector (2 
            downto 0));
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal X_Logic0_port, flag_reg1, mux1_reg1_31_port, mux1_reg1_30_port, 
      mux1_reg1_29_port, mux1_reg1_28_port, mux1_reg1_27_port, 
      mux1_reg1_26_port, mux1_reg1_25_port, mux1_reg1_24_port, 
      mux1_reg1_23_port, mux1_reg1_22_port, mux1_reg1_21_port, 
      mux1_reg1_20_port, mux1_reg1_19_port, mux1_reg1_18_port, 
      mux1_reg1_17_port, mux1_reg1_16_port, mux1_reg1_15_port, 
      mux1_reg1_14_port, mux1_reg1_13_port, mux1_reg1_12_port, 
      mux1_reg1_11_port, mux1_reg1_10_port, mux1_reg1_9_port, mux1_reg1_8_port,
      mux1_reg1_7_port, mux1_reg1_6_port, mux1_reg1_5_port, mux1_reg1_4_port, 
      mux1_reg1_3_port, mux1_reg1_2_port, mux1_reg1_1_port, mux1_reg1_0_port, 
      mux2_reg1_31_port, mux2_reg1_30_port, mux2_reg1_29_port, 
      mux2_reg1_28_port, mux2_reg1_27_port, mux2_reg1_26_port, 
      mux2_reg1_25_port, mux2_reg1_24_port, mux2_reg1_23_port, 
      mux2_reg1_22_port, mux2_reg1_21_port, mux2_reg1_20_port, 
      mux2_reg1_19_port, mux2_reg1_18_port, mux2_reg1_17_port, 
      mux2_reg1_16_port, mux2_reg1_15_port, mux2_reg1_14_port, 
      mux2_reg1_13_port, mux2_reg1_12_port, mux2_reg1_11_port, 
      mux2_reg1_10_port, mux2_reg1_9_port, mux2_reg1_8_port, mux2_reg1_7_port, 
      mux2_reg1_6_port, mux2_reg1_5_port, mux2_reg1_4_port, mux2_reg1_3_port, 
      mux2_reg1_2_port, mux2_reg1_1_port, mux2_reg1_0_port, A4_reg1_31_port, 
      A4_reg1_30_port, A4_reg1_29_port, A4_reg1_28_port, A4_reg1_27_port, 
      A4_reg1_26_port, A4_reg1_25_port, A4_reg1_24_port, A4_reg1_23_port, 
      A4_reg1_22_port, A4_reg1_21_port, A4_reg1_20_port, A4_reg1_19_port, 
      A4_reg1_18_port, A4_reg1_17_port, A4_reg1_16_port, A4_reg1_15_port, 
      A4_reg1_14_port, A4_reg1_13_port, A4_reg1_12_port, A4_reg1_11_port, 
      A4_reg1_10_port, A4_reg1_9_port, A4_reg1_8_port, A4_reg1_7_port, 
      A4_reg1_6_port, A4_reg1_5_port, A4_reg1_4_port, A4_reg1_3_port, 
      A4_reg1_2_port, A4_reg1_1_port, A4_reg1_0_port, flag_reg2, 
      mux_reg2_31_port, mux_reg2_30_port, mux_reg2_29_port, mux_reg2_28_port, 
      mux_reg2_27_port, mux_reg2_26_port, mux_reg2_25_port, mux_reg2_24_port, 
      mux_reg2_23_port, mux_reg2_22_port, mux_reg2_21_port, mux_reg2_20_port, 
      mux_reg2_19_port, mux_reg2_18_port, mux_reg2_17_port, mux_reg2_16_port, 
      mux_reg2_15_port, mux_reg2_14_port, mux_reg2_13_port, mux_reg2_12_port, 
      mux_reg2_11_port, mux_reg2_10_port, mux_reg2_9_port, mux_reg2_8_port, 
      mux_reg2_7_port, mux_reg2_6_port, mux_reg2_5_port, mux_reg2_4_port, 
      mux_reg2_3_port, mux_reg2_2_port, mux_reg2_1_port, mux_reg2_0_port, 
      sum_reg2_63_port, sum_reg2_62_port, sum_reg2_61_port, sum_reg2_60_port, 
      sum_reg2_59_port, sum_reg2_58_port, sum_reg2_57_port, sum_reg2_56_port, 
      sum_reg2_55_port, sum_reg2_54_port, sum_reg2_53_port, sum_reg2_52_port, 
      sum_reg2_51_port, sum_reg2_50_port, sum_reg2_49_port, sum_reg2_48_port, 
      sum_reg2_47_port, sum_reg2_46_port, sum_reg2_45_port, sum_reg2_44_port, 
      sum_reg2_43_port, sum_reg2_42_port, sum_reg2_41_port, sum_reg2_40_port, 
      sum_reg2_39_port, sum_reg2_38_port, sum_reg2_37_port, sum_reg2_36_port, 
      sum_reg2_35_port, sum_reg2_34_port, sum_reg2_33_port, sum_reg2_32_port, 
      sum_reg2_31_port, sum_reg2_30_port, sum_reg2_29_port, sum_reg2_28_port, 
      sum_reg2_27_port, sum_reg2_26_port, sum_reg2_25_port, sum_reg2_24_port, 
      sum_reg2_23_port, sum_reg2_22_port, sum_reg2_21_port, sum_reg2_20_port, 
      sum_reg2_19_port, sum_reg2_18_port, sum_reg2_17_port, sum_reg2_16_port, 
      sum_reg2_15_port, sum_reg2_14_port, sum_reg2_13_port, sum_reg2_12_port, 
      sum_reg2_11_port, sum_reg2_10_port, sum_reg2_9_port, sum_reg2_8_port, 
      sum_reg2_7_port, sum_reg2_6_port, sum_reg2_5_port, sum_reg2_4_port, 
      sum_reg2_3_port, sum_reg2_2_port, sum_reg2_1_port, sum_reg2_0_port, 
      A4_reg2_31_port, A4_reg2_30_port, A4_reg2_29_port, A4_reg2_28_port, 
      A4_reg2_27_port, A4_reg2_26_port, A4_reg2_25_port, A4_reg2_24_port, 
      A4_reg2_23_port, A4_reg2_22_port, A4_reg2_21_port, A4_reg2_20_port, 
      A4_reg2_19_port, A4_reg2_18_port, A4_reg2_17_port, A4_reg2_16_port, 
      A4_reg2_15_port, A4_reg2_14_port, A4_reg2_13_port, A4_reg2_12_port, 
      A4_reg2_11_port, A4_reg2_10_port, A4_reg2_9_port, A4_reg2_8_port, 
      A4_reg2_7_port, A4_reg2_6_port, A4_reg2_5_port, A4_reg2_4_port, 
      A4_reg2_3_port, A4_reg2_2_port, A4_reg2_1_port, A4_reg2_0_port, 
      mux_reg3_31_port, mux_reg3_30_port, mux_reg3_29_port, mux_reg3_28_port, 
      mux_reg3_27_port, mux_reg3_26_port, mux_reg3_25_port, mux_reg3_24_port, 
      mux_reg3_23_port, mux_reg3_22_port, mux_reg3_21_port, mux_reg3_20_port, 
      mux_reg3_19_port, mux_reg3_18_port, mux_reg3_17_port, mux_reg3_16_port, 
      mux_reg3_15_port, mux_reg3_14_port, mux_reg3_13_port, mux_reg3_12_port, 
      mux_reg3_11_port, mux_reg3_10_port, mux_reg3_9_port, mux_reg3_8_port, 
      mux_reg3_7_port, mux_reg3_6_port, mux_reg3_5_port, mux_reg3_4_port, 
      mux_reg3_3_port, mux_reg3_2_port, mux_reg3_1_port, mux_reg3_0_port, 
      sum_reg3_63_port, sum_reg3_62_port, sum_reg3_61_port, sum_reg3_60_port, 
      sum_reg3_59_port, sum_reg3_58_port, sum_reg3_57_port, sum_reg3_56_port, 
      sum_reg3_55_port, sum_reg3_54_port, sum_reg3_53_port, sum_reg3_52_port, 
      sum_reg3_51_port, sum_reg3_50_port, sum_reg3_49_port, sum_reg3_48_port, 
      sum_reg3_47_port, sum_reg3_46_port, sum_reg3_45_port, sum_reg3_44_port, 
      sum_reg3_43_port, sum_reg3_42_port, sum_reg3_41_port, sum_reg3_40_port, 
      sum_reg3_39_port, sum_reg3_38_port, sum_reg3_37_port, sum_reg3_36_port, 
      sum_reg3_35_port, sum_reg3_34_port, sum_reg3_33_port, sum_reg3_32_port, 
      sum_reg3_31_port, sum_reg3_30_port, sum_reg3_29_port, sum_reg3_28_port, 
      sum_reg3_27_port, sum_reg3_26_port, sum_reg3_25_port, sum_reg3_24_port, 
      sum_reg3_23_port, sum_reg3_22_port, sum_reg3_21_port, sum_reg3_20_port, 
      sum_reg3_19_port, sum_reg3_18_port, sum_reg3_17_port, sum_reg3_16_port, 
      sum_reg3_15_port, sum_reg3_14_port, sum_reg3_13_port, sum_reg3_12_port, 
      sum_reg3_11_port, sum_reg3_10_port, sum_reg3_9_port, sum_reg3_8_port, 
      sum_reg3_7_port, sum_reg3_6_port, sum_reg3_5_port, sum_reg3_4_port, 
      sum_reg3_3_port, sum_reg3_2_port, sum_reg3_1_port, sum_reg3_0_port, 
      enc_reg21_2_port, enc_reg21_1_port, enc_reg21_0_port, enc_reg31_2_port, 
      enc_reg31_1_port, enc_reg31_0_port, enc_reg32_2_port, enc_reg32_1_port, 
      enc_reg32_0_port, mux1_out_31_port, mux1_out_30_port, mux1_out_29_port, 
      mux1_out_28_port, mux1_out_27_port, mux1_out_26_port, mux1_out_25_port, 
      mux1_out_24_port, mux1_out_23_port, mux1_out_22_port, mux1_out_21_port, 
      mux1_out_20_port, mux1_out_19_port, mux1_out_18_port, mux1_out_17_port, 
      mux1_out_16_port, mux1_out_15_port, mux1_out_14_port, mux1_out_13_port, 
      mux1_out_12_port, mux1_out_11_port, mux1_out_10_port, mux1_out_9_port, 
      mux1_out_8_port, mux1_out_7_port, mux1_out_6_port, mux1_out_5_port, 
      mux1_out_4_port, mux1_out_3_port, mux1_out_2_port, mux1_out_1_port, 
      mux1_out_0_port, mux2_out_31_port, mux2_out_30_port, mux2_out_29_port, 
      mux2_out_28_port, mux2_out_27_port, mux2_out_26_port, mux2_out_25_port, 
      mux2_out_24_port, mux2_out_23_port, mux2_out_22_port, mux2_out_21_port, 
      mux2_out_20_port, mux2_out_19_port, mux2_out_18_port, mux2_out_17_port, 
      mux2_out_16_port, mux2_out_15_port, mux2_out_14_port, mux2_out_13_port, 
      mux2_out_12_port, mux2_out_11_port, mux2_out_10_port, mux2_out_9_port, 
      mux2_out_8_port, mux2_out_7_port, mux2_out_6_port, mux2_out_5_port, 
      mux2_out_4_port, mux2_out_3_port, mux2_out_2_port, mux2_out_1_port, 
      mux2_out_0_port, s_8A_1_31_port, s_8A_1_30_port, s_8A_1_29_port, 
      s_8A_1_28_port, s_8A_1_27_port, s_8A_1_26_port, s_8A_1_25_port, 
      s_8A_1_24_port, s_8A_1_23_port, s_8A_1_22_port, s_8A_1_21_port, 
      s_8A_1_20_port, s_8A_1_19_port, s_8A_1_18_port, s_8A_1_17_port, 
      s_8A_1_16_port, s_8A_1_15_port, s_8A_1_14_port, s_8A_1_13_port, 
      s_8A_1_12_port, s_8A_1_11_port, s_8A_1_10_port, s_8A_1_9_port, 
      s_8A_1_8_port, s_8A_1_7_port, s_8A_1_6_port, s_8A_1_5_port, s_8A_1_4_port
      , s_8A_1_3_port, s_8A_1_2_port, s_8A_1_1_port, s_8A_1_0_port, 
      mux_2_out_31_port, mux_2_out_30_port, mux_2_out_29_port, 
      mux_2_out_28_port, mux_2_out_27_port, mux_2_out_26_port, 
      mux_2_out_25_port, mux_2_out_24_port, mux_2_out_23_port, 
      mux_2_out_22_port, mux_2_out_21_port, mux_2_out_20_port, 
      mux_2_out_19_port, mux_2_out_18_port, mux_2_out_17_port, 
      mux_2_out_16_port, mux_2_out_15_port, mux_2_out_14_port, 
      mux_2_out_13_port, mux_2_out_12_port, mux_2_out_11_port, 
      mux_2_out_10_port, mux_2_out_9_port, mux_2_out_8_port, mux_2_out_7_port, 
      mux_2_out_6_port, mux_2_out_5_port, mux_2_out_4_port, mux_2_out_3_port, 
      mux_2_out_2_port, mux_2_out_1_port, mux_2_out_0_port, sum_2_out_63_port, 
      sum_2_out_62_port, sum_2_out_61_port, sum_2_out_60_port, 
      sum_2_out_59_port, sum_2_out_58_port, sum_2_out_57_port, 
      sum_2_out_56_port, sum_2_out_55_port, sum_2_out_54_port, 
      sum_2_out_53_port, sum_2_out_52_port, sum_2_out_51_port, 
      sum_2_out_50_port, sum_2_out_49_port, sum_2_out_48_port, 
      sum_2_out_47_port, sum_2_out_46_port, sum_2_out_45_port, 
      sum_2_out_44_port, sum_2_out_43_port, sum_2_out_42_port, 
      sum_2_out_41_port, sum_2_out_40_port, sum_2_out_39_port, 
      sum_2_out_38_port, sum_2_out_37_port, sum_2_out_36_port, 
      sum_2_out_35_port, sum_2_out_34_port, sum_2_out_33_port, 
      sum_2_out_32_port, sum_2_out_31_port, sum_2_out_30_port, 
      sum_2_out_29_port, sum_2_out_28_port, sum_2_out_27_port, 
      sum_2_out_26_port, sum_2_out_25_port, sum_2_out_24_port, 
      sum_2_out_23_port, sum_2_out_22_port, sum_2_out_21_port, 
      sum_2_out_20_port, sum_2_out_19_port, sum_2_out_18_port, 
      sum_2_out_17_port, sum_2_out_16_port, sum_2_out_15_port, 
      sum_2_out_14_port, sum_2_out_13_port, sum_2_out_12_port, 
      sum_2_out_11_port, sum_2_out_10_port, sum_2_out_9_port, sum_2_out_8_port,
      sum_2_out_7_port, sum_2_out_6_port, sum_2_out_5_port, sum_2_out_4_port, 
      sum_2_out_3_port, sum_2_out_2_port, sum_2_out_1_port, sum_2_out_0_port, 
      s_2A_2_31_port, s_2A_2_30_port, s_2A_2_29_port, s_2A_2_28_port, 
      s_2A_2_27_port, s_2A_2_26_port, s_2A_2_25_port, s_2A_2_24_port, 
      s_2A_2_23_port, s_2A_2_22_port, s_2A_2_21_port, s_2A_2_20_port, 
      s_2A_2_19_port, s_2A_2_18_port, s_2A_2_17_port, s_2A_2_16_port, 
      s_2A_2_15_port, s_2A_2_14_port, s_2A_2_13_port, s_2A_2_12_port, 
      s_2A_2_11_port, s_2A_2_10_port, s_2A_2_9_port, s_2A_2_8_port, 
      s_2A_2_7_port, s_2A_2_6_port, s_2A_2_5_port, s_2A_2_4_port, s_2A_2_3_port
      , s_2A_2_2_port, s_2A_2_1_port, s_2A_2_0_port, mux_3_out_31_port, 
      mux_3_out_30_port, mux_3_out_29_port, mux_3_out_28_port, 
      mux_3_out_27_port, mux_3_out_26_port, mux_3_out_25_port, 
      mux_3_out_24_port, mux_3_out_23_port, mux_3_out_22_port, 
      mux_3_out_21_port, mux_3_out_20_port, mux_3_out_19_port, 
      mux_3_out_18_port, mux_3_out_17_port, mux_3_out_16_port, 
      mux_3_out_15_port, mux_3_out_14_port, mux_3_out_13_port, 
      mux_3_out_12_port, mux_3_out_11_port, mux_3_out_10_port, mux_3_out_9_port
      , mux_3_out_8_port, mux_3_out_7_port, mux_3_out_6_port, mux_3_out_5_port,
      mux_3_out_4_port, mux_3_out_3_port, mux_3_out_2_port, mux_3_out_1_port, 
      mux_3_out_0_port, sum_3_out_63_port, sum_3_out_62_port, sum_3_out_61_port
      , sum_3_out_60_port, sum_3_out_59_port, sum_3_out_58_port, 
      sum_3_out_57_port, sum_3_out_56_port, sum_3_out_55_port, 
      sum_3_out_54_port, sum_3_out_53_port, sum_3_out_52_port, 
      sum_3_out_51_port, sum_3_out_50_port, sum_3_out_49_port, 
      sum_3_out_48_port, sum_3_out_47_port, sum_3_out_46_port, 
      sum_3_out_45_port, sum_3_out_44_port, sum_3_out_43_port, 
      sum_3_out_42_port, sum_3_out_41_port, sum_3_out_40_port, 
      sum_3_out_39_port, sum_3_out_38_port, sum_3_out_37_port, 
      sum_3_out_36_port, sum_3_out_35_port, sum_3_out_34_port, 
      sum_3_out_33_port, sum_3_out_32_port, sum_3_out_31_port, 
      sum_3_out_30_port, sum_3_out_29_port, sum_3_out_28_port, 
      sum_3_out_27_port, sum_3_out_26_port, sum_3_out_25_port, 
      sum_3_out_24_port, sum_3_out_23_port, sum_3_out_22_port, 
      sum_3_out_21_port, sum_3_out_20_port, sum_3_out_19_port, 
      sum_3_out_18_port, sum_3_out_17_port, sum_3_out_16_port, 
      sum_3_out_15_port, sum_3_out_14_port, sum_3_out_13_port, 
      sum_3_out_12_port, sum_3_out_11_port, sum_3_out_10_port, sum_3_out_9_port
      , sum_3_out_8_port, sum_3_out_7_port, sum_3_out_6_port, sum_3_out_5_port,
      sum_3_out_4_port, sum_3_out_3_port, sum_3_out_2_port, sum_3_out_1_port, 
      sum_3_out_0_port, s_sel_3_2_port, s_sel_3_1_port, s_sel_3_0_port, 
      s_sel_2_2_port, s_sel_2_1_port, s_sel_2_0_port, s_sel_1_2_port, 
      s_sel_1_1_port, s_sel_1_0_port, s_sel_0_2_port, s_sel_0_1_port, 
      s_sel_0_0_port, s_2A_1_31_port, s_2A_1_30_port, s_2A_1_29_port, 
      s_2A_1_28_port, s_2A_1_27_port, s_2A_1_26_port, s_2A_1_25_port, 
      s_2A_1_24_port, s_2A_1_23_port, s_2A_1_22_port, s_2A_1_21_port, 
      s_2A_1_20_port, s_2A_1_19_port, s_2A_1_18_port, s_2A_1_17_port, 
      s_2A_1_16_port, s_2A_1_15_port, s_2A_1_14_port, s_2A_1_13_port, 
      s_2A_1_12_port, s_2A_1_11_port, s_2A_1_10_port, s_2A_1_9_port, 
      s_2A_1_8_port, s_2A_1_7_port, s_2A_1_6_port, s_2A_1_5_port, s_2A_1_4_port
      , s_2A_1_3_port, s_2A_1_2_port, s_2A_1_1_port, s_2A_1_0_port, 
      s_4A_1_31_port, s_4A_1_30_port, s_4A_1_29_port, s_4A_1_28_port, 
      s_4A_1_27_port, s_4A_1_26_port, s_4A_1_25_port, s_4A_1_24_port, 
      s_4A_1_23_port, s_4A_1_22_port, s_4A_1_21_port, s_4A_1_20_port, 
      s_4A_1_19_port, s_4A_1_18_port, s_4A_1_17_port, s_4A_1_16_port, 
      s_4A_1_15_port, s_4A_1_14_port, s_4A_1_13_port, s_4A_1_12_port, 
      s_4A_1_11_port, s_4A_1_10_port, s_4A_1_9_port, s_4A_1_8_port, 
      s_4A_1_7_port, s_4A_1_6_port, s_4A_1_5_port, s_4A_1_4_port, s_4A_1_3_port
      , s_4A_1_2_port, s_4A_1_1_port, s_4A_1_0_port, s_A_neg_31_port, 
      s_A_neg_30_port, s_A_neg_29_port, s_A_neg_28_port, s_A_neg_27_port, 
      s_A_neg_26_port, s_A_neg_25_port, s_A_neg_24_port, s_A_neg_23_port, 
      s_A_neg_22_port, s_A_neg_21_port, s_A_neg_20_port, s_A_neg_19_port, 
      s_A_neg_18_port, s_A_neg_17_port, s_A_neg_16_port, s_A_neg_15_port, 
      s_A_neg_14_port, s_A_neg_13_port, s_A_neg_12_port, s_A_neg_11_port, 
      s_A_neg_10_port, s_A_neg_9_port, s_A_neg_8_port, s_A_neg_7_port, 
      s_A_neg_6_port, s_A_neg_5_port, s_A_neg_4_port, s_A_neg_3_port, 
      s_A_neg_2_port, s_A_neg_1_port, s_A_neg_0_port, s_2A_1_neg_31_port, 
      s_2A_1_neg_30_port, s_2A_1_neg_29_port, s_2A_1_neg_28_port, 
      s_2A_1_neg_27_port, s_2A_1_neg_26_port, s_2A_1_neg_25_port, 
      s_2A_1_neg_24_port, s_2A_1_neg_23_port, s_2A_1_neg_22_port, 
      s_2A_1_neg_21_port, s_2A_1_neg_20_port, s_2A_1_neg_19_port, 
      s_2A_1_neg_18_port, s_2A_1_neg_17_port, s_2A_1_neg_16_port, 
      s_2A_1_neg_15_port, s_2A_1_neg_14_port, s_2A_1_neg_13_port, 
      s_2A_1_neg_12_port, s_2A_1_neg_11_port, s_2A_1_neg_10_port, 
      s_2A_1_neg_9_port, s_2A_1_neg_8_port, s_2A_1_neg_7_port, 
      s_2A_1_neg_6_port, s_2A_1_neg_5_port, s_2A_1_neg_4_port, 
      s_2A_1_neg_3_port, s_2A_1_neg_2_port, s_2A_1_neg_1_port, 
      s_2A_1_neg_0_port, s_4A_1_neg_31_port, s_4A_1_neg_30_port, 
      s_4A_1_neg_29_port, s_4A_1_neg_28_port, s_4A_1_neg_27_port, 
      s_4A_1_neg_26_port, s_4A_1_neg_25_port, s_4A_1_neg_24_port, 
      s_4A_1_neg_23_port, s_4A_1_neg_22_port, s_4A_1_neg_21_port, 
      s_4A_1_neg_20_port, s_4A_1_neg_19_port, s_4A_1_neg_18_port, 
      s_4A_1_neg_17_port, s_4A_1_neg_16_port, s_4A_1_neg_15_port, 
      s_4A_1_neg_14_port, s_4A_1_neg_13_port, s_4A_1_neg_12_port, 
      s_4A_1_neg_11_port, s_4A_1_neg_10_port, s_4A_1_neg_9_port, 
      s_4A_1_neg_8_port, s_4A_1_neg_7_port, s_4A_1_neg_6_port, 
      s_4A_1_neg_5_port, s_4A_1_neg_4_port, s_4A_1_neg_3_port, 
      s_4A_1_neg_2_port, s_4A_1_neg_1_port, s_4A_1_neg_0_port, 
      s_8A_1_neg_31_port, s_8A_1_neg_30_port, s_8A_1_neg_29_port, 
      s_8A_1_neg_28_port, s_8A_1_neg_27_port, s_8A_1_neg_26_port, 
      s_8A_1_neg_25_port, s_8A_1_neg_24_port, s_8A_1_neg_23_port, 
      s_8A_1_neg_22_port, s_8A_1_neg_21_port, s_8A_1_neg_20_port, 
      s_8A_1_neg_19_port, s_8A_1_neg_18_port, s_8A_1_neg_17_port, 
      s_8A_1_neg_16_port, s_8A_1_neg_15_port, s_8A_1_neg_14_port, 
      s_8A_1_neg_13_port, s_8A_1_neg_12_port, s_8A_1_neg_11_port, 
      s_8A_1_neg_10_port, s_8A_1_neg_9_port, s_8A_1_neg_8_port, 
      s_8A_1_neg_7_port, s_8A_1_neg_6_port, s_8A_1_neg_5_port, 
      s_8A_1_neg_4_port, s_8A_1_neg_3_port, s_8A_1_neg_2_port, 
      s_8A_1_neg_1_port, s_8A_1_neg_0_port, s_A_2_31_port, s_A_2_30_port, 
      s_A_2_29_port, s_A_2_28_port, s_A_2_27_port, s_A_2_26_port, s_A_2_25_port
      , s_A_2_24_port, s_A_2_23_port, s_A_2_22_port, s_A_2_21_port, 
      s_A_2_20_port, s_A_2_19_port, s_A_2_18_port, s_A_2_17_port, s_A_2_16_port
      , s_A_2_15_port, s_A_2_14_port, s_A_2_13_port, s_A_2_12_port, 
      s_A_2_11_port, s_A_2_10_port, s_A_2_9_port, s_A_2_8_port, s_A_2_7_port, 
      s_A_2_6_port, s_A_2_5_port, s_A_2_4_port, s_A_2_3_port, s_A_2_2_port, 
      s_A_2_1_port, s_A_2_0_port, s_A_2_neg_31_port, s_A_2_neg_30_port, 
      s_A_2_neg_29_port, s_A_2_neg_28_port, s_A_2_neg_27_port, 
      s_A_2_neg_26_port, s_A_2_neg_25_port, s_A_2_neg_24_port, 
      s_A_2_neg_23_port, s_A_2_neg_22_port, s_A_2_neg_21_port, 
      s_A_2_neg_20_port, s_A_2_neg_19_port, s_A_2_neg_18_port, 
      s_A_2_neg_17_port, s_A_2_neg_16_port, s_A_2_neg_15_port, 
      s_A_2_neg_14_port, s_A_2_neg_13_port, s_A_2_neg_12_port, 
      s_A_2_neg_11_port, s_A_2_neg_10_port, s_A_2_neg_9_port, s_A_2_neg_8_port,
      s_A_2_neg_7_port, s_A_2_neg_6_port, s_A_2_neg_5_port, s_A_2_neg_4_port, 
      s_A_2_neg_3_port, s_A_2_neg_2_port, s_A_2_neg_1_port, s_A_2_neg_0_port, 
      s_2A_2_neg_31_port, s_2A_2_neg_30_port, s_2A_2_neg_29_port, 
      s_2A_2_neg_28_port, s_2A_2_neg_27_port, s_2A_2_neg_26_port, 
      s_2A_2_neg_25_port, s_2A_2_neg_24_port, s_2A_2_neg_23_port, 
      s_2A_2_neg_22_port, s_2A_2_neg_21_port, s_2A_2_neg_20_port, 
      s_2A_2_neg_19_port, s_2A_2_neg_18_port, s_2A_2_neg_17_port, 
      s_2A_2_neg_16_port, s_2A_2_neg_15_port, s_2A_2_neg_14_port, 
      s_2A_2_neg_13_port, s_2A_2_neg_12_port, s_2A_2_neg_11_port, 
      s_2A_2_neg_10_port, s_2A_2_neg_9_port, s_2A_2_neg_8_port, 
      s_2A_2_neg_7_port, s_2A_2_neg_6_port, s_2A_2_neg_5_port, 
      s_2A_2_neg_4_port, s_2A_2_neg_3_port, s_2A_2_neg_2_port, 
      s_2A_2_neg_1_port, s_2A_2_neg_0_port, s_A_3_31_port, s_A_3_30_port, 
      s_A_3_29_port, s_A_3_28_port, s_A_3_27_port, s_A_3_26_port, s_A_3_25_port
      , s_A_3_24_port, s_A_3_23_port, s_A_3_22_port, s_A_3_21_port, 
      s_A_3_20_port, s_A_3_19_port, s_A_3_18_port, s_A_3_17_port, s_A_3_16_port
      , s_A_3_15_port, s_A_3_14_port, s_A_3_13_port, s_A_3_12_port, 
      s_A_3_11_port, s_A_3_10_port, s_A_3_9_port, s_A_3_8_port, s_A_3_7_port, 
      s_A_3_6_port, s_A_3_5_port, s_A_3_4_port, s_A_3_3_port, s_A_3_2_port, 
      s_A_3_1_port, s_A_3_0_port, s_2A_3_31_port, s_2A_3_30_port, 
      s_2A_3_29_port, s_2A_3_28_port, s_2A_3_27_port, s_2A_3_26_port, 
      s_2A_3_25_port, s_2A_3_24_port, s_2A_3_23_port, s_2A_3_22_port, 
      s_2A_3_21_port, s_2A_3_20_port, s_2A_3_19_port, s_2A_3_18_port, 
      s_2A_3_17_port, s_2A_3_16_port, s_2A_3_15_port, s_2A_3_14_port, 
      s_2A_3_13_port, s_2A_3_12_port, s_2A_3_11_port, s_2A_3_10_port, 
      s_2A_3_9_port, s_2A_3_8_port, s_2A_3_7_port, s_2A_3_6_port, s_2A_3_5_port
      , s_2A_3_4_port, s_2A_3_3_port, s_2A_3_2_port, s_2A_3_1_port, 
      s_2A_3_0_port, s_A_3_neg_31_port, s_A_3_neg_30_port, s_A_3_neg_29_port, 
      s_A_3_neg_28_port, s_A_3_neg_27_port, s_A_3_neg_26_port, 
      s_A_3_neg_25_port, s_A_3_neg_24_port, s_A_3_neg_23_port, 
      s_A_3_neg_22_port, s_A_3_neg_21_port, s_A_3_neg_20_port, 
      s_A_3_neg_19_port, s_A_3_neg_18_port, s_A_3_neg_17_port, 
      s_A_3_neg_16_port, s_A_3_neg_15_port, s_A_3_neg_14_port, 
      s_A_3_neg_13_port, s_A_3_neg_12_port, s_A_3_neg_11_port, 
      s_A_3_neg_10_port, s_A_3_neg_9_port, s_A_3_neg_8_port, s_A_3_neg_7_port, 
      s_A_3_neg_6_port, s_A_3_neg_5_port, s_A_3_neg_4_port, s_A_3_neg_3_port, 
      s_A_3_neg_2_port, s_A_3_neg_1_port, s_A_3_neg_0_port, s_2A_3_neg_31_port,
      s_2A_3_neg_30_port, s_2A_3_neg_29_port, s_2A_3_neg_28_port, 
      s_2A_3_neg_27_port, s_2A_3_neg_26_port, s_2A_3_neg_25_port, 
      s_2A_3_neg_24_port, s_2A_3_neg_23_port, s_2A_3_neg_22_port, 
      s_2A_3_neg_21_port, s_2A_3_neg_20_port, s_2A_3_neg_19_port, 
      s_2A_3_neg_18_port, s_2A_3_neg_17_port, s_2A_3_neg_16_port, 
      s_2A_3_neg_15_port, s_2A_3_neg_14_port, s_2A_3_neg_13_port, 
      s_2A_3_neg_12_port, s_2A_3_neg_11_port, s_2A_3_neg_10_port, 
      s_2A_3_neg_9_port, s_2A_3_neg_8_port, s_2A_3_neg_7_port, 
      s_2A_3_neg_6_port, s_2A_3_neg_5_port, s_2A_3_neg_4_port, 
      s_2A_3_neg_3_port, s_2A_3_neg_2_port, s_2A_3_neg_1_port, 
      s_2A_3_neg_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13
      , n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, 
      n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42
      , n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, 
      n57, n58, n59, n60, n_1575, n_1576, n_1577, n_1578, n_1579, n_1580, 
      n_1581, n_1582, n_1583, n_1584, n_1585, n_1586, n_1587, n_1588, n_1589, 
      n_1590, n_1591, n_1592, n_1593, n_1594, n_1595, n_1596, n_1597, n_1598, 
      n_1599, n_1600, n_1601, n_1602, n_1603, n_1604, n_1605, n_1606, n_1607, 
      n_1608, n_1609, n_1610, n_1611, n_1612, n_1613, n_1614, n_1615, n_1616, 
      n_1617, n_1618, n_1619, n_1620, n_1621, n_1622, n_1623, n_1624, n_1625, 
      n_1626, n_1627, n_1628, n_1629, n_1630, n_1631, n_1632, n_1633, n_1634, 
      n_1635, n_1636, n_1637, n_1638, n_1639, n_1640, n_1641, n_1642, n_1643, 
      n_1644, n_1645, n_1646, n_1647, n_1648, n_1649, n_1650, n_1651, n_1652, 
      n_1653, n_1654, n_1655, n_1656, n_1657, n_1658, n_1659, n_1660, n_1661, 
      n_1662, n_1663, n_1664, n_1665, n_1666, n_1667, n_1668, n_1669, n_1670, 
      n_1671, n_1672, n_1673, n_1674, n_1675, n_1676, n_1677, n_1678, n_1679, 
      n_1680, n_1681, n_1682, n_1683, n_1684, n_1685, n_1686, n_1687, n_1688, 
      n_1689, n_1690, n_1691, n_1692, n_1693, n_1694, n_1695, n_1696, n_1697, 
      n_1698, n_1699, n_1700, n_1701, n_1702, n_1703, n_1704, n_1705, n_1706, 
      n_1707, n_1708, n_1709, n_1710, n_1711, n_1712, n_1713, n_1714, n_1715, 
      n_1716, n_1717, n_1718, n_1719, n_1720, n_1721, n_1722, n_1723, n_1724, 
      n_1725, n_1726, n_1727, n_1728, n_1729, n_1730, n_1731, n_1732, n_1733, 
      n_1734, n_1735, n_1736, n_1737, n_1738, n_1739, n_1740, n_1741, n_1742, 
      n_1743, n_1744, n_1745, n_1746, n_1747, n_1748, n_1749, n_1750, n_1751, 
      n_1752, n_1753, n_1754, n_1755, n_1756, n_1757, n_1758, n_1759, n_1760, 
      n_1761, n_1762, n_1763, n_1764, n_1765, n_1766, n_1767, n_1768, n_1769, 
      n_1770, n_1771, n_1772, n_1773, n_1774, n_1775, n_1776, n_1777, n_1778, 
      n_1779, n_1780, n_1781, n_1782, n_1783, n_1784, n_1785, n_1786, n_1787, 
      n_1788, n_1789, n_1790, n_1791, n_1792, n_1793, n_1794, n_1795, n_1796, 
      n_1797, n_1798, n_1799, n_1800, n_1801, n_1802, n_1803, n_1804, n_1805, 
      n_1806, n_1807, n_1808, n_1809, n_1810, n_1811, n_1812, n_1813, n_1814, 
      n_1815, n_1816, n_1817, n_1818, n_1819, n_1820, n_1821, n_1822, n_1823, 
      n_1824, n_1825, n_1826, n_1827, n_1828, n_1829, n_1830, n_1831, n_1832, 
      n_1833, n_1834, n_1835, n_1836, n_1837, n_1838, n_1839, n_1840, n_1841, 
      n_1842, n_1843, n_1844, n_1845, n_1846, n_1847, n_1848, n_1849, n_1850, 
      n_1851, n_1852, n_1853, n_1854, n_1855, n_1856, n_1857, n_1858, n_1859, 
      n_1860, n_1861, n_1862, n_1863, n_1864, n_1865, n_1866, n_1867, n_1868, 
      n_1869, n_1870, n_1871, n_1872, n_1873, n_1874, n_1875, n_1876, n_1877, 
      n_1878, n_1879, n_1880, n_1881, n_1882, n_1883, n_1884, n_1885, n_1886, 
      n_1887, n_1888, n_1889, n_1890, n_1891, n_1892, n_1893, n_1894, n_1895, 
      n_1896, n_1897, n_1898, n_1899, n_1900, n_1901, n_1902, n_1903, n_1904, 
      n_1905, n_1906, n_1907, n_1908, n_1909, n_1910, n_1911, n_1912, n_1913, 
      n_1914, n_1915, n_1916, n_1917, n_1918, n_1919 : std_logic;

begin
   
   X_Logic0_port <= '0';
   flag_reg1_reg : DFFR_X1 port map( D => mulin_flag, CK => CLK, RN => n60, Q 
                           => flag_reg1, QN => n_1575);
   mux1_reg1_reg_31_inst : DFFR_X1 port map( D => mux1_out_31_port, CK => CLK, 
                           RN => n60, Q => mux1_reg1_31_port, QN => n_1576);
   mux1_reg1_reg_30_inst : DFFR_X1 port map( D => mux1_out_30_port, CK => CLK, 
                           RN => n59, Q => mux1_reg1_30_port, QN => n_1577);
   mux1_reg1_reg_29_inst : DFFR_X1 port map( D => mux1_out_29_port, CK => CLK, 
                           RN => n59, Q => mux1_reg1_29_port, QN => n_1578);
   mux1_reg1_reg_28_inst : DFFR_X1 port map( D => mux1_out_28_port, CK => CLK, 
                           RN => n59, Q => mux1_reg1_28_port, QN => n_1579);
   mux1_reg1_reg_27_inst : DFFR_X1 port map( D => mux1_out_27_port, CK => CLK, 
                           RN => n59, Q => mux1_reg1_27_port, QN => n_1580);
   mux1_reg1_reg_26_inst : DFFR_X1 port map( D => mux1_out_26_port, CK => CLK, 
                           RN => n59, Q => mux1_reg1_26_port, QN => n_1581);
   mux1_reg1_reg_25_inst : DFFR_X1 port map( D => mux1_out_25_port, CK => CLK, 
                           RN => n59, Q => mux1_reg1_25_port, QN => n_1582);
   mux1_reg1_reg_24_inst : DFFR_X1 port map( D => mux1_out_24_port, CK => CLK, 
                           RN => n59, Q => mux1_reg1_24_port, QN => n_1583);
   mux1_reg1_reg_23_inst : DFFR_X1 port map( D => mux1_out_23_port, CK => CLK, 
                           RN => n59, Q => mux1_reg1_23_port, QN => n_1584);
   mux1_reg1_reg_22_inst : DFFR_X1 port map( D => mux1_out_22_port, CK => CLK, 
                           RN => n59, Q => mux1_reg1_22_port, QN => n_1585);
   mux1_reg1_reg_21_inst : DFFR_X1 port map( D => mux1_out_21_port, CK => CLK, 
                           RN => n59, Q => mux1_reg1_21_port, QN => n_1586);
   mux1_reg1_reg_20_inst : DFFR_X1 port map( D => mux1_out_20_port, CK => CLK, 
                           RN => n59, Q => mux1_reg1_20_port, QN => n_1587);
   mux1_reg1_reg_19_inst : DFFR_X1 port map( D => mux1_out_19_port, CK => CLK, 
                           RN => n58, Q => mux1_reg1_19_port, QN => n_1588);
   mux1_reg1_reg_18_inst : DFFR_X1 port map( D => mux1_out_18_port, CK => CLK, 
                           RN => n58, Q => mux1_reg1_18_port, QN => n_1589);
   mux1_reg1_reg_17_inst : DFFR_X1 port map( D => mux1_out_17_port, CK => CLK, 
                           RN => n58, Q => mux1_reg1_17_port, QN => n_1590);
   mux1_reg1_reg_16_inst : DFFR_X1 port map( D => mux1_out_16_port, CK => CLK, 
                           RN => n58, Q => mux1_reg1_16_port, QN => n_1591);
   mux1_reg1_reg_15_inst : DFFR_X1 port map( D => mux1_out_15_port, CK => CLK, 
                           RN => n58, Q => mux1_reg1_15_port, QN => n_1592);
   mux1_reg1_reg_14_inst : DFFR_X1 port map( D => mux1_out_14_port, CK => CLK, 
                           RN => n58, Q => mux1_reg1_14_port, QN => n_1593);
   mux1_reg1_reg_13_inst : DFFR_X1 port map( D => mux1_out_13_port, CK => CLK, 
                           RN => n58, Q => mux1_reg1_13_port, QN => n_1594);
   mux1_reg1_reg_12_inst : DFFR_X1 port map( D => mux1_out_12_port, CK => CLK, 
                           RN => n58, Q => mux1_reg1_12_port, QN => n_1595);
   mux1_reg1_reg_11_inst : DFFR_X1 port map( D => mux1_out_11_port, CK => CLK, 
                           RN => n58, Q => mux1_reg1_11_port, QN => n_1596);
   mux1_reg1_reg_10_inst : DFFR_X1 port map( D => mux1_out_10_port, CK => CLK, 
                           RN => n58, Q => mux1_reg1_10_port, QN => n_1597);
   mux1_reg1_reg_9_inst : DFFR_X1 port map( D => mux1_out_9_port, CK => CLK, RN
                           => n58, Q => mux1_reg1_9_port, QN => n_1598);
   mux1_reg1_reg_8_inst : DFFR_X1 port map( D => mux1_out_8_port, CK => CLK, RN
                           => n57, Q => mux1_reg1_8_port, QN => n_1599);
   mux1_reg1_reg_7_inst : DFFR_X1 port map( D => mux1_out_7_port, CK => CLK, RN
                           => n57, Q => mux1_reg1_7_port, QN => n_1600);
   mux1_reg1_reg_6_inst : DFFR_X1 port map( D => mux1_out_6_port, CK => CLK, RN
                           => n57, Q => mux1_reg1_6_port, QN => n_1601);
   mux1_reg1_reg_5_inst : DFFR_X1 port map( D => mux1_out_5_port, CK => CLK, RN
                           => n57, Q => mux1_reg1_5_port, QN => n_1602);
   mux1_reg1_reg_4_inst : DFFR_X1 port map( D => mux1_out_4_port, CK => CLK, RN
                           => n57, Q => mux1_reg1_4_port, QN => n_1603);
   mux1_reg1_reg_3_inst : DFFR_X1 port map( D => mux1_out_3_port, CK => CLK, RN
                           => n57, Q => mux1_reg1_3_port, QN => n_1604);
   mux1_reg1_reg_2_inst : DFFR_X1 port map( D => mux1_out_2_port, CK => CLK, RN
                           => n57, Q => mux1_reg1_2_port, QN => n_1605);
   mux1_reg1_reg_1_inst : DFFR_X1 port map( D => mux1_out_1_port, CK => CLK, RN
                           => n57, Q => mux1_reg1_1_port, QN => n_1606);
   mux1_reg1_reg_0_inst : DFFR_X1 port map( D => mux1_out_0_port, CK => CLK, RN
                           => n57, Q => mux1_reg1_0_port, QN => n_1607);
   mux2_reg1_reg_31_inst : DFFR_X1 port map( D => mux2_out_31_port, CK => CLK, 
                           RN => n57, Q => mux2_reg1_31_port, QN => n_1608);
   mux2_reg1_reg_30_inst : DFFR_X1 port map( D => mux2_out_30_port, CK => CLK, 
                           RN => n57, Q => mux2_reg1_30_port, QN => n_1609);
   mux2_reg1_reg_29_inst : DFFR_X1 port map( D => mux2_out_29_port, CK => CLK, 
                           RN => n56, Q => mux2_reg1_29_port, QN => n_1610);
   mux2_reg1_reg_28_inst : DFFR_X1 port map( D => mux2_out_28_port, CK => CLK, 
                           RN => n56, Q => mux2_reg1_28_port, QN => n_1611);
   mux2_reg1_reg_27_inst : DFFR_X1 port map( D => mux2_out_27_port, CK => CLK, 
                           RN => n56, Q => mux2_reg1_27_port, QN => n_1612);
   mux2_reg1_reg_26_inst : DFFR_X1 port map( D => mux2_out_26_port, CK => CLK, 
                           RN => n56, Q => mux2_reg1_26_port, QN => n_1613);
   mux2_reg1_reg_25_inst : DFFR_X1 port map( D => mux2_out_25_port, CK => CLK, 
                           RN => n56, Q => mux2_reg1_25_port, QN => n_1614);
   mux2_reg1_reg_24_inst : DFFR_X1 port map( D => mux2_out_24_port, CK => CLK, 
                           RN => n56, Q => mux2_reg1_24_port, QN => n_1615);
   mux2_reg1_reg_23_inst : DFFR_X1 port map( D => mux2_out_23_port, CK => CLK, 
                           RN => n56, Q => mux2_reg1_23_port, QN => n_1616);
   mux2_reg1_reg_22_inst : DFFR_X1 port map( D => mux2_out_22_port, CK => CLK, 
                           RN => n56, Q => mux2_reg1_22_port, QN => n_1617);
   mux2_reg1_reg_21_inst : DFFR_X1 port map( D => mux2_out_21_port, CK => CLK, 
                           RN => n56, Q => mux2_reg1_21_port, QN => n_1618);
   mux2_reg1_reg_20_inst : DFFR_X1 port map( D => mux2_out_20_port, CK => CLK, 
                           RN => n56, Q => mux2_reg1_20_port, QN => n_1619);
   mux2_reg1_reg_19_inst : DFFR_X1 port map( D => mux2_out_19_port, CK => CLK, 
                           RN => n56, Q => mux2_reg1_19_port, QN => n_1620);
   mux2_reg1_reg_18_inst : DFFR_X1 port map( D => mux2_out_18_port, CK => CLK, 
                           RN => n55, Q => mux2_reg1_18_port, QN => n_1621);
   mux2_reg1_reg_17_inst : DFFR_X1 port map( D => mux2_out_17_port, CK => CLK, 
                           RN => n55, Q => mux2_reg1_17_port, QN => n_1622);
   mux2_reg1_reg_16_inst : DFFR_X1 port map( D => mux2_out_16_port, CK => CLK, 
                           RN => n55, Q => mux2_reg1_16_port, QN => n_1623);
   mux2_reg1_reg_15_inst : DFFR_X1 port map( D => mux2_out_15_port, CK => CLK, 
                           RN => n55, Q => mux2_reg1_15_port, QN => n_1624);
   mux2_reg1_reg_14_inst : DFFR_X1 port map( D => mux2_out_14_port, CK => CLK, 
                           RN => n55, Q => mux2_reg1_14_port, QN => n_1625);
   mux2_reg1_reg_13_inst : DFFR_X1 port map( D => mux2_out_13_port, CK => CLK, 
                           RN => n55, Q => mux2_reg1_13_port, QN => n_1626);
   mux2_reg1_reg_12_inst : DFFR_X1 port map( D => mux2_out_12_port, CK => CLK, 
                           RN => n55, Q => mux2_reg1_12_port, QN => n_1627);
   mux2_reg1_reg_11_inst : DFFR_X1 port map( D => mux2_out_11_port, CK => CLK, 
                           RN => n55, Q => mux2_reg1_11_port, QN => n_1628);
   mux2_reg1_reg_10_inst : DFFR_X1 port map( D => mux2_out_10_port, CK => CLK, 
                           RN => n55, Q => mux2_reg1_10_port, QN => n_1629);
   mux2_reg1_reg_9_inst : DFFR_X1 port map( D => mux2_out_9_port, CK => CLK, RN
                           => n55, Q => mux2_reg1_9_port, QN => n_1630);
   mux2_reg1_reg_8_inst : DFFR_X1 port map( D => mux2_out_8_port, CK => CLK, RN
                           => n55, Q => mux2_reg1_8_port, QN => n_1631);
   mux2_reg1_reg_7_inst : DFFR_X1 port map( D => mux2_out_7_port, CK => CLK, RN
                           => n54, Q => mux2_reg1_7_port, QN => n_1632);
   mux2_reg1_reg_6_inst : DFFR_X1 port map( D => mux2_out_6_port, CK => CLK, RN
                           => n54, Q => mux2_reg1_6_port, QN => n_1633);
   mux2_reg1_reg_5_inst : DFFR_X1 port map( D => mux2_out_5_port, CK => CLK, RN
                           => n54, Q => mux2_reg1_5_port, QN => n_1634);
   mux2_reg1_reg_4_inst : DFFR_X1 port map( D => mux2_out_4_port, CK => CLK, RN
                           => n54, Q => mux2_reg1_4_port, QN => n_1635);
   mux2_reg1_reg_3_inst : DFFR_X1 port map( D => mux2_out_3_port, CK => CLK, RN
                           => n54, Q => mux2_reg1_3_port, QN => n_1636);
   mux2_reg1_reg_2_inst : DFFR_X1 port map( D => mux2_out_2_port, CK => CLK, RN
                           => n54, Q => mux2_reg1_2_port, QN => n_1637);
   mux2_reg1_reg_1_inst : DFFR_X1 port map( D => mux2_out_1_port, CK => CLK, RN
                           => n54, Q => mux2_reg1_1_port, QN => n_1638);
   mux2_reg1_reg_0_inst : DFFR_X1 port map( D => mux2_out_0_port, CK => CLK, RN
                           => n54, Q => mux2_reg1_0_port, QN => n_1639);
   A4_reg1_reg_31_inst : DFFR_X1 port map( D => s_8A_1_31_port, CK => CLK, RN 
                           => n54, Q => A4_reg1_31_port, QN => n_1640);
   A4_reg1_reg_30_inst : DFFR_X1 port map( D => s_8A_1_30_port, CK => CLK, RN 
                           => n54, Q => A4_reg1_30_port, QN => n_1641);
   A4_reg1_reg_29_inst : DFFR_X1 port map( D => s_8A_1_29_port, CK => CLK, RN 
                           => n54, Q => A4_reg1_29_port, QN => n_1642);
   A4_reg1_reg_28_inst : DFFR_X1 port map( D => s_8A_1_28_port, CK => CLK, RN 
                           => n53, Q => A4_reg1_28_port, QN => n_1643);
   A4_reg1_reg_27_inst : DFFR_X1 port map( D => s_8A_1_27_port, CK => CLK, RN 
                           => n53, Q => A4_reg1_27_port, QN => n_1644);
   A4_reg1_reg_26_inst : DFFR_X1 port map( D => s_8A_1_26_port, CK => CLK, RN 
                           => n53, Q => A4_reg1_26_port, QN => n_1645);
   A4_reg1_reg_25_inst : DFFR_X1 port map( D => s_8A_1_25_port, CK => CLK, RN 
                           => n53, Q => A4_reg1_25_port, QN => n_1646);
   A4_reg1_reg_24_inst : DFFR_X1 port map( D => s_8A_1_24_port, CK => CLK, RN 
                           => n53, Q => A4_reg1_24_port, QN => n_1647);
   A4_reg1_reg_23_inst : DFFR_X1 port map( D => s_8A_1_23_port, CK => CLK, RN 
                           => n53, Q => A4_reg1_23_port, QN => n_1648);
   A4_reg1_reg_22_inst : DFFR_X1 port map( D => s_8A_1_22_port, CK => CLK, RN 
                           => n53, Q => A4_reg1_22_port, QN => n_1649);
   A4_reg1_reg_21_inst : DFFR_X1 port map( D => s_8A_1_21_port, CK => CLK, RN 
                           => n53, Q => A4_reg1_21_port, QN => n_1650);
   A4_reg1_reg_20_inst : DFFR_X1 port map( D => s_8A_1_20_port, CK => CLK, RN 
                           => n53, Q => A4_reg1_20_port, QN => n_1651);
   A4_reg1_reg_19_inst : DFFR_X1 port map( D => s_8A_1_19_port, CK => CLK, RN 
                           => n53, Q => A4_reg1_19_port, QN => n_1652);
   A4_reg1_reg_18_inst : DFFR_X1 port map( D => s_8A_1_18_port, CK => CLK, RN 
                           => n53, Q => A4_reg1_18_port, QN => n_1653);
   A4_reg1_reg_17_inst : DFFR_X1 port map( D => s_8A_1_17_port, CK => CLK, RN 
                           => n52, Q => A4_reg1_17_port, QN => n_1654);
   A4_reg1_reg_16_inst : DFFR_X1 port map( D => s_8A_1_16_port, CK => CLK, RN 
                           => n52, Q => A4_reg1_16_port, QN => n_1655);
   A4_reg1_reg_15_inst : DFFR_X1 port map( D => s_8A_1_15_port, CK => CLK, RN 
                           => n52, Q => A4_reg1_15_port, QN => n_1656);
   A4_reg1_reg_14_inst : DFFR_X1 port map( D => s_8A_1_14_port, CK => CLK, RN 
                           => n52, Q => A4_reg1_14_port, QN => n_1657);
   A4_reg1_reg_13_inst : DFFR_X1 port map( D => s_8A_1_13_port, CK => CLK, RN 
                           => n52, Q => A4_reg1_13_port, QN => n_1658);
   A4_reg1_reg_12_inst : DFFR_X1 port map( D => s_8A_1_12_port, CK => CLK, RN 
                           => n52, Q => A4_reg1_12_port, QN => n_1659);
   A4_reg1_reg_11_inst : DFFR_X1 port map( D => s_8A_1_11_port, CK => CLK, RN 
                           => n52, Q => A4_reg1_11_port, QN => n_1660);
   A4_reg1_reg_10_inst : DFFR_X1 port map( D => s_8A_1_10_port, CK => CLK, RN 
                           => n52, Q => A4_reg1_10_port, QN => n_1661);
   A4_reg1_reg_9_inst : DFFR_X1 port map( D => s_8A_1_9_port, CK => CLK, RN => 
                           n52, Q => A4_reg1_9_port, QN => n_1662);
   A4_reg1_reg_8_inst : DFFR_X1 port map( D => s_8A_1_8_port, CK => CLK, RN => 
                           n52, Q => A4_reg1_8_port, QN => n_1663);
   A4_reg1_reg_7_inst : DFFR_X1 port map( D => s_8A_1_7_port, CK => CLK, RN => 
                           n52, Q => A4_reg1_7_port, QN => n_1664);
   A4_reg1_reg_6_inst : DFFR_X1 port map( D => s_8A_1_6_port, CK => CLK, RN => 
                           n51, Q => A4_reg1_6_port, QN => n_1665);
   A4_reg1_reg_5_inst : DFFR_X1 port map( D => s_8A_1_5_port, CK => CLK, RN => 
                           n51, Q => A4_reg1_5_port, QN => n_1666);
   A4_reg1_reg_4_inst : DFFR_X1 port map( D => s_8A_1_4_port, CK => CLK, RN => 
                           n51, Q => A4_reg1_4_port, QN => n_1667);
   A4_reg1_reg_3_inst : DFFR_X1 port map( D => s_8A_1_3_port, CK => CLK, RN => 
                           n51, Q => A4_reg1_3_port, QN => n_1668);
   flag_reg2_reg : DFFR_X1 port map( D => flag_reg1, CK => CLK, RN => n51, Q =>
                           flag_reg2, QN => n_1669);
   sum_reg2_reg_63_inst : DFFR_X1 port map( D => sum_2_out_63_port, CK => CLK, 
                           RN => n51, Q => sum_reg2_63_port, QN => n_1670);
   sum_reg2_reg_62_inst : DFFR_X1 port map( D => sum_2_out_62_port, CK => CLK, 
                           RN => n51, Q => sum_reg2_62_port, QN => n_1671);
   sum_reg2_reg_61_inst : DFFR_X1 port map( D => sum_2_out_61_port, CK => CLK, 
                           RN => n51, Q => sum_reg2_61_port, QN => n_1672);
   sum_reg2_reg_60_inst : DFFR_X1 port map( D => sum_2_out_60_port, CK => CLK, 
                           RN => n50, Q => sum_reg2_60_port, QN => n_1673);
   sum_reg2_reg_59_inst : DFFR_X1 port map( D => sum_2_out_59_port, CK => CLK, 
                           RN => n50, Q => sum_reg2_59_port, QN => n_1674);
   sum_reg2_reg_58_inst : DFFR_X1 port map( D => sum_2_out_58_port, CK => CLK, 
                           RN => n50, Q => sum_reg2_58_port, QN => n_1675);
   sum_reg2_reg_57_inst : DFFR_X1 port map( D => sum_2_out_57_port, CK => CLK, 
                           RN => n50, Q => sum_reg2_57_port, QN => n_1676);
   sum_reg2_reg_56_inst : DFFR_X1 port map( D => sum_2_out_56_port, CK => CLK, 
                           RN => n50, Q => sum_reg2_56_port, QN => n_1677);
   sum_reg2_reg_55_inst : DFFR_X1 port map( D => sum_2_out_55_port, CK => CLK, 
                           RN => n50, Q => sum_reg2_55_port, QN => n_1678);
   sum_reg2_reg_54_inst : DFFR_X1 port map( D => sum_2_out_54_port, CK => CLK, 
                           RN => n50, Q => sum_reg2_54_port, QN => n_1679);
   sum_reg2_reg_53_inst : DFFR_X1 port map( D => sum_2_out_53_port, CK => CLK, 
                           RN => n50, Q => sum_reg2_53_port, QN => n_1680);
   sum_reg2_reg_52_inst : DFFR_X1 port map( D => sum_2_out_52_port, CK => CLK, 
                           RN => n50, Q => sum_reg2_52_port, QN => n_1681);
   sum_reg2_reg_51_inst : DFFR_X1 port map( D => sum_2_out_51_port, CK => CLK, 
                           RN => n50, Q => sum_reg2_51_port, QN => n_1682);
   sum_reg2_reg_50_inst : DFFR_X1 port map( D => sum_2_out_50_port, CK => CLK, 
                           RN => n50, Q => sum_reg2_50_port, QN => n_1683);
   sum_reg2_reg_49_inst : DFFR_X1 port map( D => sum_2_out_49_port, CK => CLK, 
                           RN => n49, Q => sum_reg2_49_port, QN => n_1684);
   sum_reg2_reg_48_inst : DFFR_X1 port map( D => sum_2_out_48_port, CK => CLK, 
                           RN => n49, Q => sum_reg2_48_port, QN => n_1685);
   sum_reg2_reg_47_inst : DFFR_X1 port map( D => sum_2_out_47_port, CK => CLK, 
                           RN => n49, Q => sum_reg2_47_port, QN => n_1686);
   sum_reg2_reg_46_inst : DFFR_X1 port map( D => sum_2_out_46_port, CK => CLK, 
                           RN => n49, Q => sum_reg2_46_port, QN => n_1687);
   sum_reg2_reg_45_inst : DFFR_X1 port map( D => sum_2_out_45_port, CK => CLK, 
                           RN => n49, Q => sum_reg2_45_port, QN => n_1688);
   sum_reg2_reg_44_inst : DFFR_X1 port map( D => sum_2_out_44_port, CK => CLK, 
                           RN => n49, Q => sum_reg2_44_port, QN => n_1689);
   sum_reg2_reg_43_inst : DFFR_X1 port map( D => sum_2_out_43_port, CK => CLK, 
                           RN => n49, Q => sum_reg2_43_port, QN => n_1690);
   sum_reg2_reg_42_inst : DFFR_X1 port map( D => sum_2_out_42_port, CK => CLK, 
                           RN => n49, Q => sum_reg2_42_port, QN => n_1691);
   sum_reg2_reg_41_inst : DFFR_X1 port map( D => sum_2_out_41_port, CK => CLK, 
                           RN => n49, Q => sum_reg2_41_port, QN => n_1692);
   sum_reg2_reg_40_inst : DFFR_X1 port map( D => sum_2_out_40_port, CK => CLK, 
                           RN => n49, Q => sum_reg2_40_port, QN => n_1693);
   sum_reg2_reg_39_inst : DFFR_X1 port map( D => sum_2_out_39_port, CK => CLK, 
                           RN => n49, Q => sum_reg2_39_port, QN => n_1694);
   sum_reg2_reg_38_inst : DFFR_X1 port map( D => sum_2_out_38_port, CK => CLK, 
                           RN => n48, Q => sum_reg2_38_port, QN => n_1695);
   sum_reg2_reg_37_inst : DFFR_X1 port map( D => sum_2_out_37_port, CK => CLK, 
                           RN => n48, Q => sum_reg2_37_port, QN => n_1696);
   sum_reg2_reg_36_inst : DFFR_X1 port map( D => sum_2_out_36_port, CK => CLK, 
                           RN => n48, Q => sum_reg2_36_port, QN => n_1697);
   sum_reg2_reg_35_inst : DFFR_X1 port map( D => sum_2_out_35_port, CK => CLK, 
                           RN => n48, Q => sum_reg2_35_port, QN => n_1698);
   sum_reg2_reg_34_inst : DFFR_X1 port map( D => sum_2_out_34_port, CK => CLK, 
                           RN => n48, Q => sum_reg2_34_port, QN => n_1699);
   sum_reg2_reg_33_inst : DFFR_X1 port map( D => sum_2_out_33_port, CK => CLK, 
                           RN => n48, Q => sum_reg2_33_port, QN => n_1700);
   sum_reg2_reg_32_inst : DFFR_X1 port map( D => sum_2_out_32_port, CK => CLK, 
                           RN => n48, Q => sum_reg2_32_port, QN => n_1701);
   sum_reg2_reg_31_inst : DFFR_X1 port map( D => sum_2_out_31_port, CK => CLK, 
                           RN => n48, Q => sum_reg2_31_port, QN => n_1702);
   sum_reg2_reg_30_inst : DFFR_X1 port map( D => sum_2_out_30_port, CK => CLK, 
                           RN => n48, Q => sum_reg2_30_port, QN => n_1703);
   sum_reg2_reg_29_inst : DFFR_X1 port map( D => sum_2_out_29_port, CK => CLK, 
                           RN => n48, Q => sum_reg2_29_port, QN => n_1704);
   sum_reg2_reg_28_inst : DFFR_X1 port map( D => sum_2_out_28_port, CK => CLK, 
                           RN => n48, Q => sum_reg2_28_port, QN => n_1705);
   sum_reg2_reg_27_inst : DFFR_X1 port map( D => sum_2_out_27_port, CK => CLK, 
                           RN => n47, Q => sum_reg2_27_port, QN => n_1706);
   sum_reg2_reg_26_inst : DFFR_X1 port map( D => sum_2_out_26_port, CK => CLK, 
                           RN => n47, Q => sum_reg2_26_port, QN => n_1707);
   sum_reg2_reg_25_inst : DFFR_X1 port map( D => sum_2_out_25_port, CK => CLK, 
                           RN => n47, Q => sum_reg2_25_port, QN => n_1708);
   sum_reg2_reg_24_inst : DFFR_X1 port map( D => sum_2_out_24_port, CK => CLK, 
                           RN => n47, Q => sum_reg2_24_port, QN => n_1709);
   sum_reg2_reg_23_inst : DFFR_X1 port map( D => sum_2_out_23_port, CK => CLK, 
                           RN => n47, Q => sum_reg2_23_port, QN => n_1710);
   sum_reg2_reg_22_inst : DFFR_X1 port map( D => sum_2_out_22_port, CK => CLK, 
                           RN => n47, Q => sum_reg2_22_port, QN => n_1711);
   sum_reg2_reg_21_inst : DFFR_X1 port map( D => sum_2_out_21_port, CK => CLK, 
                           RN => n47, Q => sum_reg2_21_port, QN => n_1712);
   sum_reg2_reg_20_inst : DFFR_X1 port map( D => sum_2_out_20_port, CK => CLK, 
                           RN => n47, Q => sum_reg2_20_port, QN => n_1713);
   sum_reg2_reg_19_inst : DFFR_X1 port map( D => sum_2_out_19_port, CK => CLK, 
                           RN => n47, Q => sum_reg2_19_port, QN => n_1714);
   sum_reg2_reg_18_inst : DFFR_X1 port map( D => sum_2_out_18_port, CK => CLK, 
                           RN => n47, Q => sum_reg2_18_port, QN => n_1715);
   sum_reg2_reg_17_inst : DFFR_X1 port map( D => sum_2_out_17_port, CK => CLK, 
                           RN => n47, Q => sum_reg2_17_port, QN => n_1716);
   sum_reg2_reg_16_inst : DFFR_X1 port map( D => sum_2_out_16_port, CK => CLK, 
                           RN => n46, Q => sum_reg2_16_port, QN => n_1717);
   sum_reg2_reg_15_inst : DFFR_X1 port map( D => sum_2_out_15_port, CK => CLK, 
                           RN => n46, Q => sum_reg2_15_port, QN => n_1718);
   sum_reg2_reg_14_inst : DFFR_X1 port map( D => sum_2_out_14_port, CK => CLK, 
                           RN => n46, Q => sum_reg2_14_port, QN => n_1719);
   sum_reg2_reg_13_inst : DFFR_X1 port map( D => sum_2_out_13_port, CK => CLK, 
                           RN => n46, Q => sum_reg2_13_port, QN => n_1720);
   sum_reg2_reg_12_inst : DFFR_X1 port map( D => sum_2_out_12_port, CK => CLK, 
                           RN => n46, Q => sum_reg2_12_port, QN => n_1721);
   sum_reg2_reg_11_inst : DFFR_X1 port map( D => sum_2_out_11_port, CK => CLK, 
                           RN => n46, Q => sum_reg2_11_port, QN => n_1722);
   sum_reg2_reg_10_inst : DFFR_X1 port map( D => sum_2_out_10_port, CK => CLK, 
                           RN => n46, Q => sum_reg2_10_port, QN => n_1723);
   sum_reg2_reg_9_inst : DFFR_X1 port map( D => sum_2_out_9_port, CK => CLK, RN
                           => n46, Q => sum_reg2_9_port, QN => n_1724);
   sum_reg2_reg_8_inst : DFFR_X1 port map( D => sum_2_out_8_port, CK => CLK, RN
                           => n46, Q => sum_reg2_8_port, QN => n_1725);
   sum_reg2_reg_7_inst : DFFR_X1 port map( D => sum_2_out_7_port, CK => CLK, RN
                           => n46, Q => sum_reg2_7_port, QN => n_1726);
   sum_reg2_reg_6_inst : DFFR_X1 port map( D => sum_2_out_6_port, CK => CLK, RN
                           => n46, Q => sum_reg2_6_port, QN => n_1727);
   sum_reg2_reg_5_inst : DFFR_X1 port map( D => sum_2_out_5_port, CK => CLK, RN
                           => n45, Q => sum_reg2_5_port, QN => n_1728);
   sum_reg2_reg_4_inst : DFFR_X1 port map( D => sum_2_out_4_port, CK => CLK, RN
                           => n45, Q => sum_reg2_4_port, QN => n_1729);
   sum_reg2_reg_3_inst : DFFR_X1 port map( D => sum_2_out_3_port, CK => CLK, RN
                           => n45, Q => sum_reg2_3_port, QN => n_1730);
   sum_reg2_reg_2_inst : DFFR_X1 port map( D => sum_2_out_2_port, CK => CLK, RN
                           => n45, Q => sum_reg2_2_port, QN => n_1731);
   sum_reg2_reg_1_inst : DFFR_X1 port map( D => sum_2_out_1_port, CK => CLK, RN
                           => n45, Q => sum_reg2_1_port, QN => n_1732);
   sum_reg2_reg_0_inst : DFFR_X1 port map( D => sum_2_out_0_port, CK => CLK, RN
                           => n45, Q => sum_reg2_0_port, QN => n_1733);
   A4_reg2_reg_31_inst : DFFR_X1 port map( D => s_2A_2_31_port, CK => CLK, RN 
                           => n45, Q => A4_reg2_31_port, QN => n_1734);
   A4_reg2_reg_30_inst : DFFR_X1 port map( D => s_2A_2_30_port, CK => CLK, RN 
                           => n45, Q => A4_reg2_30_port, QN => n_1735);
   A4_reg2_reg_29_inst : DFFR_X1 port map( D => s_2A_2_29_port, CK => CLK, RN 
                           => n45, Q => A4_reg2_29_port, QN => n_1736);
   A4_reg2_reg_28_inst : DFFR_X1 port map( D => s_2A_2_28_port, CK => CLK, RN 
                           => n45, Q => A4_reg2_28_port, QN => n_1737);
   A4_reg2_reg_27_inst : DFFR_X1 port map( D => s_2A_2_27_port, CK => CLK, RN 
                           => n45, Q => A4_reg2_27_port, QN => n_1738);
   A4_reg2_reg_26_inst : DFFR_X1 port map( D => s_2A_2_26_port, CK => CLK, RN 
                           => n44, Q => A4_reg2_26_port, QN => n_1739);
   A4_reg2_reg_25_inst : DFFR_X1 port map( D => s_2A_2_25_port, CK => CLK, RN 
                           => n44, Q => A4_reg2_25_port, QN => n_1740);
   A4_reg2_reg_24_inst : DFFR_X1 port map( D => s_2A_2_24_port, CK => CLK, RN 
                           => n44, Q => A4_reg2_24_port, QN => n_1741);
   A4_reg2_reg_23_inst : DFFR_X1 port map( D => s_2A_2_23_port, CK => CLK, RN 
                           => n44, Q => A4_reg2_23_port, QN => n_1742);
   A4_reg2_reg_22_inst : DFFR_X1 port map( D => s_2A_2_22_port, CK => CLK, RN 
                           => n44, Q => A4_reg2_22_port, QN => n_1743);
   A4_reg2_reg_21_inst : DFFR_X1 port map( D => s_2A_2_21_port, CK => CLK, RN 
                           => n44, Q => A4_reg2_21_port, QN => n_1744);
   A4_reg2_reg_20_inst : DFFR_X1 port map( D => s_2A_2_20_port, CK => CLK, RN 
                           => n44, Q => A4_reg2_20_port, QN => n_1745);
   A4_reg2_reg_19_inst : DFFR_X1 port map( D => s_2A_2_19_port, CK => CLK, RN 
                           => n44, Q => A4_reg2_19_port, QN => n_1746);
   A4_reg2_reg_18_inst : DFFR_X1 port map( D => s_2A_2_18_port, CK => CLK, RN 
                           => n44, Q => A4_reg2_18_port, QN => n_1747);
   A4_reg2_reg_17_inst : DFFR_X1 port map( D => s_2A_2_17_port, CK => CLK, RN 
                           => n44, Q => A4_reg2_17_port, QN => n_1748);
   A4_reg2_reg_16_inst : DFFR_X1 port map( D => s_2A_2_16_port, CK => CLK, RN 
                           => n44, Q => A4_reg2_16_port, QN => n_1749);
   A4_reg2_reg_15_inst : DFFR_X1 port map( D => s_2A_2_15_port, CK => CLK, RN 
                           => n43, Q => A4_reg2_15_port, QN => n_1750);
   A4_reg2_reg_14_inst : DFFR_X1 port map( D => s_2A_2_14_port, CK => CLK, RN 
                           => n43, Q => A4_reg2_14_port, QN => n_1751);
   A4_reg2_reg_13_inst : DFFR_X1 port map( D => s_2A_2_13_port, CK => CLK, RN 
                           => n43, Q => A4_reg2_13_port, QN => n_1752);
   A4_reg2_reg_12_inst : DFFR_X1 port map( D => s_2A_2_12_port, CK => CLK, RN 
                           => n43, Q => A4_reg2_12_port, QN => n_1753);
   A4_reg2_reg_11_inst : DFFR_X1 port map( D => s_2A_2_11_port, CK => CLK, RN 
                           => n43, Q => A4_reg2_11_port, QN => n_1754);
   A4_reg2_reg_10_inst : DFFR_X1 port map( D => s_2A_2_10_port, CK => CLK, RN 
                           => n43, Q => A4_reg2_10_port, QN => n_1755);
   A4_reg2_reg_9_inst : DFFR_X1 port map( D => s_2A_2_9_port, CK => CLK, RN => 
                           n43, Q => A4_reg2_9_port, QN => n_1756);
   A4_reg2_reg_8_inst : DFFR_X1 port map( D => s_2A_2_8_port, CK => CLK, RN => 
                           n43, Q => A4_reg2_8_port, QN => n_1757);
   A4_reg2_reg_7_inst : DFFR_X1 port map( D => s_2A_2_7_port, CK => CLK, RN => 
                           n43, Q => A4_reg2_7_port, QN => n_1758);
   A4_reg2_reg_6_inst : DFFR_X1 port map( D => s_2A_2_6_port, CK => CLK, RN => 
                           n43, Q => A4_reg2_6_port, QN => n_1759);
   A4_reg2_reg_5_inst : DFFR_X1 port map( D => s_2A_2_5_port, CK => CLK, RN => 
                           n43, Q => A4_reg2_5_port, QN => n_1760);
   A4_reg2_reg_4_inst : DFFR_X1 port map( D => s_2A_2_4_port, CK => CLK, RN => 
                           n42, Q => A4_reg2_4_port, QN => n_1761);
   A4_reg2_reg_3_inst : DFFR_X1 port map( D => s_2A_2_3_port, CK => CLK, RN => 
                           n42, Q => A4_reg2_3_port, QN => n_1762);
   A4_reg2_reg_2_inst : DFFR_X1 port map( D => s_2A_2_2_port, CK => CLK, RN => 
                           n42, Q => A4_reg2_2_port, QN => n_1763);
   flag_reg3_reg : DFFR_X1 port map( D => flag_reg2, CK => CLK, RN => n42, Q =>
                           MULready, QN => n_1764);
   enc_reg21_reg_2_inst : DFFR_X1 port map( D => s_sel_2_2_port, CK => CLK, RN 
                           => n42, Q => enc_reg21_2_port, QN => n_1765);
   enc_reg21_reg_1_inst : DFFR_X1 port map( D => s_sel_2_1_port, CK => CLK, RN 
                           => n42, Q => enc_reg21_1_port, QN => n_1766);
   enc_reg21_reg_0_inst : DFFR_X1 port map( D => s_sel_2_0_port, CK => CLK, RN 
                           => n42, Q => enc_reg21_0_port, QN => n_1767);
   mux_reg2_reg_0_inst : DFFR_X1 port map( D => mux_2_out_0_port, CK => CLK, RN
                           => n42, Q => mux_reg2_0_port, QN => n_1768);
   mux_reg2_reg_1_inst : DFFR_X1 port map( D => mux_2_out_1_port, CK => CLK, RN
                           => n42, Q => mux_reg2_1_port, QN => n_1769);
   mux_reg2_reg_2_inst : DFFR_X1 port map( D => mux_2_out_2_port, CK => CLK, RN
                           => n41, Q => mux_reg2_2_port, QN => n_1770);
   mux_reg2_reg_3_inst : DFFR_X1 port map( D => mux_2_out_3_port, CK => CLK, RN
                           => n41, Q => mux_reg2_3_port, QN => n_1771);
   mux_reg2_reg_4_inst : DFFR_X1 port map( D => mux_2_out_4_port, CK => CLK, RN
                           => n41, Q => mux_reg2_4_port, QN => n_1772);
   mux_reg2_reg_5_inst : DFFR_X1 port map( D => mux_2_out_5_port, CK => CLK, RN
                           => n41, Q => mux_reg2_5_port, QN => n_1773);
   mux_reg2_reg_6_inst : DFFR_X1 port map( D => mux_2_out_6_port, CK => CLK, RN
                           => n41, Q => mux_reg2_6_port, QN => n_1774);
   mux_reg2_reg_7_inst : DFFR_X1 port map( D => mux_2_out_7_port, CK => CLK, RN
                           => n41, Q => mux_reg2_7_port, QN => n_1775);
   mux_reg2_reg_8_inst : DFFR_X1 port map( D => mux_2_out_8_port, CK => CLK, RN
                           => n41, Q => mux_reg2_8_port, QN => n_1776);
   mux_reg2_reg_9_inst : DFFR_X1 port map( D => mux_2_out_9_port, CK => CLK, RN
                           => n41, Q => mux_reg2_9_port, QN => n_1777);
   mux_reg2_reg_10_inst : DFFR_X1 port map( D => mux_2_out_10_port, CK => CLK, 
                           RN => n41, Q => mux_reg2_10_port, QN => n_1778);
   mux_reg2_reg_11_inst : DFFR_X1 port map( D => mux_2_out_11_port, CK => CLK, 
                           RN => n41, Q => mux_reg2_11_port, QN => n_1779);
   mux_reg2_reg_12_inst : DFFR_X1 port map( D => mux_2_out_12_port, CK => CLK, 
                           RN => n41, Q => mux_reg2_12_port, QN => n_1780);
   mux_reg2_reg_13_inst : DFFR_X1 port map( D => mux_2_out_13_port, CK => CLK, 
                           RN => n40, Q => mux_reg2_13_port, QN => n_1781);
   mux_reg2_reg_14_inst : DFFR_X1 port map( D => mux_2_out_14_port, CK => CLK, 
                           RN => n40, Q => mux_reg2_14_port, QN => n_1782);
   mux_reg2_reg_15_inst : DFFR_X1 port map( D => mux_2_out_15_port, CK => CLK, 
                           RN => n40, Q => mux_reg2_15_port, QN => n_1783);
   mux_reg2_reg_16_inst : DFFR_X1 port map( D => mux_2_out_16_port, CK => CLK, 
                           RN => n40, Q => mux_reg2_16_port, QN => n_1784);
   mux_reg2_reg_17_inst : DFFR_X1 port map( D => mux_2_out_17_port, CK => CLK, 
                           RN => n40, Q => mux_reg2_17_port, QN => n_1785);
   mux_reg2_reg_18_inst : DFFR_X1 port map( D => mux_2_out_18_port, CK => CLK, 
                           RN => n40, Q => mux_reg2_18_port, QN => n_1786);
   mux_reg2_reg_19_inst : DFFR_X1 port map( D => mux_2_out_19_port, CK => CLK, 
                           RN => n40, Q => mux_reg2_19_port, QN => n_1787);
   mux_reg2_reg_20_inst : DFFR_X1 port map( D => mux_2_out_20_port, CK => CLK, 
                           RN => n40, Q => mux_reg2_20_port, QN => n_1788);
   mux_reg2_reg_21_inst : DFFR_X1 port map( D => mux_2_out_21_port, CK => CLK, 
                           RN => n40, Q => mux_reg2_21_port, QN => n_1789);
   mux_reg2_reg_22_inst : DFFR_X1 port map( D => mux_2_out_22_port, CK => CLK, 
                           RN => n40, Q => mux_reg2_22_port, QN => n_1790);
   mux_reg2_reg_23_inst : DFFR_X1 port map( D => mux_2_out_23_port, CK => CLK, 
                           RN => n40, Q => mux_reg2_23_port, QN => n_1791);
   mux_reg2_reg_24_inst : DFFR_X1 port map( D => mux_2_out_24_port, CK => CLK, 
                           RN => n39, Q => mux_reg2_24_port, QN => n_1792);
   mux_reg2_reg_25_inst : DFFR_X1 port map( D => mux_2_out_25_port, CK => CLK, 
                           RN => n39, Q => mux_reg2_25_port, QN => n_1793);
   mux_reg2_reg_26_inst : DFFR_X1 port map( D => mux_2_out_26_port, CK => CLK, 
                           RN => n39, Q => mux_reg2_26_port, QN => n_1794);
   mux_reg2_reg_27_inst : DFFR_X1 port map( D => mux_2_out_27_port, CK => CLK, 
                           RN => n39, Q => mux_reg2_27_port, QN => n_1795);
   mux_reg2_reg_28_inst : DFFR_X1 port map( D => mux_2_out_28_port, CK => CLK, 
                           RN => n39, Q => mux_reg2_28_port, QN => n_1796);
   mux_reg2_reg_29_inst : DFFR_X1 port map( D => mux_2_out_29_port, CK => CLK, 
                           RN => n39, Q => mux_reg2_29_port, QN => n_1797);
   mux_reg2_reg_30_inst : DFFR_X1 port map( D => mux_2_out_30_port, CK => CLK, 
                           RN => n39, Q => mux_reg2_30_port, QN => n_1798);
   mux_reg2_reg_31_inst : DFFR_X1 port map( D => mux_2_out_31_port, CK => CLK, 
                           RN => n39, Q => mux_reg2_31_port, QN => n_1799);
   sum_reg3_reg_0_inst : DFFR_X1 port map( D => sum_3_out_0_port, CK => CLK, RN
                           => n39, Q => sum_reg3_0_port, QN => n_1800);
   sum_reg3_reg_1_inst : DFFR_X1 port map( D => sum_3_out_1_port, CK => CLK, RN
                           => n39, Q => sum_reg3_1_port, QN => n_1801);
   sum_reg3_reg_2_inst : DFFR_X1 port map( D => sum_3_out_2_port, CK => CLK, RN
                           => n39, Q => sum_reg3_2_port, QN => n_1802);
   sum_reg3_reg_3_inst : DFFR_X1 port map( D => sum_3_out_3_port, CK => CLK, RN
                           => n38, Q => sum_reg3_3_port, QN => n_1803);
   sum_reg3_reg_4_inst : DFFR_X1 port map( D => sum_3_out_4_port, CK => CLK, RN
                           => n38, Q => sum_reg3_4_port, QN => n_1804);
   sum_reg3_reg_5_inst : DFFR_X1 port map( D => sum_3_out_5_port, CK => CLK, RN
                           => n38, Q => sum_reg3_5_port, QN => n_1805);
   sum_reg3_reg_6_inst : DFFR_X1 port map( D => sum_3_out_6_port, CK => CLK, RN
                           => n38, Q => sum_reg3_6_port, QN => n_1806);
   sum_reg3_reg_7_inst : DFFR_X1 port map( D => sum_3_out_7_port, CK => CLK, RN
                           => n38, Q => sum_reg3_7_port, QN => n_1807);
   sum_reg3_reg_8_inst : DFFR_X1 port map( D => sum_3_out_8_port, CK => CLK, RN
                           => n38, Q => sum_reg3_8_port, QN => n_1808);
   sum_reg3_reg_9_inst : DFFR_X1 port map( D => sum_3_out_9_port, CK => CLK, RN
                           => n38, Q => sum_reg3_9_port, QN => n_1809);
   sum_reg3_reg_10_inst : DFFR_X1 port map( D => sum_3_out_10_port, CK => CLK, 
                           RN => n38, Q => sum_reg3_10_port, QN => n_1810);
   sum_reg3_reg_11_inst : DFFR_X1 port map( D => sum_3_out_11_port, CK => CLK, 
                           RN => n38, Q => sum_reg3_11_port, QN => n_1811);
   sum_reg3_reg_12_inst : DFFR_X1 port map( D => sum_3_out_12_port, CK => CLK, 
                           RN => n38, Q => sum_reg3_12_port, QN => n_1812);
   sum_reg3_reg_13_inst : DFFR_X1 port map( D => sum_3_out_13_port, CK => CLK, 
                           RN => n38, Q => sum_reg3_13_port, QN => n_1813);
   sum_reg3_reg_14_inst : DFFR_X1 port map( D => sum_3_out_14_port, CK => CLK, 
                           RN => n37, Q => sum_reg3_14_port, QN => n_1814);
   sum_reg3_reg_15_inst : DFFR_X1 port map( D => sum_3_out_15_port, CK => CLK, 
                           RN => n37, Q => sum_reg3_15_port, QN => n_1815);
   sum_reg3_reg_16_inst : DFFR_X1 port map( D => sum_3_out_16_port, CK => CLK, 
                           RN => n37, Q => sum_reg3_16_port, QN => n_1816);
   sum_reg3_reg_17_inst : DFFR_X1 port map( D => sum_3_out_17_port, CK => CLK, 
                           RN => n37, Q => sum_reg3_17_port, QN => n_1817);
   sum_reg3_reg_18_inst : DFFR_X1 port map( D => sum_3_out_18_port, CK => CLK, 
                           RN => n37, Q => sum_reg3_18_port, QN => n_1818);
   sum_reg3_reg_19_inst : DFFR_X1 port map( D => sum_3_out_19_port, CK => CLK, 
                           RN => n37, Q => sum_reg3_19_port, QN => n_1819);
   sum_reg3_reg_20_inst : DFFR_X1 port map( D => sum_3_out_20_port, CK => CLK, 
                           RN => n37, Q => sum_reg3_20_port, QN => n_1820);
   sum_reg3_reg_21_inst : DFFR_X1 port map( D => sum_3_out_21_port, CK => CLK, 
                           RN => n37, Q => sum_reg3_21_port, QN => n_1821);
   sum_reg3_reg_22_inst : DFFR_X1 port map( D => sum_3_out_22_port, CK => CLK, 
                           RN => n37, Q => sum_reg3_22_port, QN => n_1822);
   sum_reg3_reg_23_inst : DFFR_X1 port map( D => sum_3_out_23_port, CK => CLK, 
                           RN => n37, Q => sum_reg3_23_port, QN => n_1823);
   sum_reg3_reg_24_inst : DFFR_X1 port map( D => sum_3_out_24_port, CK => CLK, 
                           RN => n37, Q => sum_reg3_24_port, QN => n_1824);
   sum_reg3_reg_25_inst : DFFR_X1 port map( D => sum_3_out_25_port, CK => CLK, 
                           RN => n36, Q => sum_reg3_25_port, QN => n_1825);
   sum_reg3_reg_26_inst : DFFR_X1 port map( D => sum_3_out_26_port, CK => CLK, 
                           RN => n36, Q => sum_reg3_26_port, QN => n_1826);
   sum_reg3_reg_27_inst : DFFR_X1 port map( D => sum_3_out_27_port, CK => CLK, 
                           RN => n36, Q => sum_reg3_27_port, QN => n_1827);
   sum_reg3_reg_28_inst : DFFR_X1 port map( D => sum_3_out_28_port, CK => CLK, 
                           RN => n36, Q => sum_reg3_28_port, QN => n_1828);
   sum_reg3_reg_29_inst : DFFR_X1 port map( D => sum_3_out_29_port, CK => CLK, 
                           RN => n36, Q => sum_reg3_29_port, QN => n_1829);
   sum_reg3_reg_30_inst : DFFR_X1 port map( D => sum_3_out_30_port, CK => CLK, 
                           RN => n36, Q => sum_reg3_30_port, QN => n_1830);
   sum_reg3_reg_31_inst : DFFR_X1 port map( D => sum_3_out_31_port, CK => CLK, 
                           RN => n36, Q => sum_reg3_31_port, QN => n_1831);
   sum_reg3_reg_32_inst : DFFR_X1 port map( D => sum_3_out_32_port, CK => CLK, 
                           RN => n36, Q => sum_reg3_32_port, QN => n_1832);
   sum_reg3_reg_33_inst : DFFR_X1 port map( D => sum_3_out_33_port, CK => CLK, 
                           RN => n36, Q => sum_reg3_33_port, QN => n_1833);
   sum_reg3_reg_34_inst : DFFR_X1 port map( D => sum_3_out_34_port, CK => CLK, 
                           RN => n36, Q => sum_reg3_34_port, QN => n_1834);
   sum_reg3_reg_35_inst : DFFR_X1 port map( D => sum_3_out_35_port, CK => CLK, 
                           RN => n36, Q => sum_reg3_35_port, QN => n_1835);
   sum_reg3_reg_36_inst : DFFR_X1 port map( D => sum_3_out_36_port, CK => CLK, 
                           RN => n35, Q => sum_reg3_36_port, QN => n_1836);
   sum_reg3_reg_37_inst : DFFR_X1 port map( D => sum_3_out_37_port, CK => CLK, 
                           RN => n35, Q => sum_reg3_37_port, QN => n_1837);
   sum_reg3_reg_38_inst : DFFR_X1 port map( D => sum_3_out_38_port, CK => CLK, 
                           RN => n35, Q => sum_reg3_38_port, QN => n_1838);
   sum_reg3_reg_39_inst : DFFR_X1 port map( D => sum_3_out_39_port, CK => CLK, 
                           RN => n35, Q => sum_reg3_39_port, QN => n_1839);
   sum_reg3_reg_40_inst : DFFR_X1 port map( D => sum_3_out_40_port, CK => CLK, 
                           RN => n35, Q => sum_reg3_40_port, QN => n_1840);
   sum_reg3_reg_41_inst : DFFR_X1 port map( D => sum_3_out_41_port, CK => CLK, 
                           RN => n35, Q => sum_reg3_41_port, QN => n_1841);
   sum_reg3_reg_42_inst : DFFR_X1 port map( D => sum_3_out_42_port, CK => CLK, 
                           RN => n35, Q => sum_reg3_42_port, QN => n_1842);
   sum_reg3_reg_43_inst : DFFR_X1 port map( D => sum_3_out_43_port, CK => CLK, 
                           RN => n35, Q => sum_reg3_43_port, QN => n_1843);
   sum_reg3_reg_44_inst : DFFR_X1 port map( D => sum_3_out_44_port, CK => CLK, 
                           RN => n35, Q => sum_reg3_44_port, QN => n_1844);
   sum_reg3_reg_45_inst : DFFR_X1 port map( D => sum_3_out_45_port, CK => CLK, 
                           RN => n35, Q => sum_reg3_45_port, QN => n_1845);
   sum_reg3_reg_46_inst : DFFR_X1 port map( D => sum_3_out_46_port, CK => CLK, 
                           RN => n35, Q => sum_reg3_46_port, QN => n_1846);
   sum_reg3_reg_47_inst : DFFR_X1 port map( D => sum_3_out_47_port, CK => CLK, 
                           RN => n34, Q => sum_reg3_47_port, QN => n_1847);
   sum_reg3_reg_48_inst : DFFR_X1 port map( D => sum_3_out_48_port, CK => CLK, 
                           RN => n34, Q => sum_reg3_48_port, QN => n_1848);
   sum_reg3_reg_49_inst : DFFR_X1 port map( D => sum_3_out_49_port, CK => CLK, 
                           RN => n34, Q => sum_reg3_49_port, QN => n_1849);
   sum_reg3_reg_50_inst : DFFR_X1 port map( D => sum_3_out_50_port, CK => CLK, 
                           RN => n34, Q => sum_reg3_50_port, QN => n_1850);
   sum_reg3_reg_51_inst : DFFR_X1 port map( D => sum_3_out_51_port, CK => CLK, 
                           RN => n34, Q => sum_reg3_51_port, QN => n_1851);
   sum_reg3_reg_52_inst : DFFR_X1 port map( D => sum_3_out_52_port, CK => CLK, 
                           RN => n34, Q => sum_reg3_52_port, QN => n_1852);
   sum_reg3_reg_53_inst : DFFR_X1 port map( D => sum_3_out_53_port, CK => CLK, 
                           RN => n34, Q => sum_reg3_53_port, QN => n_1853);
   sum_reg3_reg_54_inst : DFFR_X1 port map( D => sum_3_out_54_port, CK => CLK, 
                           RN => n34, Q => sum_reg3_54_port, QN => n_1854);
   sum_reg3_reg_55_inst : DFFR_X1 port map( D => sum_3_out_55_port, CK => CLK, 
                           RN => n34, Q => sum_reg3_55_port, QN => n_1855);
   sum_reg3_reg_56_inst : DFFR_X1 port map( D => sum_3_out_56_port, CK => CLK, 
                           RN => n34, Q => sum_reg3_56_port, QN => n_1856);
   sum_reg3_reg_57_inst : DFFR_X1 port map( D => sum_3_out_57_port, CK => CLK, 
                           RN => n34, Q => sum_reg3_57_port, QN => n_1857);
   sum_reg3_reg_58_inst : DFFR_X1 port map( D => sum_3_out_58_port, CK => CLK, 
                           RN => n33, Q => sum_reg3_58_port, QN => n_1858);
   sum_reg3_reg_59_inst : DFFR_X1 port map( D => sum_3_out_59_port, CK => CLK, 
                           RN => n33, Q => sum_reg3_59_port, QN => n_1859);
   sum_reg3_reg_60_inst : DFFR_X1 port map( D => sum_3_out_60_port, CK => CLK, 
                           RN => n33, Q => sum_reg3_60_port, QN => n_1860);
   sum_reg3_reg_61_inst : DFFR_X1 port map( D => sum_3_out_61_port, CK => CLK, 
                           RN => n33, Q => sum_reg3_61_port, QN => n_1861);
   sum_reg3_reg_62_inst : DFFR_X1 port map( D => sum_3_out_62_port, CK => CLK, 
                           RN => n33, Q => sum_reg3_62_port, QN => n_1862);
   sum_reg3_reg_63_inst : DFFR_X1 port map( D => sum_3_out_63_port, CK => CLK, 
                           RN => n33, Q => sum_reg3_63_port, QN => n_1863);
   enc_reg31_reg_2_inst : DFFR_X1 port map( D => s_sel_3_2_port, CK => CLK, RN 
                           => n33, Q => enc_reg31_2_port, QN => n_1864);
   enc_reg32_reg_2_inst : DFFR_X1 port map( D => enc_reg31_2_port, CK => CLK, 
                           RN => n33, Q => enc_reg32_2_port, QN => n_1865);
   enc_reg31_reg_1_inst : DFFR_X1 port map( D => s_sel_3_1_port, CK => CLK, RN 
                           => n33, Q => enc_reg31_1_port, QN => n_1866);
   enc_reg32_reg_1_inst : DFFR_X1 port map( D => enc_reg31_1_port, CK => CLK, 
                           RN => n33, Q => enc_reg32_1_port, QN => n_1867);
   enc_reg31_reg_0_inst : DFFR_X1 port map( D => s_sel_3_0_port, CK => CLK, RN 
                           => n33, Q => enc_reg31_0_port, QN => n_1868);
   enc_reg32_reg_0_inst : DFFR_X1 port map( D => enc_reg31_0_port, CK => CLK, 
                           RN => n32, Q => enc_reg32_0_port, QN => n_1869);
   mux_reg3_reg_0_inst : DFFR_X1 port map( D => mux_3_out_0_port, CK => CLK, RN
                           => n32, Q => mux_reg3_0_port, QN => n_1870);
   mux_reg3_reg_1_inst : DFFR_X1 port map( D => mux_3_out_1_port, CK => CLK, RN
                           => n32, Q => mux_reg3_1_port, QN => n_1871);
   mux_reg3_reg_2_inst : DFFR_X1 port map( D => mux_3_out_2_port, CK => CLK, RN
                           => n32, Q => mux_reg3_2_port, QN => n_1872);
   mux_reg3_reg_3_inst : DFFR_X1 port map( D => mux_3_out_3_port, CK => CLK, RN
                           => n32, Q => mux_reg3_3_port, QN => n_1873);
   mux_reg3_reg_4_inst : DFFR_X1 port map( D => mux_3_out_4_port, CK => CLK, RN
                           => n32, Q => mux_reg3_4_port, QN => n_1874);
   mux_reg3_reg_5_inst : DFFR_X1 port map( D => mux_3_out_5_port, CK => CLK, RN
                           => n32, Q => mux_reg3_5_port, QN => n_1875);
   mux_reg3_reg_6_inst : DFFR_X1 port map( D => mux_3_out_6_port, CK => CLK, RN
                           => n32, Q => mux_reg3_6_port, QN => n_1876);
   mux_reg3_reg_7_inst : DFFR_X1 port map( D => mux_3_out_7_port, CK => CLK, RN
                           => n32, Q => mux_reg3_7_port, QN => n_1877);
   mux_reg3_reg_8_inst : DFFR_X1 port map( D => mux_3_out_8_port, CK => CLK, RN
                           => n32, Q => mux_reg3_8_port, QN => n_1878);
   mux_reg3_reg_9_inst : DFFR_X1 port map( D => mux_3_out_9_port, CK => CLK, RN
                           => n32, Q => mux_reg3_9_port, QN => n_1879);
   mux_reg3_reg_10_inst : DFFR_X1 port map( D => mux_3_out_10_port, CK => CLK, 
                           RN => n31, Q => mux_reg3_10_port, QN => n_1880);
   mux_reg3_reg_11_inst : DFFR_X1 port map( D => mux_3_out_11_port, CK => CLK, 
                           RN => n31, Q => mux_reg3_11_port, QN => n_1881);
   mux_reg3_reg_12_inst : DFFR_X1 port map( D => mux_3_out_12_port, CK => CLK, 
                           RN => n31, Q => mux_reg3_12_port, QN => n_1882);
   mux_reg3_reg_13_inst : DFFR_X1 port map( D => mux_3_out_13_port, CK => CLK, 
                           RN => n31, Q => mux_reg3_13_port, QN => n_1883);
   mux_reg3_reg_14_inst : DFFR_X1 port map( D => mux_3_out_14_port, CK => CLK, 
                           RN => n31, Q => mux_reg3_14_port, QN => n_1884);
   mux_reg3_reg_15_inst : DFFR_X1 port map( D => mux_3_out_15_port, CK => CLK, 
                           RN => n31, Q => mux_reg3_15_port, QN => n_1885);
   mux_reg3_reg_16_inst : DFFR_X1 port map( D => mux_3_out_16_port, CK => CLK, 
                           RN => n31, Q => mux_reg3_16_port, QN => n_1886);
   mux_reg3_reg_17_inst : DFFR_X1 port map( D => mux_3_out_17_port, CK => CLK, 
                           RN => n31, Q => mux_reg3_17_port, QN => n_1887);
   mux_reg3_reg_18_inst : DFFR_X1 port map( D => mux_3_out_18_port, CK => CLK, 
                           RN => n31, Q => mux_reg3_18_port, QN => n_1888);
   mux_reg3_reg_19_inst : DFFR_X1 port map( D => mux_3_out_19_port, CK => CLK, 
                           RN => n31, Q => mux_reg3_19_port, QN => n_1889);
   mux_reg3_reg_20_inst : DFFR_X1 port map( D => mux_3_out_20_port, CK => CLK, 
                           RN => n31, Q => mux_reg3_20_port, QN => n_1890);
   mux_reg3_reg_21_inst : DFFR_X1 port map( D => mux_3_out_21_port, CK => CLK, 
                           RN => n30, Q => mux_reg3_21_port, QN => n_1891);
   mux_reg3_reg_22_inst : DFFR_X1 port map( D => mux_3_out_22_port, CK => CLK, 
                           RN => n30, Q => mux_reg3_22_port, QN => n_1892);
   mux_reg3_reg_23_inst : DFFR_X1 port map( D => mux_3_out_23_port, CK => CLK, 
                           RN => n30, Q => mux_reg3_23_port, QN => n_1893);
   mux_reg3_reg_24_inst : DFFR_X1 port map( D => mux_3_out_24_port, CK => CLK, 
                           RN => n30, Q => mux_reg3_24_port, QN => n_1894);
   mux_reg3_reg_25_inst : DFFR_X1 port map( D => mux_3_out_25_port, CK => CLK, 
                           RN => n30, Q => mux_reg3_25_port, QN => n_1895);
   mux_reg3_reg_26_inst : DFFR_X1 port map( D => mux_3_out_26_port, CK => CLK, 
                           RN => n30, Q => mux_reg3_26_port, QN => n_1896);
   mux_reg3_reg_27_inst : DFFR_X1 port map( D => mux_3_out_27_port, CK => CLK, 
                           RN => n30, Q => mux_reg3_27_port, QN => n_1897);
   mux_reg3_reg_28_inst : DFFR_X1 port map( D => mux_3_out_28_port, CK => CLK, 
                           RN => n30, Q => mux_reg3_28_port, QN => n_1898);
   mux_reg3_reg_29_inst : DFFR_X1 port map( D => mux_3_out_29_port, CK => CLK, 
                           RN => n30, Q => mux_reg3_29_port, QN => n_1899);
   mux_reg3_reg_30_inst : DFFR_X1 port map( D => mux_3_out_30_port, CK => CLK, 
                           RN => n30, Q => mux_reg3_30_port, QN => n_1900);
   mux_reg3_reg_31_inst : DFFR_X1 port map( D => mux_3_out_31_port, CK => CLK, 
                           RN => n30, Q => mux_reg3_31_port, QN => n_1901);
   enc_0 : enc33_0 port map( A(2) => B(1), A(1) => B(0), A(0) => X_Logic0_port,
                           Y(2) => s_sel_0_2_port, Y(1) => s_sel_0_1_port, Y(0)
                           => s_sel_0_0_port);
   enc_1 : enc33_3 port map( A(2) => B(3), A(1) => B(2), A(0) => B(1), Y(2) => 
                           s_sel_1_2_port, Y(1) => s_sel_1_1_port, Y(0) => 
                           s_sel_1_0_port);
   enc_2 : enc33_2 port map( A(2) => B(5), A(1) => B(4), A(0) => B(3), Y(2) => 
                           s_sel_2_2_port, Y(1) => s_sel_2_1_port, Y(0) => 
                           s_sel_2_0_port);
   enc_3 : enc33_1 port map( A(2) => B(7), A(1) => B(6), A(0) => B(5), Y(2) => 
                           s_sel_3_2_port, Y(1) => s_sel_3_1_port, Y(0) => 
                           s_sel_3_0_port);
   shift2A : shl1_NBIT32_0 port map( A(31) => n18, A(30) => A(30), A(29) => 
                           A(29), A(28) => A(28), A(27) => A(27), A(26) => 
                           A(26), A(25) => A(25), A(24) => A(24), A(23) => 
                           A(23), A(22) => A(22), A(21) => A(21), A(20) => 
                           A(20), A(19) => A(19), A(18) => A(18), A(17) => 
                           A(17), A(16) => A(16), A(15) => A(15), A(14) => 
                           A(14), A(13) => A(13), A(12) => A(12), A(11) => 
                           A(11), A(10) => A(10), A(9) => A(9), A(8) => A(8), 
                           A(7) => A(7), A(6) => A(6), A(5) => A(5), A(4) => 
                           A(4), A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), Y(31) => s_2A_1_31_port, Y(30) => 
                           s_2A_1_30_port, Y(29) => s_2A_1_29_port, Y(28) => 
                           s_2A_1_28_port, Y(27) => s_2A_1_27_port, Y(26) => 
                           s_2A_1_26_port, Y(25) => s_2A_1_25_port, Y(24) => 
                           s_2A_1_24_port, Y(23) => s_2A_1_23_port, Y(22) => 
                           s_2A_1_22_port, Y(21) => s_2A_1_21_port, Y(20) => 
                           s_2A_1_20_port, Y(19) => s_2A_1_19_port, Y(18) => 
                           s_2A_1_18_port, Y(17) => s_2A_1_17_port, Y(16) => 
                           s_2A_1_16_port, Y(15) => s_2A_1_15_port, Y(14) => 
                           s_2A_1_14_port, Y(13) => s_2A_1_13_port, Y(12) => 
                           s_2A_1_12_port, Y(11) => s_2A_1_11_port, Y(10) => 
                           s_2A_1_10_port, Y(9) => s_2A_1_9_port, Y(8) => 
                           s_2A_1_8_port, Y(7) => s_2A_1_7_port, Y(6) => 
                           s_2A_1_6_port, Y(5) => s_2A_1_5_port, Y(4) => 
                           s_2A_1_4_port, Y(3) => s_2A_1_3_port, Y(2) => 
                           s_2A_1_2_port, Y(1) => s_2A_1_1_port, Y(0) => n_1902
                           );
   shift4A : shl2_NBIT32_0 port map( A(31) => n18, A(30) => A(30), A(29) => 
                           A(29), A(28) => A(28), A(27) => A(27), A(26) => 
                           A(26), A(25) => A(25), A(24) => A(24), A(23) => 
                           A(23), A(22) => A(22), A(21) => A(21), A(20) => 
                           A(20), A(19) => A(19), A(18) => A(18), A(17) => 
                           A(17), A(16) => A(16), A(15) => A(15), A(14) => 
                           A(14), A(13) => A(13), A(12) => A(12), A(11) => 
                           A(11), A(10) => A(10), A(9) => A(9), A(8) => A(8), 
                           A(7) => A(7), A(6) => A(6), A(5) => A(5), A(4) => 
                           A(4), A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), Y(31) => s_4A_1_31_port, Y(30) => 
                           s_4A_1_30_port, Y(29) => s_4A_1_29_port, Y(28) => 
                           s_4A_1_28_port, Y(27) => s_4A_1_27_port, Y(26) => 
                           s_4A_1_26_port, Y(25) => s_4A_1_25_port, Y(24) => 
                           s_4A_1_24_port, Y(23) => s_4A_1_23_port, Y(22) => 
                           s_4A_1_22_port, Y(21) => s_4A_1_21_port, Y(20) => 
                           s_4A_1_20_port, Y(19) => s_4A_1_19_port, Y(18) => 
                           s_4A_1_18_port, Y(17) => s_4A_1_17_port, Y(16) => 
                           s_4A_1_16_port, Y(15) => s_4A_1_15_port, Y(14) => 
                           s_4A_1_14_port, Y(13) => s_4A_1_13_port, Y(12) => 
                           s_4A_1_12_port, Y(11) => s_4A_1_11_port, Y(10) => 
                           s_4A_1_10_port, Y(9) => s_4A_1_9_port, Y(8) => 
                           s_4A_1_8_port, Y(7) => s_4A_1_7_port, Y(6) => 
                           s_4A_1_6_port, Y(5) => s_4A_1_5_port, Y(4) => 
                           s_4A_1_4_port, Y(3) => s_4A_1_3_port, Y(2) => 
                           s_4A_1_2_port, Y(1) => n_1903, Y(0) => n_1904);
   shift8A : shl3_NBIT32 port map( A(31) => n18, A(30) => A(30), A(29) => A(29)
                           , A(28) => A(28), A(27) => A(27), A(26) => A(26), 
                           A(25) => A(25), A(24) => A(24), A(23) => A(23), 
                           A(22) => A(22), A(21) => A(21), A(20) => A(20), 
                           A(19) => A(19), A(18) => A(18), A(17) => A(17), 
                           A(16) => A(16), A(15) => A(15), A(14) => A(14), 
                           A(13) => A(13), A(12) => A(12), A(11) => A(11), 
                           A(10) => A(10), A(9) => A(9), A(8) => A(8), A(7) => 
                           A(7), A(6) => A(6), A(5) => A(5), A(4) => A(4), A(3)
                           => A(3), A(2) => A(2), A(1) => A(1), A(0) => A(0), 
                           Y(31) => s_8A_1_31_port, Y(30) => s_8A_1_30_port, 
                           Y(29) => s_8A_1_29_port, Y(28) => s_8A_1_28_port, 
                           Y(27) => s_8A_1_27_port, Y(26) => s_8A_1_26_port, 
                           Y(25) => s_8A_1_25_port, Y(24) => s_8A_1_24_port, 
                           Y(23) => s_8A_1_23_port, Y(22) => s_8A_1_22_port, 
                           Y(21) => s_8A_1_21_port, Y(20) => s_8A_1_20_port, 
                           Y(19) => s_8A_1_19_port, Y(18) => s_8A_1_18_port, 
                           Y(17) => s_8A_1_17_port, Y(16) => s_8A_1_16_port, 
                           Y(15) => s_8A_1_15_port, Y(14) => s_8A_1_14_port, 
                           Y(13) => s_8A_1_13_port, Y(12) => s_8A_1_12_port, 
                           Y(11) => s_8A_1_11_port, Y(10) => s_8A_1_10_port, 
                           Y(9) => s_8A_1_9_port, Y(8) => s_8A_1_8_port, Y(7) 
                           => s_8A_1_7_port, Y(6) => s_8A_1_6_port, Y(5) => 
                           s_8A_1_5_port, Y(4) => s_8A_1_4_port, Y(3) => 
                           s_8A_1_3_port, Y(2) => n_1905, Y(1) => n_1906, Y(0) 
                           => n_1907);
   neg1 : negate_NBIT32_0 port map( A(31) => n18, A(30) => A(30), A(29) => 
                           A(29), A(28) => A(28), A(27) => A(27), A(26) => 
                           A(26), A(25) => A(25), A(24) => A(24), A(23) => 
                           A(23), A(22) => A(22), A(21) => A(21), A(20) => 
                           A(20), A(19) => A(19), A(18) => A(18), A(17) => 
                           A(17), A(16) => A(16), A(15) => A(15), A(14) => 
                           A(14), A(13) => A(13), A(12) => A(12), A(11) => 
                           A(11), A(10) => A(10), A(9) => A(9), A(8) => A(8), 
                           A(7) => A(7), A(6) => A(6), A(5) => A(5), A(4) => 
                           A(4), A(3) => A(3), A(2) => A(2), A(1) => A(1), A(0)
                           => A(0), Y(31) => s_A_neg_31_port, Y(30) => 
                           s_A_neg_30_port, Y(29) => s_A_neg_29_port, Y(28) => 
                           s_A_neg_28_port, Y(27) => s_A_neg_27_port, Y(26) => 
                           s_A_neg_26_port, Y(25) => s_A_neg_25_port, Y(24) => 
                           s_A_neg_24_port, Y(23) => s_A_neg_23_port, Y(22) => 
                           s_A_neg_22_port, Y(21) => s_A_neg_21_port, Y(20) => 
                           s_A_neg_20_port, Y(19) => s_A_neg_19_port, Y(18) => 
                           s_A_neg_18_port, Y(17) => s_A_neg_17_port, Y(16) => 
                           s_A_neg_16_port, Y(15) => s_A_neg_15_port, Y(14) => 
                           s_A_neg_14_port, Y(13) => s_A_neg_13_port, Y(12) => 
                           s_A_neg_12_port, Y(11) => s_A_neg_11_port, Y(10) => 
                           s_A_neg_10_port, Y(9) => s_A_neg_9_port, Y(8) => 
                           s_A_neg_8_port, Y(7) => s_A_neg_7_port, Y(6) => 
                           s_A_neg_6_port, Y(5) => s_A_neg_5_port, Y(4) => 
                           s_A_neg_4_port, Y(3) => s_A_neg_3_port, Y(2) => 
                           s_A_neg_2_port, Y(1) => s_A_neg_1_port, Y(0) => 
                           s_A_neg_0_port);
   neg2 : negate_NBIT32_7 port map( A(31) => s_2A_1_31_port, A(30) => 
                           s_2A_1_30_port, A(29) => s_2A_1_29_port, A(28) => 
                           s_2A_1_28_port, A(27) => s_2A_1_27_port, A(26) => 
                           s_2A_1_26_port, A(25) => s_2A_1_25_port, A(24) => 
                           s_2A_1_24_port, A(23) => s_2A_1_23_port, A(22) => 
                           s_2A_1_22_port, A(21) => s_2A_1_21_port, A(20) => 
                           s_2A_1_20_port, A(19) => s_2A_1_19_port, A(18) => 
                           s_2A_1_18_port, A(17) => s_2A_1_17_port, A(16) => 
                           s_2A_1_16_port, A(15) => s_2A_1_15_port, A(14) => 
                           s_2A_1_14_port, A(13) => s_2A_1_13_port, A(12) => 
                           s_2A_1_12_port, A(11) => s_2A_1_11_port, A(10) => 
                           s_2A_1_10_port, A(9) => s_2A_1_9_port, A(8) => 
                           s_2A_1_8_port, A(7) => s_2A_1_7_port, A(6) => 
                           s_2A_1_6_port, A(5) => s_2A_1_5_port, A(4) => 
                           s_2A_1_4_port, A(3) => s_2A_1_3_port, A(2) => 
                           s_2A_1_2_port, A(1) => s_2A_1_1_port, A(0) => 
                           s_2A_1_0_port, Y(31) => s_2A_1_neg_31_port, Y(30) =>
                           s_2A_1_neg_30_port, Y(29) => s_2A_1_neg_29_port, 
                           Y(28) => s_2A_1_neg_28_port, Y(27) => 
                           s_2A_1_neg_27_port, Y(26) => s_2A_1_neg_26_port, 
                           Y(25) => s_2A_1_neg_25_port, Y(24) => 
                           s_2A_1_neg_24_port, Y(23) => s_2A_1_neg_23_port, 
                           Y(22) => s_2A_1_neg_22_port, Y(21) => 
                           s_2A_1_neg_21_port, Y(20) => s_2A_1_neg_20_port, 
                           Y(19) => s_2A_1_neg_19_port, Y(18) => 
                           s_2A_1_neg_18_port, Y(17) => s_2A_1_neg_17_port, 
                           Y(16) => s_2A_1_neg_16_port, Y(15) => 
                           s_2A_1_neg_15_port, Y(14) => s_2A_1_neg_14_port, 
                           Y(13) => s_2A_1_neg_13_port, Y(12) => 
                           s_2A_1_neg_12_port, Y(11) => s_2A_1_neg_11_port, 
                           Y(10) => s_2A_1_neg_10_port, Y(9) => 
                           s_2A_1_neg_9_port, Y(8) => s_2A_1_neg_8_port, Y(7) 
                           => s_2A_1_neg_7_port, Y(6) => s_2A_1_neg_6_port, 
                           Y(5) => s_2A_1_neg_5_port, Y(4) => s_2A_1_neg_4_port
                           , Y(3) => s_2A_1_neg_3_port, Y(2) => 
                           s_2A_1_neg_2_port, Y(1) => s_2A_1_neg_1_port, Y(0) 
                           => s_2A_1_neg_0_port);
   neg3 : negate_NBIT32_6 port map( A(31) => s_4A_1_31_port, A(30) => 
                           s_4A_1_30_port, A(29) => s_4A_1_29_port, A(28) => 
                           s_4A_1_28_port, A(27) => s_4A_1_27_port, A(26) => 
                           s_4A_1_26_port, A(25) => s_4A_1_25_port, A(24) => 
                           s_4A_1_24_port, A(23) => s_4A_1_23_port, A(22) => 
                           s_4A_1_22_port, A(21) => s_4A_1_21_port, A(20) => 
                           s_4A_1_20_port, A(19) => s_4A_1_19_port, A(18) => 
                           s_4A_1_18_port, A(17) => s_4A_1_17_port, A(16) => 
                           s_4A_1_16_port, A(15) => s_4A_1_15_port, A(14) => 
                           s_4A_1_14_port, A(13) => s_4A_1_13_port, A(12) => 
                           s_4A_1_12_port, A(11) => s_4A_1_11_port, A(10) => 
                           s_4A_1_10_port, A(9) => s_4A_1_9_port, A(8) => 
                           s_4A_1_8_port, A(7) => s_4A_1_7_port, A(6) => 
                           s_4A_1_6_port, A(5) => s_4A_1_5_port, A(4) => 
                           s_4A_1_4_port, A(3) => s_4A_1_3_port, A(2) => 
                           s_4A_1_2_port, A(1) => s_4A_1_1_port, A(0) => 
                           s_4A_1_0_port, Y(31) => s_4A_1_neg_31_port, Y(30) =>
                           s_4A_1_neg_30_port, Y(29) => s_4A_1_neg_29_port, 
                           Y(28) => s_4A_1_neg_28_port, Y(27) => 
                           s_4A_1_neg_27_port, Y(26) => s_4A_1_neg_26_port, 
                           Y(25) => s_4A_1_neg_25_port, Y(24) => 
                           s_4A_1_neg_24_port, Y(23) => s_4A_1_neg_23_port, 
                           Y(22) => s_4A_1_neg_22_port, Y(21) => 
                           s_4A_1_neg_21_port, Y(20) => s_4A_1_neg_20_port, 
                           Y(19) => s_4A_1_neg_19_port, Y(18) => 
                           s_4A_1_neg_18_port, Y(17) => s_4A_1_neg_17_port, 
                           Y(16) => s_4A_1_neg_16_port, Y(15) => 
                           s_4A_1_neg_15_port, Y(14) => s_4A_1_neg_14_port, 
                           Y(13) => s_4A_1_neg_13_port, Y(12) => 
                           s_4A_1_neg_12_port, Y(11) => s_4A_1_neg_11_port, 
                           Y(10) => s_4A_1_neg_10_port, Y(9) => 
                           s_4A_1_neg_9_port, Y(8) => s_4A_1_neg_8_port, Y(7) 
                           => s_4A_1_neg_7_port, Y(6) => s_4A_1_neg_6_port, 
                           Y(5) => s_4A_1_neg_5_port, Y(4) => s_4A_1_neg_4_port
                           , Y(3) => s_4A_1_neg_3_port, Y(2) => 
                           s_4A_1_neg_2_port, Y(1) => s_4A_1_neg_1_port, Y(0) 
                           => s_4A_1_neg_0_port);
   neg4 : negate_NBIT32_5 port map( A(31) => s_8A_1_31_port, A(30) => 
                           s_8A_1_30_port, A(29) => s_8A_1_29_port, A(28) => 
                           s_8A_1_28_port, A(27) => s_8A_1_27_port, A(26) => 
                           s_8A_1_26_port, A(25) => s_8A_1_25_port, A(24) => 
                           s_8A_1_24_port, A(23) => s_8A_1_23_port, A(22) => 
                           s_8A_1_22_port, A(21) => s_8A_1_21_port, A(20) => 
                           s_8A_1_20_port, A(19) => s_8A_1_19_port, A(18) => 
                           s_8A_1_18_port, A(17) => s_8A_1_17_port, A(16) => 
                           s_8A_1_16_port, A(15) => s_8A_1_15_port, A(14) => 
                           s_8A_1_14_port, A(13) => s_8A_1_13_port, A(12) => 
                           s_8A_1_12_port, A(11) => s_8A_1_11_port, A(10) => 
                           s_8A_1_10_port, A(9) => s_8A_1_9_port, A(8) => 
                           s_8A_1_8_port, A(7) => s_8A_1_7_port, A(6) => 
                           s_8A_1_6_port, A(5) => s_8A_1_5_port, A(4) => 
                           s_8A_1_4_port, A(3) => s_8A_1_3_port, A(2) => 
                           s_8A_1_2_port, A(1) => s_8A_1_1_port, A(0) => 
                           s_8A_1_0_port, Y(31) => s_8A_1_neg_31_port, Y(30) =>
                           s_8A_1_neg_30_port, Y(29) => s_8A_1_neg_29_port, 
                           Y(28) => s_8A_1_neg_28_port, Y(27) => 
                           s_8A_1_neg_27_port, Y(26) => s_8A_1_neg_26_port, 
                           Y(25) => s_8A_1_neg_25_port, Y(24) => 
                           s_8A_1_neg_24_port, Y(23) => s_8A_1_neg_23_port, 
                           Y(22) => s_8A_1_neg_22_port, Y(21) => 
                           s_8A_1_neg_21_port, Y(20) => s_8A_1_neg_20_port, 
                           Y(19) => s_8A_1_neg_19_port, Y(18) => 
                           s_8A_1_neg_18_port, Y(17) => s_8A_1_neg_17_port, 
                           Y(16) => s_8A_1_neg_16_port, Y(15) => 
                           s_8A_1_neg_15_port, Y(14) => s_8A_1_neg_14_port, 
                           Y(13) => s_8A_1_neg_13_port, Y(12) => 
                           s_8A_1_neg_12_port, Y(11) => s_8A_1_neg_11_port, 
                           Y(10) => s_8A_1_neg_10_port, Y(9) => 
                           s_8A_1_neg_9_port, Y(8) => s_8A_1_neg_8_port, Y(7) 
                           => s_8A_1_neg_7_port, Y(6) => s_8A_1_neg_6_port, 
                           Y(5) => s_8A_1_neg_5_port, Y(4) => s_8A_1_neg_4_port
                           , Y(3) => s_8A_1_neg_3_port, Y(2) => 
                           s_8A_1_neg_2_port, Y(1) => s_8A_1_neg_1_port, Y(0) 
                           => s_8A_1_neg_0_port);
   mux1 : mux51_gen_NBIT32_0 port map( A0(31) => X_Logic0_port, A0(30) => 
                           X_Logic0_port, A0(29) => X_Logic0_port, A0(28) => 
                           X_Logic0_port, A0(27) => X_Logic0_port, A0(26) => 
                           X_Logic0_port, A0(25) => X_Logic0_port, A0(24) => 
                           X_Logic0_port, A0(23) => X_Logic0_port, A0(22) => 
                           X_Logic0_port, A0(21) => X_Logic0_port, A0(20) => 
                           X_Logic0_port, A0(19) => X_Logic0_port, A0(18) => 
                           X_Logic0_port, A0(17) => X_Logic0_port, A0(16) => 
                           X_Logic0_port, A0(15) => X_Logic0_port, A0(14) => 
                           X_Logic0_port, A0(13) => X_Logic0_port, A0(12) => 
                           X_Logic0_port, A0(11) => X_Logic0_port, A0(10) => 
                           X_Logic0_port, A0(9) => X_Logic0_port, A0(8) => 
                           X_Logic0_port, A0(7) => X_Logic0_port, A0(6) => 
                           X_Logic0_port, A0(5) => X_Logic0_port, A0(4) => 
                           X_Logic0_port, A0(3) => X_Logic0_port, A0(2) => 
                           X_Logic0_port, A0(1) => X_Logic0_port, A0(0) => 
                           X_Logic0_port, A1(31) => n18, A1(30) => A(30), 
                           A1(29) => A(29), A1(28) => A(28), A1(27) => A(27), 
                           A1(26) => A(26), A1(25) => A(25), A1(24) => A(24), 
                           A1(23) => A(23), A1(22) => A(22), A1(21) => A(21), 
                           A1(20) => A(20), A1(19) => A(19), A1(18) => A(18), 
                           A1(17) => A(17), A1(16) => A(16), A1(15) => A(15), 
                           A1(14) => A(14), A1(13) => A(13), A1(12) => A(12), 
                           A1(11) => A(11), A1(10) => A(10), A1(9) => A(9), 
                           A1(8) => A(8), A1(7) => A(7), A1(6) => A(6), A1(5) 
                           => A(5), A1(4) => A(4), A1(3) => A(3), A1(2) => A(2)
                           , A1(1) => A(1), A1(0) => A(0), A2(31) => 
                           s_A_neg_31_port, A2(30) => s_A_neg_30_port, A2(29) 
                           => s_A_neg_29_port, A2(28) => s_A_neg_28_port, 
                           A2(27) => s_A_neg_27_port, A2(26) => s_A_neg_26_port
                           , A2(25) => s_A_neg_25_port, A2(24) => 
                           s_A_neg_24_port, A2(23) => s_A_neg_23_port, A2(22) 
                           => s_A_neg_22_port, A2(21) => s_A_neg_21_port, 
                           A2(20) => s_A_neg_20_port, A2(19) => s_A_neg_19_port
                           , A2(18) => s_A_neg_18_port, A2(17) => 
                           s_A_neg_17_port, A2(16) => s_A_neg_16_port, A2(15) 
                           => s_A_neg_15_port, A2(14) => s_A_neg_14_port, 
                           A2(13) => s_A_neg_13_port, A2(12) => s_A_neg_12_port
                           , A2(11) => s_A_neg_11_port, A2(10) => 
                           s_A_neg_10_port, A2(9) => s_A_neg_9_port, A2(8) => 
                           s_A_neg_8_port, A2(7) => s_A_neg_7_port, A2(6) => 
                           s_A_neg_6_port, A2(5) => s_A_neg_5_port, A2(4) => 
                           s_A_neg_4_port, A2(3) => s_A_neg_3_port, A2(2) => 
                           s_A_neg_2_port, A2(1) => s_A_neg_1_port, A2(0) => 
                           s_A_neg_0_port, A3(31) => s_2A_1_31_port, A3(30) => 
                           s_2A_1_30_port, A3(29) => s_2A_1_29_port, A3(28) => 
                           s_2A_1_28_port, A3(27) => s_2A_1_27_port, A3(26) => 
                           s_2A_1_26_port, A3(25) => s_2A_1_25_port, A3(24) => 
                           s_2A_1_24_port, A3(23) => s_2A_1_23_port, A3(22) => 
                           s_2A_1_22_port, A3(21) => s_2A_1_21_port, A3(20) => 
                           s_2A_1_20_port, A3(19) => s_2A_1_19_port, A3(18) => 
                           s_2A_1_18_port, A3(17) => s_2A_1_17_port, A3(16) => 
                           s_2A_1_16_port, A3(15) => s_2A_1_15_port, A3(14) => 
                           s_2A_1_14_port, A3(13) => s_2A_1_13_port, A3(12) => 
                           s_2A_1_12_port, A3(11) => s_2A_1_11_port, A3(10) => 
                           s_2A_1_10_port, A3(9) => s_2A_1_9_port, A3(8) => 
                           s_2A_1_8_port, A3(7) => s_2A_1_7_port, A3(6) => 
                           s_2A_1_6_port, A3(5) => s_2A_1_5_port, A3(4) => 
                           s_2A_1_4_port, A3(3) => s_2A_1_3_port, A3(2) => 
                           s_2A_1_2_port, A3(1) => s_2A_1_1_port, A3(0) => 
                           s_2A_1_0_port, A4(31) => s_2A_1_neg_31_port, A4(30) 
                           => s_2A_1_neg_30_port, A4(29) => s_2A_1_neg_29_port,
                           A4(28) => s_2A_1_neg_28_port, A4(27) => 
                           s_2A_1_neg_27_port, A4(26) => s_2A_1_neg_26_port, 
                           A4(25) => s_2A_1_neg_25_port, A4(24) => 
                           s_2A_1_neg_24_port, A4(23) => s_2A_1_neg_23_port, 
                           A4(22) => s_2A_1_neg_22_port, A4(21) => 
                           s_2A_1_neg_21_port, A4(20) => s_2A_1_neg_20_port, 
                           A4(19) => s_2A_1_neg_19_port, A4(18) => 
                           s_2A_1_neg_18_port, A4(17) => s_2A_1_neg_17_port, 
                           A4(16) => s_2A_1_neg_16_port, A4(15) => 
                           s_2A_1_neg_15_port, A4(14) => s_2A_1_neg_14_port, 
                           A4(13) => s_2A_1_neg_13_port, A4(12) => 
                           s_2A_1_neg_12_port, A4(11) => s_2A_1_neg_11_port, 
                           A4(10) => s_2A_1_neg_10_port, A4(9) => 
                           s_2A_1_neg_9_port, A4(8) => s_2A_1_neg_8_port, A4(7)
                           => s_2A_1_neg_7_port, A4(6) => s_2A_1_neg_6_port, 
                           A4(5) => s_2A_1_neg_5_port, A4(4) => 
                           s_2A_1_neg_4_port, A4(3) => s_2A_1_neg_3_port, A4(2)
                           => s_2A_1_neg_2_port, A4(1) => s_2A_1_neg_1_port, 
                           A4(0) => s_2A_1_neg_0_port, SEL(2) => s_sel_0_2_port
                           , SEL(1) => s_sel_0_1_port, SEL(0) => s_sel_0_0_port
                           , Y(31) => mux1_out_31_port, Y(30) => 
                           mux1_out_30_port, Y(29) => mux1_out_29_port, Y(28) 
                           => mux1_out_28_port, Y(27) => mux1_out_27_port, 
                           Y(26) => mux1_out_26_port, Y(25) => mux1_out_25_port
                           , Y(24) => mux1_out_24_port, Y(23) => 
                           mux1_out_23_port, Y(22) => mux1_out_22_port, Y(21) 
                           => mux1_out_21_port, Y(20) => mux1_out_20_port, 
                           Y(19) => mux1_out_19_port, Y(18) => mux1_out_18_port
                           , Y(17) => mux1_out_17_port, Y(16) => 
                           mux1_out_16_port, Y(15) => mux1_out_15_port, Y(14) 
                           => mux1_out_14_port, Y(13) => mux1_out_13_port, 
                           Y(12) => mux1_out_12_port, Y(11) => mux1_out_11_port
                           , Y(10) => mux1_out_10_port, Y(9) => mux1_out_9_port
                           , Y(8) => mux1_out_8_port, Y(7) => mux1_out_7_port, 
                           Y(6) => mux1_out_6_port, Y(5) => mux1_out_5_port, 
                           Y(4) => mux1_out_4_port, Y(3) => mux1_out_3_port, 
                           Y(2) => mux1_out_2_port, Y(1) => mux1_out_1_port, 
                           Y(0) => mux1_out_0_port);
   mux2 : mux51_gen_NBIT32_3 port map( A0(31) => X_Logic0_port, A0(30) => 
                           X_Logic0_port, A0(29) => X_Logic0_port, A0(28) => 
                           X_Logic0_port, A0(27) => X_Logic0_port, A0(26) => 
                           X_Logic0_port, A0(25) => X_Logic0_port, A0(24) => 
                           X_Logic0_port, A0(23) => X_Logic0_port, A0(22) => 
                           X_Logic0_port, A0(21) => X_Logic0_port, A0(20) => 
                           X_Logic0_port, A0(19) => X_Logic0_port, A0(18) => 
                           X_Logic0_port, A0(17) => X_Logic0_port, A0(16) => 
                           X_Logic0_port, A0(15) => X_Logic0_port, A0(14) => 
                           X_Logic0_port, A0(13) => X_Logic0_port, A0(12) => 
                           X_Logic0_port, A0(11) => X_Logic0_port, A0(10) => 
                           X_Logic0_port, A0(9) => X_Logic0_port, A0(8) => 
                           X_Logic0_port, A0(7) => X_Logic0_port, A0(6) => 
                           X_Logic0_port, A0(5) => X_Logic0_port, A0(4) => 
                           X_Logic0_port, A0(3) => X_Logic0_port, A0(2) => 
                           X_Logic0_port, A0(1) => X_Logic0_port, A0(0) => 
                           X_Logic0_port, A1(31) => s_4A_1_31_port, A1(30) => 
                           s_4A_1_30_port, A1(29) => s_4A_1_29_port, A1(28) => 
                           s_4A_1_28_port, A1(27) => s_4A_1_27_port, A1(26) => 
                           s_4A_1_26_port, A1(25) => s_4A_1_25_port, A1(24) => 
                           s_4A_1_24_port, A1(23) => s_4A_1_23_port, A1(22) => 
                           s_4A_1_22_port, A1(21) => s_4A_1_21_port, A1(20) => 
                           s_4A_1_20_port, A1(19) => s_4A_1_19_port, A1(18) => 
                           s_4A_1_18_port, A1(17) => s_4A_1_17_port, A1(16) => 
                           s_4A_1_16_port, A1(15) => s_4A_1_15_port, A1(14) => 
                           s_4A_1_14_port, A1(13) => s_4A_1_13_port, A1(12) => 
                           s_4A_1_12_port, A1(11) => s_4A_1_11_port, A1(10) => 
                           s_4A_1_10_port, A1(9) => s_4A_1_9_port, A1(8) => 
                           s_4A_1_8_port, A1(7) => s_4A_1_7_port, A1(6) => 
                           s_4A_1_6_port, A1(5) => s_4A_1_5_port, A1(4) => 
                           s_4A_1_4_port, A1(3) => s_4A_1_3_port, A1(2) => 
                           s_4A_1_2_port, A1(1) => s_4A_1_1_port, A1(0) => 
                           s_4A_1_0_port, A2(31) => s_4A_1_neg_31_port, A2(30) 
                           => s_4A_1_neg_30_port, A2(29) => s_4A_1_neg_29_port,
                           A2(28) => s_4A_1_neg_28_port, A2(27) => 
                           s_4A_1_neg_27_port, A2(26) => s_4A_1_neg_26_port, 
                           A2(25) => s_4A_1_neg_25_port, A2(24) => 
                           s_4A_1_neg_24_port, A2(23) => s_4A_1_neg_23_port, 
                           A2(22) => s_4A_1_neg_22_port, A2(21) => 
                           s_4A_1_neg_21_port, A2(20) => s_4A_1_neg_20_port, 
                           A2(19) => s_4A_1_neg_19_port, A2(18) => 
                           s_4A_1_neg_18_port, A2(17) => s_4A_1_neg_17_port, 
                           A2(16) => s_4A_1_neg_16_port, A2(15) => 
                           s_4A_1_neg_15_port, A2(14) => s_4A_1_neg_14_port, 
                           A2(13) => s_4A_1_neg_13_port, A2(12) => 
                           s_4A_1_neg_12_port, A2(11) => s_4A_1_neg_11_port, 
                           A2(10) => s_4A_1_neg_10_port, A2(9) => 
                           s_4A_1_neg_9_port, A2(8) => s_4A_1_neg_8_port, A2(7)
                           => s_4A_1_neg_7_port, A2(6) => s_4A_1_neg_6_port, 
                           A2(5) => s_4A_1_neg_5_port, A2(4) => 
                           s_4A_1_neg_4_port, A2(3) => s_4A_1_neg_3_port, A2(2)
                           => s_4A_1_neg_2_port, A2(1) => s_4A_1_neg_1_port, 
                           A2(0) => s_4A_1_neg_0_port, A3(31) => s_8A_1_31_port
                           , A3(30) => s_8A_1_30_port, A3(29) => s_8A_1_29_port
                           , A3(28) => s_8A_1_28_port, A3(27) => s_8A_1_27_port
                           , A3(26) => s_8A_1_26_port, A3(25) => s_8A_1_25_port
                           , A3(24) => s_8A_1_24_port, A3(23) => s_8A_1_23_port
                           , A3(22) => s_8A_1_22_port, A3(21) => s_8A_1_21_port
                           , A3(20) => s_8A_1_20_port, A3(19) => s_8A_1_19_port
                           , A3(18) => s_8A_1_18_port, A3(17) => s_8A_1_17_port
                           , A3(16) => s_8A_1_16_port, A3(15) => s_8A_1_15_port
                           , A3(14) => s_8A_1_14_port, A3(13) => s_8A_1_13_port
                           , A3(12) => s_8A_1_12_port, A3(11) => s_8A_1_11_port
                           , A3(10) => s_8A_1_10_port, A3(9) => s_8A_1_9_port, 
                           A3(8) => s_8A_1_8_port, A3(7) => s_8A_1_7_port, 
                           A3(6) => s_8A_1_6_port, A3(5) => s_8A_1_5_port, 
                           A3(4) => s_8A_1_4_port, A3(3) => s_8A_1_3_port, 
                           A3(2) => s_8A_1_2_port, A3(1) => s_8A_1_1_port, 
                           A3(0) => s_8A_1_0_port, A4(31) => s_8A_1_neg_31_port
                           , A4(30) => s_8A_1_neg_30_port, A4(29) => 
                           s_8A_1_neg_29_port, A4(28) => s_8A_1_neg_28_port, 
                           A4(27) => s_8A_1_neg_27_port, A4(26) => 
                           s_8A_1_neg_26_port, A4(25) => s_8A_1_neg_25_port, 
                           A4(24) => s_8A_1_neg_24_port, A4(23) => 
                           s_8A_1_neg_23_port, A4(22) => s_8A_1_neg_22_port, 
                           A4(21) => s_8A_1_neg_21_port, A4(20) => 
                           s_8A_1_neg_20_port, A4(19) => s_8A_1_neg_19_port, 
                           A4(18) => s_8A_1_neg_18_port, A4(17) => 
                           s_8A_1_neg_17_port, A4(16) => s_8A_1_neg_16_port, 
                           A4(15) => s_8A_1_neg_15_port, A4(14) => 
                           s_8A_1_neg_14_port, A4(13) => s_8A_1_neg_13_port, 
                           A4(12) => s_8A_1_neg_12_port, A4(11) => 
                           s_8A_1_neg_11_port, A4(10) => s_8A_1_neg_10_port, 
                           A4(9) => s_8A_1_neg_9_port, A4(8) => 
                           s_8A_1_neg_8_port, A4(7) => s_8A_1_neg_7_port, A4(6)
                           => s_8A_1_neg_6_port, A4(5) => s_8A_1_neg_5_port, 
                           A4(4) => s_8A_1_neg_4_port, A4(3) => 
                           s_8A_1_neg_3_port, A4(2) => s_8A_1_neg_2_port, A4(1)
                           => s_8A_1_neg_1_port, A4(0) => s_8A_1_neg_0_port, 
                           SEL(2) => s_sel_1_2_port, SEL(1) => s_sel_1_1_port, 
                           SEL(0) => s_sel_1_0_port, Y(31) => mux2_out_31_port,
                           Y(30) => mux2_out_30_port, Y(29) => mux2_out_29_port
                           , Y(28) => mux2_out_28_port, Y(27) => 
                           mux2_out_27_port, Y(26) => mux2_out_26_port, Y(25) 
                           => mux2_out_25_port, Y(24) => mux2_out_24_port, 
                           Y(23) => mux2_out_23_port, Y(22) => mux2_out_22_port
                           , Y(21) => mux2_out_21_port, Y(20) => 
                           mux2_out_20_port, Y(19) => mux2_out_19_port, Y(18) 
                           => mux2_out_18_port, Y(17) => mux2_out_17_port, 
                           Y(16) => mux2_out_16_port, Y(15) => mux2_out_15_port
                           , Y(14) => mux2_out_14_port, Y(13) => 
                           mux2_out_13_port, Y(12) => mux2_out_12_port, Y(11) 
                           => mux2_out_11_port, Y(10) => mux2_out_10_port, Y(9)
                           => mux2_out_9_port, Y(8) => mux2_out_8_port, Y(7) =>
                           mux2_out_7_port, Y(6) => mux2_out_6_port, Y(5) => 
                           mux2_out_5_port, Y(4) => mux2_out_4_port, Y(3) => 
                           mux2_out_3_port, Y(2) => mux2_out_2_port, Y(1) => 
                           mux2_out_1_port, Y(0) => mux2_out_0_port);
   shift2A_2 : shl1_NBIT32_2 port map( A(31) => A4_reg1_31_port, A(30) => 
                           A4_reg1_30_port, A(29) => A4_reg1_29_port, A(28) => 
                           A4_reg1_28_port, A(27) => A4_reg1_27_port, A(26) => 
                           A4_reg1_26_port, A(25) => A4_reg1_25_port, A(24) => 
                           A4_reg1_24_port, A(23) => A4_reg1_23_port, A(22) => 
                           A4_reg1_22_port, A(21) => A4_reg1_21_port, A(20) => 
                           A4_reg1_20_port, A(19) => A4_reg1_19_port, A(18) => 
                           A4_reg1_18_port, A(17) => A4_reg1_17_port, A(16) => 
                           A4_reg1_16_port, A(15) => A4_reg1_15_port, A(14) => 
                           A4_reg1_14_port, A(13) => A4_reg1_13_port, A(12) => 
                           A4_reg1_12_port, A(11) => A4_reg1_11_port, A(10) => 
                           A4_reg1_10_port, A(9) => A4_reg1_9_port, A(8) => 
                           A4_reg1_8_port, A(7) => A4_reg1_7_port, A(6) => 
                           A4_reg1_6_port, A(5) => A4_reg1_5_port, A(4) => 
                           A4_reg1_4_port, A(3) => A4_reg1_3_port, A(2) => 
                           A4_reg1_2_port, A(1) => A4_reg1_1_port, A(0) => 
                           A4_reg1_0_port, Y(31) => s_A_2_31_port, Y(30) => 
                           s_A_2_30_port, Y(29) => s_A_2_29_port, Y(28) => 
                           s_A_2_28_port, Y(27) => s_A_2_27_port, Y(26) => 
                           s_A_2_26_port, Y(25) => s_A_2_25_port, Y(24) => 
                           s_A_2_24_port, Y(23) => s_A_2_23_port, Y(22) => 
                           s_A_2_22_port, Y(21) => s_A_2_21_port, Y(20) => 
                           s_A_2_20_port, Y(19) => s_A_2_19_port, Y(18) => 
                           s_A_2_18_port, Y(17) => s_A_2_17_port, Y(16) => 
                           s_A_2_16_port, Y(15) => s_A_2_15_port, Y(14) => 
                           s_A_2_14_port, Y(13) => s_A_2_13_port, Y(12) => 
                           s_A_2_12_port, Y(11) => s_A_2_11_port, Y(10) => 
                           s_A_2_10_port, Y(9) => s_A_2_9_port, Y(8) => 
                           s_A_2_8_port, Y(7) => s_A_2_7_port, Y(6) => 
                           s_A_2_6_port, Y(5) => s_A_2_5_port, Y(4) => 
                           s_A_2_4_port, Y(3) => s_A_2_3_port, Y(2) => 
                           s_A_2_2_port, Y(1) => s_A_2_1_port, Y(0) => n_1908);
   shift4A_2 : shl2_NBIT32_2 port map( A(31) => A4_reg1_31_port, A(30) => 
                           A4_reg1_30_port, A(29) => A4_reg1_29_port, A(28) => 
                           A4_reg1_28_port, A(27) => A4_reg1_27_port, A(26) => 
                           A4_reg1_26_port, A(25) => A4_reg1_25_port, A(24) => 
                           A4_reg1_24_port, A(23) => A4_reg1_23_port, A(22) => 
                           A4_reg1_22_port, A(21) => A4_reg1_21_port, A(20) => 
                           A4_reg1_20_port, A(19) => A4_reg1_19_port, A(18) => 
                           A4_reg1_18_port, A(17) => A4_reg1_17_port, A(16) => 
                           A4_reg1_16_port, A(15) => A4_reg1_15_port, A(14) => 
                           A4_reg1_14_port, A(13) => A4_reg1_13_port, A(12) => 
                           A4_reg1_12_port, A(11) => A4_reg1_11_port, A(10) => 
                           A4_reg1_10_port, A(9) => A4_reg1_9_port, A(8) => 
                           A4_reg1_8_port, A(7) => A4_reg1_7_port, A(6) => 
                           A4_reg1_6_port, A(5) => A4_reg1_5_port, A(4) => 
                           A4_reg1_4_port, A(3) => A4_reg1_3_port, A(2) => 
                           A4_reg1_2_port, A(1) => A4_reg1_1_port, A(0) => 
                           A4_reg1_0_port, Y(31) => s_2A_2_31_port, Y(30) => 
                           s_2A_2_30_port, Y(29) => s_2A_2_29_port, Y(28) => 
                           s_2A_2_28_port, Y(27) => s_2A_2_27_port, Y(26) => 
                           s_2A_2_26_port, Y(25) => s_2A_2_25_port, Y(24) => 
                           s_2A_2_24_port, Y(23) => s_2A_2_23_port, Y(22) => 
                           s_2A_2_22_port, Y(21) => s_2A_2_21_port, Y(20) => 
                           s_2A_2_20_port, Y(19) => s_2A_2_19_port, Y(18) => 
                           s_2A_2_18_port, Y(17) => s_2A_2_17_port, Y(16) => 
                           s_2A_2_16_port, Y(15) => s_2A_2_15_port, Y(14) => 
                           s_2A_2_14_port, Y(13) => s_2A_2_13_port, Y(12) => 
                           s_2A_2_12_port, Y(11) => s_2A_2_11_port, Y(10) => 
                           s_2A_2_10_port, Y(9) => s_2A_2_9_port, Y(8) => 
                           s_2A_2_8_port, Y(7) => s_2A_2_7_port, Y(6) => 
                           s_2A_2_6_port, Y(5) => s_2A_2_5_port, Y(4) => 
                           s_2A_2_4_port, Y(3) => s_2A_2_3_port, Y(2) => 
                           s_2A_2_2_port, Y(1) => n_1909, Y(0) => n_1910);
   neg5 : negate_NBIT32_4 port map( A(31) => s_A_2_31_port, A(30) => 
                           s_A_2_30_port, A(29) => s_A_2_29_port, A(28) => 
                           s_A_2_28_port, A(27) => s_A_2_27_port, A(26) => 
                           s_A_2_26_port, A(25) => s_A_2_25_port, A(24) => 
                           s_A_2_24_port, A(23) => s_A_2_23_port, A(22) => 
                           s_A_2_22_port, A(21) => s_A_2_21_port, A(20) => 
                           s_A_2_20_port, A(19) => s_A_2_19_port, A(18) => 
                           s_A_2_18_port, A(17) => s_A_2_17_port, A(16) => 
                           s_A_2_16_port, A(15) => s_A_2_15_port, A(14) => 
                           s_A_2_14_port, A(13) => s_A_2_13_port, A(12) => 
                           s_A_2_12_port, A(11) => s_A_2_11_port, A(10) => 
                           s_A_2_10_port, A(9) => s_A_2_9_port, A(8) => 
                           s_A_2_8_port, A(7) => s_A_2_7_port, A(6) => 
                           s_A_2_6_port, A(5) => s_A_2_5_port, A(4) => 
                           s_A_2_4_port, A(3) => s_A_2_3_port, A(2) => 
                           s_A_2_2_port, A(1) => s_A_2_1_port, A(0) => 
                           s_A_2_0_port, Y(31) => s_A_2_neg_31_port, Y(30) => 
                           s_A_2_neg_30_port, Y(29) => s_A_2_neg_29_port, Y(28)
                           => s_A_2_neg_28_port, Y(27) => s_A_2_neg_27_port, 
                           Y(26) => s_A_2_neg_26_port, Y(25) => 
                           s_A_2_neg_25_port, Y(24) => s_A_2_neg_24_port, Y(23)
                           => s_A_2_neg_23_port, Y(22) => s_A_2_neg_22_port, 
                           Y(21) => s_A_2_neg_21_port, Y(20) => 
                           s_A_2_neg_20_port, Y(19) => s_A_2_neg_19_port, Y(18)
                           => s_A_2_neg_18_port, Y(17) => s_A_2_neg_17_port, 
                           Y(16) => s_A_2_neg_16_port, Y(15) => 
                           s_A_2_neg_15_port, Y(14) => s_A_2_neg_14_port, Y(13)
                           => s_A_2_neg_13_port, Y(12) => s_A_2_neg_12_port, 
                           Y(11) => s_A_2_neg_11_port, Y(10) => 
                           s_A_2_neg_10_port, Y(9) => s_A_2_neg_9_port, Y(8) =>
                           s_A_2_neg_8_port, Y(7) => s_A_2_neg_7_port, Y(6) => 
                           s_A_2_neg_6_port, Y(5) => s_A_2_neg_5_port, Y(4) => 
                           s_A_2_neg_4_port, Y(3) => s_A_2_neg_3_port, Y(2) => 
                           s_A_2_neg_2_port, Y(1) => s_A_2_neg_1_port, Y(0) => 
                           s_A_2_neg_0_port);
   neg6 : negate_NBIT32_3 port map( A(31) => s_2A_2_31_port, A(30) => 
                           s_2A_2_30_port, A(29) => s_2A_2_29_port, A(28) => 
                           s_2A_2_28_port, A(27) => s_2A_2_27_port, A(26) => 
                           s_2A_2_26_port, A(25) => s_2A_2_25_port, A(24) => 
                           s_2A_2_24_port, A(23) => s_2A_2_23_port, A(22) => 
                           s_2A_2_22_port, A(21) => s_2A_2_21_port, A(20) => 
                           s_2A_2_20_port, A(19) => s_2A_2_19_port, A(18) => 
                           s_2A_2_18_port, A(17) => s_2A_2_17_port, A(16) => 
                           s_2A_2_16_port, A(15) => s_2A_2_15_port, A(14) => 
                           s_2A_2_14_port, A(13) => s_2A_2_13_port, A(12) => 
                           s_2A_2_12_port, A(11) => s_2A_2_11_port, A(10) => 
                           s_2A_2_10_port, A(9) => s_2A_2_9_port, A(8) => 
                           s_2A_2_8_port, A(7) => s_2A_2_7_port, A(6) => 
                           s_2A_2_6_port, A(5) => s_2A_2_5_port, A(4) => 
                           s_2A_2_4_port, A(3) => s_2A_2_3_port, A(2) => 
                           s_2A_2_2_port, A(1) => s_2A_2_1_port, A(0) => 
                           s_2A_2_0_port, Y(31) => s_2A_2_neg_31_port, Y(30) =>
                           s_2A_2_neg_30_port, Y(29) => s_2A_2_neg_29_port, 
                           Y(28) => s_2A_2_neg_28_port, Y(27) => 
                           s_2A_2_neg_27_port, Y(26) => s_2A_2_neg_26_port, 
                           Y(25) => s_2A_2_neg_25_port, Y(24) => 
                           s_2A_2_neg_24_port, Y(23) => s_2A_2_neg_23_port, 
                           Y(22) => s_2A_2_neg_22_port, Y(21) => 
                           s_2A_2_neg_21_port, Y(20) => s_2A_2_neg_20_port, 
                           Y(19) => s_2A_2_neg_19_port, Y(18) => 
                           s_2A_2_neg_18_port, Y(17) => s_2A_2_neg_17_port, 
                           Y(16) => s_2A_2_neg_16_port, Y(15) => 
                           s_2A_2_neg_15_port, Y(14) => s_2A_2_neg_14_port, 
                           Y(13) => s_2A_2_neg_13_port, Y(12) => 
                           s_2A_2_neg_12_port, Y(11) => s_2A_2_neg_11_port, 
                           Y(10) => s_2A_2_neg_10_port, Y(9) => 
                           s_2A_2_neg_9_port, Y(8) => s_2A_2_neg_8_port, Y(7) 
                           => s_2A_2_neg_7_port, Y(6) => s_2A_2_neg_6_port, 
                           Y(5) => s_2A_2_neg_5_port, Y(4) => s_2A_2_neg_4_port
                           , Y(3) => s_2A_2_neg_3_port, Y(2) => 
                           s_2A_2_neg_2_port, Y(1) => s_2A_2_neg_1_port, Y(0) 
                           => s_2A_2_neg_0_port);
   mux3 : mux51_gen_NBIT32_2 port map( A0(31) => X_Logic0_port, A0(30) => 
                           X_Logic0_port, A0(29) => X_Logic0_port, A0(28) => 
                           X_Logic0_port, A0(27) => X_Logic0_port, A0(26) => 
                           X_Logic0_port, A0(25) => X_Logic0_port, A0(24) => 
                           X_Logic0_port, A0(23) => X_Logic0_port, A0(22) => 
                           X_Logic0_port, A0(21) => X_Logic0_port, A0(20) => 
                           X_Logic0_port, A0(19) => X_Logic0_port, A0(18) => 
                           X_Logic0_port, A0(17) => X_Logic0_port, A0(16) => 
                           X_Logic0_port, A0(15) => X_Logic0_port, A0(14) => 
                           X_Logic0_port, A0(13) => X_Logic0_port, A0(12) => 
                           X_Logic0_port, A0(11) => X_Logic0_port, A0(10) => 
                           X_Logic0_port, A0(9) => X_Logic0_port, A0(8) => 
                           X_Logic0_port, A0(7) => X_Logic0_port, A0(6) => 
                           X_Logic0_port, A0(5) => X_Logic0_port, A0(4) => 
                           X_Logic0_port, A0(3) => X_Logic0_port, A0(2) => 
                           X_Logic0_port, A0(1) => X_Logic0_port, A0(0) => 
                           X_Logic0_port, A1(31) => s_A_2_31_port, A1(30) => 
                           s_A_2_30_port, A1(29) => s_A_2_29_port, A1(28) => 
                           s_A_2_28_port, A1(27) => s_A_2_27_port, A1(26) => 
                           s_A_2_26_port, A1(25) => s_A_2_25_port, A1(24) => 
                           s_A_2_24_port, A1(23) => s_A_2_23_port, A1(22) => 
                           s_A_2_22_port, A1(21) => s_A_2_21_port, A1(20) => 
                           s_A_2_20_port, A1(19) => s_A_2_19_port, A1(18) => 
                           s_A_2_18_port, A1(17) => s_A_2_17_port, A1(16) => 
                           s_A_2_16_port, A1(15) => s_A_2_15_port, A1(14) => 
                           s_A_2_14_port, A1(13) => s_A_2_13_port, A1(12) => 
                           s_A_2_12_port, A1(11) => s_A_2_11_port, A1(10) => 
                           s_A_2_10_port, A1(9) => s_A_2_9_port, A1(8) => 
                           s_A_2_8_port, A1(7) => s_A_2_7_port, A1(6) => 
                           s_A_2_6_port, A1(5) => s_A_2_5_port, A1(4) => 
                           s_A_2_4_port, A1(3) => s_A_2_3_port, A1(2) => 
                           s_A_2_2_port, A1(1) => s_A_2_1_port, A1(0) => 
                           s_A_2_0_port, A2(31) => s_A_2_neg_31_port, A2(30) =>
                           s_A_2_neg_30_port, A2(29) => s_A_2_neg_29_port, 
                           A2(28) => s_A_2_neg_28_port, A2(27) => 
                           s_A_2_neg_27_port, A2(26) => s_A_2_neg_26_port, 
                           A2(25) => s_A_2_neg_25_port, A2(24) => 
                           s_A_2_neg_24_port, A2(23) => s_A_2_neg_23_port, 
                           A2(22) => s_A_2_neg_22_port, A2(21) => 
                           s_A_2_neg_21_port, A2(20) => s_A_2_neg_20_port, 
                           A2(19) => s_A_2_neg_19_port, A2(18) => 
                           s_A_2_neg_18_port, A2(17) => s_A_2_neg_17_port, 
                           A2(16) => s_A_2_neg_16_port, A2(15) => 
                           s_A_2_neg_15_port, A2(14) => s_A_2_neg_14_port, 
                           A2(13) => s_A_2_neg_13_port, A2(12) => 
                           s_A_2_neg_12_port, A2(11) => s_A_2_neg_11_port, 
                           A2(10) => s_A_2_neg_10_port, A2(9) => 
                           s_A_2_neg_9_port, A2(8) => s_A_2_neg_8_port, A2(7) 
                           => s_A_2_neg_7_port, A2(6) => s_A_2_neg_6_port, 
                           A2(5) => s_A_2_neg_5_port, A2(4) => s_A_2_neg_4_port
                           , A2(3) => s_A_2_neg_3_port, A2(2) => 
                           s_A_2_neg_2_port, A2(1) => s_A_2_neg_1_port, A2(0) 
                           => s_A_2_neg_0_port, A3(31) => s_2A_2_31_port, 
                           A3(30) => s_2A_2_30_port, A3(29) => s_2A_2_29_port, 
                           A3(28) => s_2A_2_28_port, A3(27) => s_2A_2_27_port, 
                           A3(26) => s_2A_2_26_port, A3(25) => s_2A_2_25_port, 
                           A3(24) => s_2A_2_24_port, A3(23) => s_2A_2_23_port, 
                           A3(22) => s_2A_2_22_port, A3(21) => s_2A_2_21_port, 
                           A3(20) => s_2A_2_20_port, A3(19) => s_2A_2_19_port, 
                           A3(18) => s_2A_2_18_port, A3(17) => s_2A_2_17_port, 
                           A3(16) => s_2A_2_16_port, A3(15) => s_2A_2_15_port, 
                           A3(14) => s_2A_2_14_port, A3(13) => s_2A_2_13_port, 
                           A3(12) => s_2A_2_12_port, A3(11) => s_2A_2_11_port, 
                           A3(10) => s_2A_2_10_port, A3(9) => s_2A_2_9_port, 
                           A3(8) => s_2A_2_8_port, A3(7) => s_2A_2_7_port, 
                           A3(6) => s_2A_2_6_port, A3(5) => s_2A_2_5_port, 
                           A3(4) => s_2A_2_4_port, A3(3) => s_2A_2_3_port, 
                           A3(2) => s_2A_2_2_port, A3(1) => s_2A_2_1_port, 
                           A3(0) => s_2A_2_0_port, A4(31) => s_2A_2_neg_31_port
                           , A4(30) => s_2A_2_neg_30_port, A4(29) => 
                           s_2A_2_neg_29_port, A4(28) => s_2A_2_neg_28_port, 
                           A4(27) => s_2A_2_neg_27_port, A4(26) => 
                           s_2A_2_neg_26_port, A4(25) => s_2A_2_neg_25_port, 
                           A4(24) => s_2A_2_neg_24_port, A4(23) => 
                           s_2A_2_neg_23_port, A4(22) => s_2A_2_neg_22_port, 
                           A4(21) => s_2A_2_neg_21_port, A4(20) => 
                           s_2A_2_neg_20_port, A4(19) => s_2A_2_neg_19_port, 
                           A4(18) => s_2A_2_neg_18_port, A4(17) => 
                           s_2A_2_neg_17_port, A4(16) => s_2A_2_neg_16_port, 
                           A4(15) => s_2A_2_neg_15_port, A4(14) => 
                           s_2A_2_neg_14_port, A4(13) => s_2A_2_neg_13_port, 
                           A4(12) => s_2A_2_neg_12_port, A4(11) => 
                           s_2A_2_neg_11_port, A4(10) => s_2A_2_neg_10_port, 
                           A4(9) => s_2A_2_neg_9_port, A4(8) => 
                           s_2A_2_neg_8_port, A4(7) => s_2A_2_neg_7_port, A4(6)
                           => s_2A_2_neg_6_port, A4(5) => s_2A_2_neg_5_port, 
                           A4(4) => s_2A_2_neg_4_port, A4(3) => 
                           s_2A_2_neg_3_port, A4(2) => s_2A_2_neg_2_port, A4(1)
                           => s_2A_2_neg_1_port, A4(0) => s_2A_2_neg_0_port, 
                           SEL(2) => enc_reg21_2_port, SEL(1) => 
                           enc_reg21_1_port, SEL(0) => enc_reg21_0_port, Y(31) 
                           => mux_2_out_31_port, Y(30) => mux_2_out_30_port, 
                           Y(29) => mux_2_out_29_port, Y(28) => 
                           mux_2_out_28_port, Y(27) => mux_2_out_27_port, Y(26)
                           => mux_2_out_26_port, Y(25) => mux_2_out_25_port, 
                           Y(24) => mux_2_out_24_port, Y(23) => 
                           mux_2_out_23_port, Y(22) => mux_2_out_22_port, Y(21)
                           => mux_2_out_21_port, Y(20) => mux_2_out_20_port, 
                           Y(19) => mux_2_out_19_port, Y(18) => 
                           mux_2_out_18_port, Y(17) => mux_2_out_17_port, Y(16)
                           => mux_2_out_16_port, Y(15) => mux_2_out_15_port, 
                           Y(14) => mux_2_out_14_port, Y(13) => 
                           mux_2_out_13_port, Y(12) => mux_2_out_12_port, Y(11)
                           => mux_2_out_11_port, Y(10) => mux_2_out_10_port, 
                           Y(9) => mux_2_out_9_port, Y(8) => mux_2_out_8_port, 
                           Y(7) => mux_2_out_7_port, Y(6) => mux_2_out_6_port, 
                           Y(5) => mux_2_out_5_port, Y(4) => mux_2_out_4_port, 
                           Y(3) => mux_2_out_3_port, Y(2) => mux_2_out_2_port, 
                           Y(1) => mux_2_out_1_port, Y(0) => mux_2_out_0_port);
   SUM1 : P4_ADDER_NBIT64_0 port map( A(63) => n12, A(62) => n12, A(61) => n12,
                           A(60) => n12, A(59) => n12, A(58) => n13, A(57) => 
                           n13, A(56) => n13, A(55) => n13, A(54) => n13, A(53)
                           => n13, A(52) => n14, A(51) => n14, A(50) => n14, 
                           A(49) => n14, A(48) => n14, A(47) => n14, A(46) => 
                           n15, A(45) => n15, A(44) => n15, A(43) => n15, A(42)
                           => n15, A(41) => n15, A(40) => n16, A(39) => n16, 
                           A(38) => n16, A(37) => n16, A(36) => n16, A(35) => 
                           n16, A(34) => n17, A(33) => n17, A(32) => n17, A(31)
                           => n17, A(30) => mux1_reg1_30_port, A(29) => 
                           mux1_reg1_29_port, A(28) => mux1_reg1_28_port, A(27)
                           => mux1_reg1_27_port, A(26) => mux1_reg1_26_port, 
                           A(25) => mux1_reg1_25_port, A(24) => 
                           mux1_reg1_24_port, A(23) => mux1_reg1_23_port, A(22)
                           => mux1_reg1_22_port, A(21) => mux1_reg1_21_port, 
                           A(20) => mux1_reg1_20_port, A(19) => 
                           mux1_reg1_19_port, A(18) => mux1_reg1_18_port, A(17)
                           => mux1_reg1_17_port, A(16) => mux1_reg1_16_port, 
                           A(15) => mux1_reg1_15_port, A(14) => 
                           mux1_reg1_14_port, A(13) => mux1_reg1_13_port, A(12)
                           => mux1_reg1_12_port, A(11) => mux1_reg1_11_port, 
                           A(10) => mux1_reg1_10_port, A(9) => mux1_reg1_9_port
                           , A(8) => mux1_reg1_8_port, A(7) => mux1_reg1_7_port
                           , A(6) => mux1_reg1_6_port, A(5) => mux1_reg1_5_port
                           , A(4) => mux1_reg1_4_port, A(3) => mux1_reg1_3_port
                           , A(2) => mux1_reg1_2_port, A(1) => mux1_reg1_1_port
                           , A(0) => mux1_reg1_0_port, B(63) => n9, B(62) => n9
                           , B(61) => n9, B(60) => n9, B(59) => n9, B(58) => n9
                           , B(57) => n9, B(56) => n9, B(55) => n9, B(54) => n9
                           , B(53) => n9, B(52) => n8, B(51) => n8, B(50) => n8
                           , B(49) => n8, B(48) => n8, B(47) => n8, B(46) => n8
                           , B(45) => n8, B(44) => n8, B(43) => n8, B(42) => n8
                           , B(41) => n7, B(40) => n7, B(39) => n7, B(38) => n7
                           , B(37) => n7, B(36) => n7, B(35) => n7, B(34) => n7
                           , B(33) => n7, B(32) => n7, B(31) => n7, B(30) => 
                           mux2_reg1_30_port, B(29) => mux2_reg1_29_port, B(28)
                           => mux2_reg1_28_port, B(27) => mux2_reg1_27_port, 
                           B(26) => mux2_reg1_26_port, B(25) => 
                           mux2_reg1_25_port, B(24) => mux2_reg1_24_port, B(23)
                           => mux2_reg1_23_port, B(22) => mux2_reg1_22_port, 
                           B(21) => mux2_reg1_21_port, B(20) => 
                           mux2_reg1_20_port, B(19) => mux2_reg1_19_port, B(18)
                           => mux2_reg1_18_port, B(17) => mux2_reg1_17_port, 
                           B(16) => mux2_reg1_16_port, B(15) => 
                           mux2_reg1_15_port, B(14) => mux2_reg1_14_port, B(13)
                           => mux2_reg1_13_port, B(12) => mux2_reg1_12_port, 
                           B(11) => mux2_reg1_11_port, B(10) => 
                           mux2_reg1_10_port, B(9) => mux2_reg1_9_port, B(8) =>
                           mux2_reg1_8_port, B(7) => mux2_reg1_7_port, B(6) => 
                           mux2_reg1_6_port, B(5) => mux2_reg1_5_port, B(4) => 
                           mux2_reg1_4_port, B(3) => mux2_reg1_3_port, B(2) => 
                           mux2_reg1_2_port, B(1) => mux2_reg1_1_port, B(0) => 
                           mux2_reg1_0_port, Cin => X_Logic0_port, S(63) => 
                           sum_2_out_63_port, S(62) => sum_2_out_62_port, S(61)
                           => sum_2_out_61_port, S(60) => sum_2_out_60_port, 
                           S(59) => sum_2_out_59_port, S(58) => 
                           sum_2_out_58_port, S(57) => sum_2_out_57_port, S(56)
                           => sum_2_out_56_port, S(55) => sum_2_out_55_port, 
                           S(54) => sum_2_out_54_port, S(53) => 
                           sum_2_out_53_port, S(52) => sum_2_out_52_port, S(51)
                           => sum_2_out_51_port, S(50) => sum_2_out_50_port, 
                           S(49) => sum_2_out_49_port, S(48) => 
                           sum_2_out_48_port, S(47) => sum_2_out_47_port, S(46)
                           => sum_2_out_46_port, S(45) => sum_2_out_45_port, 
                           S(44) => sum_2_out_44_port, S(43) => 
                           sum_2_out_43_port, S(42) => sum_2_out_42_port, S(41)
                           => sum_2_out_41_port, S(40) => sum_2_out_40_port, 
                           S(39) => sum_2_out_39_port, S(38) => 
                           sum_2_out_38_port, S(37) => sum_2_out_37_port, S(36)
                           => sum_2_out_36_port, S(35) => sum_2_out_35_port, 
                           S(34) => sum_2_out_34_port, S(33) => 
                           sum_2_out_33_port, S(32) => sum_2_out_32_port, S(31)
                           => sum_2_out_31_port, S(30) => sum_2_out_30_port, 
                           S(29) => sum_2_out_29_port, S(28) => 
                           sum_2_out_28_port, S(27) => sum_2_out_27_port, S(26)
                           => sum_2_out_26_port, S(25) => sum_2_out_25_port, 
                           S(24) => sum_2_out_24_port, S(23) => 
                           sum_2_out_23_port, S(22) => sum_2_out_22_port, S(21)
                           => sum_2_out_21_port, S(20) => sum_2_out_20_port, 
                           S(19) => sum_2_out_19_port, S(18) => 
                           sum_2_out_18_port, S(17) => sum_2_out_17_port, S(16)
                           => sum_2_out_16_port, S(15) => sum_2_out_15_port, 
                           S(14) => sum_2_out_14_port, S(13) => 
                           sum_2_out_13_port, S(12) => sum_2_out_12_port, S(11)
                           => sum_2_out_11_port, S(10) => sum_2_out_10_port, 
                           S(9) => sum_2_out_9_port, S(8) => sum_2_out_8_port, 
                           S(7) => sum_2_out_7_port, S(6) => sum_2_out_6_port, 
                           S(5) => sum_2_out_5_port, S(4) => sum_2_out_4_port, 
                           S(3) => sum_2_out_3_port, S(2) => sum_2_out_2_port, 
                           S(1) => sum_2_out_1_port, S(0) => sum_2_out_0_port, 
                           Cout => n_1911, ovf => n_1912);
   shift2A_3 : shl1_NBIT32_1 port map( A(31) => A4_reg2_31_port, A(30) => 
                           A4_reg2_30_port, A(29) => A4_reg2_29_port, A(28) => 
                           A4_reg2_28_port, A(27) => A4_reg2_27_port, A(26) => 
                           A4_reg2_26_port, A(25) => A4_reg2_25_port, A(24) => 
                           A4_reg2_24_port, A(23) => A4_reg2_23_port, A(22) => 
                           A4_reg2_22_port, A(21) => A4_reg2_21_port, A(20) => 
                           A4_reg2_20_port, A(19) => A4_reg2_19_port, A(18) => 
                           A4_reg2_18_port, A(17) => A4_reg2_17_port, A(16) => 
                           A4_reg2_16_port, A(15) => A4_reg2_15_port, A(14) => 
                           A4_reg2_14_port, A(13) => A4_reg2_13_port, A(12) => 
                           A4_reg2_12_port, A(11) => A4_reg2_11_port, A(10) => 
                           A4_reg2_10_port, A(9) => A4_reg2_9_port, A(8) => 
                           A4_reg2_8_port, A(7) => A4_reg2_7_port, A(6) => 
                           A4_reg2_6_port, A(5) => A4_reg2_5_port, A(4) => 
                           A4_reg2_4_port, A(3) => A4_reg2_3_port, A(2) => 
                           A4_reg2_2_port, A(1) => A4_reg2_1_port, A(0) => 
                           A4_reg2_0_port, Y(31) => s_A_3_31_port, Y(30) => 
                           s_A_3_30_port, Y(29) => s_A_3_29_port, Y(28) => 
                           s_A_3_28_port, Y(27) => s_A_3_27_port, Y(26) => 
                           s_A_3_26_port, Y(25) => s_A_3_25_port, Y(24) => 
                           s_A_3_24_port, Y(23) => s_A_3_23_port, Y(22) => 
                           s_A_3_22_port, Y(21) => s_A_3_21_port, Y(20) => 
                           s_A_3_20_port, Y(19) => s_A_3_19_port, Y(18) => 
                           s_A_3_18_port, Y(17) => s_A_3_17_port, Y(16) => 
                           s_A_3_16_port, Y(15) => s_A_3_15_port, Y(14) => 
                           s_A_3_14_port, Y(13) => s_A_3_13_port, Y(12) => 
                           s_A_3_12_port, Y(11) => s_A_3_11_port, Y(10) => 
                           s_A_3_10_port, Y(9) => s_A_3_9_port, Y(8) => 
                           s_A_3_8_port, Y(7) => s_A_3_7_port, Y(6) => 
                           s_A_3_6_port, Y(5) => s_A_3_5_port, Y(4) => 
                           s_A_3_4_port, Y(3) => s_A_3_3_port, Y(2) => 
                           s_A_3_2_port, Y(1) => s_A_3_1_port, Y(0) => n_1913);
   shift4A_3 : shl2_NBIT32_1 port map( A(31) => A4_reg2_31_port, A(30) => 
                           A4_reg2_30_port, A(29) => A4_reg2_29_port, A(28) => 
                           A4_reg2_28_port, A(27) => A4_reg2_27_port, A(26) => 
                           A4_reg2_26_port, A(25) => A4_reg2_25_port, A(24) => 
                           A4_reg2_24_port, A(23) => A4_reg2_23_port, A(22) => 
                           A4_reg2_22_port, A(21) => A4_reg2_21_port, A(20) => 
                           A4_reg2_20_port, A(19) => A4_reg2_19_port, A(18) => 
                           A4_reg2_18_port, A(17) => A4_reg2_17_port, A(16) => 
                           A4_reg2_16_port, A(15) => A4_reg2_15_port, A(14) => 
                           A4_reg2_14_port, A(13) => A4_reg2_13_port, A(12) => 
                           A4_reg2_12_port, A(11) => A4_reg2_11_port, A(10) => 
                           A4_reg2_10_port, A(9) => A4_reg2_9_port, A(8) => 
                           A4_reg2_8_port, A(7) => A4_reg2_7_port, A(6) => 
                           A4_reg2_6_port, A(5) => A4_reg2_5_port, A(4) => 
                           A4_reg2_4_port, A(3) => A4_reg2_3_port, A(2) => 
                           A4_reg2_2_port, A(1) => A4_reg2_1_port, A(0) => 
                           A4_reg2_0_port, Y(31) => s_2A_3_31_port, Y(30) => 
                           s_2A_3_30_port, Y(29) => s_2A_3_29_port, Y(28) => 
                           s_2A_3_28_port, Y(27) => s_2A_3_27_port, Y(26) => 
                           s_2A_3_26_port, Y(25) => s_2A_3_25_port, Y(24) => 
                           s_2A_3_24_port, Y(23) => s_2A_3_23_port, Y(22) => 
                           s_2A_3_22_port, Y(21) => s_2A_3_21_port, Y(20) => 
                           s_2A_3_20_port, Y(19) => s_2A_3_19_port, Y(18) => 
                           s_2A_3_18_port, Y(17) => s_2A_3_17_port, Y(16) => 
                           s_2A_3_16_port, Y(15) => s_2A_3_15_port, Y(14) => 
                           s_2A_3_14_port, Y(13) => s_2A_3_13_port, Y(12) => 
                           s_2A_3_12_port, Y(11) => s_2A_3_11_port, Y(10) => 
                           s_2A_3_10_port, Y(9) => s_2A_3_9_port, Y(8) => 
                           s_2A_3_8_port, Y(7) => s_2A_3_7_port, Y(6) => 
                           s_2A_3_6_port, Y(5) => s_2A_3_5_port, Y(4) => 
                           s_2A_3_4_port, Y(3) => s_2A_3_3_port, Y(2) => 
                           s_2A_3_2_port, Y(1) => n_1914, Y(0) => n_1915);
   neg7 : negate_NBIT32_2 port map( A(31) => s_A_3_31_port, A(30) => 
                           s_A_3_30_port, A(29) => s_A_3_29_port, A(28) => 
                           s_A_3_28_port, A(27) => s_A_3_27_port, A(26) => 
                           s_A_3_26_port, A(25) => s_A_3_25_port, A(24) => 
                           s_A_3_24_port, A(23) => s_A_3_23_port, A(22) => 
                           s_A_3_22_port, A(21) => s_A_3_21_port, A(20) => 
                           s_A_3_20_port, A(19) => s_A_3_19_port, A(18) => 
                           s_A_3_18_port, A(17) => s_A_3_17_port, A(16) => 
                           s_A_3_16_port, A(15) => s_A_3_15_port, A(14) => 
                           s_A_3_14_port, A(13) => s_A_3_13_port, A(12) => 
                           s_A_3_12_port, A(11) => s_A_3_11_port, A(10) => 
                           s_A_3_10_port, A(9) => s_A_3_9_port, A(8) => 
                           s_A_3_8_port, A(7) => s_A_3_7_port, A(6) => 
                           s_A_3_6_port, A(5) => s_A_3_5_port, A(4) => 
                           s_A_3_4_port, A(3) => s_A_3_3_port, A(2) => 
                           s_A_3_2_port, A(1) => s_A_3_1_port, A(0) => 
                           s_A_3_0_port, Y(31) => s_A_3_neg_31_port, Y(30) => 
                           s_A_3_neg_30_port, Y(29) => s_A_3_neg_29_port, Y(28)
                           => s_A_3_neg_28_port, Y(27) => s_A_3_neg_27_port, 
                           Y(26) => s_A_3_neg_26_port, Y(25) => 
                           s_A_3_neg_25_port, Y(24) => s_A_3_neg_24_port, Y(23)
                           => s_A_3_neg_23_port, Y(22) => s_A_3_neg_22_port, 
                           Y(21) => s_A_3_neg_21_port, Y(20) => 
                           s_A_3_neg_20_port, Y(19) => s_A_3_neg_19_port, Y(18)
                           => s_A_3_neg_18_port, Y(17) => s_A_3_neg_17_port, 
                           Y(16) => s_A_3_neg_16_port, Y(15) => 
                           s_A_3_neg_15_port, Y(14) => s_A_3_neg_14_port, Y(13)
                           => s_A_3_neg_13_port, Y(12) => s_A_3_neg_12_port, 
                           Y(11) => s_A_3_neg_11_port, Y(10) => 
                           s_A_3_neg_10_port, Y(9) => s_A_3_neg_9_port, Y(8) =>
                           s_A_3_neg_8_port, Y(7) => s_A_3_neg_7_port, Y(6) => 
                           s_A_3_neg_6_port, Y(5) => s_A_3_neg_5_port, Y(4) => 
                           s_A_3_neg_4_port, Y(3) => s_A_3_neg_3_port, Y(2) => 
                           s_A_3_neg_2_port, Y(1) => s_A_3_neg_1_port, Y(0) => 
                           s_A_3_neg_0_port);
   neg8 : negate_NBIT32_1 port map( A(31) => s_2A_3_31_port, A(30) => 
                           s_2A_3_30_port, A(29) => s_2A_3_29_port, A(28) => 
                           s_2A_3_28_port, A(27) => s_2A_3_27_port, A(26) => 
                           s_2A_3_26_port, A(25) => s_2A_3_25_port, A(24) => 
                           s_2A_3_24_port, A(23) => s_2A_3_23_port, A(22) => 
                           s_2A_3_22_port, A(21) => s_2A_3_21_port, A(20) => 
                           s_2A_3_20_port, A(19) => s_2A_3_19_port, A(18) => 
                           s_2A_3_18_port, A(17) => s_2A_3_17_port, A(16) => 
                           s_2A_3_16_port, A(15) => s_2A_3_15_port, A(14) => 
                           s_2A_3_14_port, A(13) => s_2A_3_13_port, A(12) => 
                           s_2A_3_12_port, A(11) => s_2A_3_11_port, A(10) => 
                           s_2A_3_10_port, A(9) => s_2A_3_9_port, A(8) => 
                           s_2A_3_8_port, A(7) => s_2A_3_7_port, A(6) => 
                           s_2A_3_6_port, A(5) => s_2A_3_5_port, A(4) => 
                           s_2A_3_4_port, A(3) => s_2A_3_3_port, A(2) => 
                           s_2A_3_2_port, A(1) => s_2A_3_1_port, A(0) => 
                           s_2A_3_0_port, Y(31) => s_2A_3_neg_31_port, Y(30) =>
                           s_2A_3_neg_30_port, Y(29) => s_2A_3_neg_29_port, 
                           Y(28) => s_2A_3_neg_28_port, Y(27) => 
                           s_2A_3_neg_27_port, Y(26) => s_2A_3_neg_26_port, 
                           Y(25) => s_2A_3_neg_25_port, Y(24) => 
                           s_2A_3_neg_24_port, Y(23) => s_2A_3_neg_23_port, 
                           Y(22) => s_2A_3_neg_22_port, Y(21) => 
                           s_2A_3_neg_21_port, Y(20) => s_2A_3_neg_20_port, 
                           Y(19) => s_2A_3_neg_19_port, Y(18) => 
                           s_2A_3_neg_18_port, Y(17) => s_2A_3_neg_17_port, 
                           Y(16) => s_2A_3_neg_16_port, Y(15) => 
                           s_2A_3_neg_15_port, Y(14) => s_2A_3_neg_14_port, 
                           Y(13) => s_2A_3_neg_13_port, Y(12) => 
                           s_2A_3_neg_12_port, Y(11) => s_2A_3_neg_11_port, 
                           Y(10) => s_2A_3_neg_10_port, Y(9) => 
                           s_2A_3_neg_9_port, Y(8) => s_2A_3_neg_8_port, Y(7) 
                           => s_2A_3_neg_7_port, Y(6) => s_2A_3_neg_6_port, 
                           Y(5) => s_2A_3_neg_5_port, Y(4) => s_2A_3_neg_4_port
                           , Y(3) => s_2A_3_neg_3_port, Y(2) => 
                           s_2A_3_neg_2_port, Y(1) => s_2A_3_neg_1_port, Y(0) 
                           => s_2A_3_neg_0_port);
   mux4 : mux51_gen_NBIT32_1 port map( A0(31) => X_Logic0_port, A0(30) => 
                           X_Logic0_port, A0(29) => X_Logic0_port, A0(28) => 
                           X_Logic0_port, A0(27) => X_Logic0_port, A0(26) => 
                           X_Logic0_port, A0(25) => X_Logic0_port, A0(24) => 
                           X_Logic0_port, A0(23) => X_Logic0_port, A0(22) => 
                           X_Logic0_port, A0(21) => X_Logic0_port, A0(20) => 
                           X_Logic0_port, A0(19) => X_Logic0_port, A0(18) => 
                           X_Logic0_port, A0(17) => X_Logic0_port, A0(16) => 
                           X_Logic0_port, A0(15) => X_Logic0_port, A0(14) => 
                           X_Logic0_port, A0(13) => X_Logic0_port, A0(12) => 
                           X_Logic0_port, A0(11) => X_Logic0_port, A0(10) => 
                           X_Logic0_port, A0(9) => X_Logic0_port, A0(8) => 
                           X_Logic0_port, A0(7) => X_Logic0_port, A0(6) => 
                           X_Logic0_port, A0(5) => X_Logic0_port, A0(4) => 
                           X_Logic0_port, A0(3) => X_Logic0_port, A0(2) => 
                           X_Logic0_port, A0(1) => X_Logic0_port, A0(0) => 
                           X_Logic0_port, A1(31) => s_A_3_31_port, A1(30) => 
                           s_A_3_30_port, A1(29) => s_A_3_29_port, A1(28) => 
                           s_A_3_28_port, A1(27) => s_A_3_27_port, A1(26) => 
                           s_A_3_26_port, A1(25) => s_A_3_25_port, A1(24) => 
                           s_A_3_24_port, A1(23) => s_A_3_23_port, A1(22) => 
                           s_A_3_22_port, A1(21) => s_A_3_21_port, A1(20) => 
                           s_A_3_20_port, A1(19) => s_A_3_19_port, A1(18) => 
                           s_A_3_18_port, A1(17) => s_A_3_17_port, A1(16) => 
                           s_A_3_16_port, A1(15) => s_A_3_15_port, A1(14) => 
                           s_A_3_14_port, A1(13) => s_A_3_13_port, A1(12) => 
                           s_A_3_12_port, A1(11) => s_A_3_11_port, A1(10) => 
                           s_A_3_10_port, A1(9) => s_A_3_9_port, A1(8) => 
                           s_A_3_8_port, A1(7) => s_A_3_7_port, A1(6) => 
                           s_A_3_6_port, A1(5) => s_A_3_5_port, A1(4) => 
                           s_A_3_4_port, A1(3) => s_A_3_3_port, A1(2) => 
                           s_A_3_2_port, A1(1) => s_A_3_1_port, A1(0) => 
                           s_A_3_0_port, A2(31) => s_A_3_neg_31_port, A2(30) =>
                           s_A_3_neg_30_port, A2(29) => s_A_3_neg_29_port, 
                           A2(28) => s_A_3_neg_28_port, A2(27) => 
                           s_A_3_neg_27_port, A2(26) => s_A_3_neg_26_port, 
                           A2(25) => s_A_3_neg_25_port, A2(24) => 
                           s_A_3_neg_24_port, A2(23) => s_A_3_neg_23_port, 
                           A2(22) => s_A_3_neg_22_port, A2(21) => 
                           s_A_3_neg_21_port, A2(20) => s_A_3_neg_20_port, 
                           A2(19) => s_A_3_neg_19_port, A2(18) => 
                           s_A_3_neg_18_port, A2(17) => s_A_3_neg_17_port, 
                           A2(16) => s_A_3_neg_16_port, A2(15) => 
                           s_A_3_neg_15_port, A2(14) => s_A_3_neg_14_port, 
                           A2(13) => s_A_3_neg_13_port, A2(12) => 
                           s_A_3_neg_12_port, A2(11) => s_A_3_neg_11_port, 
                           A2(10) => s_A_3_neg_10_port, A2(9) => 
                           s_A_3_neg_9_port, A2(8) => s_A_3_neg_8_port, A2(7) 
                           => s_A_3_neg_7_port, A2(6) => s_A_3_neg_6_port, 
                           A2(5) => s_A_3_neg_5_port, A2(4) => s_A_3_neg_4_port
                           , A2(3) => s_A_3_neg_3_port, A2(2) => 
                           s_A_3_neg_2_port, A2(1) => s_A_3_neg_1_port, A2(0) 
                           => s_A_3_neg_0_port, A3(31) => s_2A_3_31_port, 
                           A3(30) => s_2A_3_30_port, A3(29) => s_2A_3_29_port, 
                           A3(28) => s_2A_3_28_port, A3(27) => s_2A_3_27_port, 
                           A3(26) => s_2A_3_26_port, A3(25) => s_2A_3_25_port, 
                           A3(24) => s_2A_3_24_port, A3(23) => s_2A_3_23_port, 
                           A3(22) => s_2A_3_22_port, A3(21) => s_2A_3_21_port, 
                           A3(20) => s_2A_3_20_port, A3(19) => s_2A_3_19_port, 
                           A3(18) => s_2A_3_18_port, A3(17) => s_2A_3_17_port, 
                           A3(16) => s_2A_3_16_port, A3(15) => s_2A_3_15_port, 
                           A3(14) => s_2A_3_14_port, A3(13) => s_2A_3_13_port, 
                           A3(12) => s_2A_3_12_port, A3(11) => s_2A_3_11_port, 
                           A3(10) => s_2A_3_10_port, A3(9) => s_2A_3_9_port, 
                           A3(8) => s_2A_3_8_port, A3(7) => s_2A_3_7_port, 
                           A3(6) => s_2A_3_6_port, A3(5) => s_2A_3_5_port, 
                           A3(4) => s_2A_3_4_port, A3(3) => s_2A_3_3_port, 
                           A3(2) => s_2A_3_2_port, A3(1) => s_2A_3_1_port, 
                           A3(0) => s_2A_3_0_port, A4(31) => s_2A_3_neg_31_port
                           , A4(30) => s_2A_3_neg_30_port, A4(29) => 
                           s_2A_3_neg_29_port, A4(28) => s_2A_3_neg_28_port, 
                           A4(27) => s_2A_3_neg_27_port, A4(26) => 
                           s_2A_3_neg_26_port, A4(25) => s_2A_3_neg_25_port, 
                           A4(24) => s_2A_3_neg_24_port, A4(23) => 
                           s_2A_3_neg_23_port, A4(22) => s_2A_3_neg_22_port, 
                           A4(21) => s_2A_3_neg_21_port, A4(20) => 
                           s_2A_3_neg_20_port, A4(19) => s_2A_3_neg_19_port, 
                           A4(18) => s_2A_3_neg_18_port, A4(17) => 
                           s_2A_3_neg_17_port, A4(16) => s_2A_3_neg_16_port, 
                           A4(15) => s_2A_3_neg_15_port, A4(14) => 
                           s_2A_3_neg_14_port, A4(13) => s_2A_3_neg_13_port, 
                           A4(12) => s_2A_3_neg_12_port, A4(11) => 
                           s_2A_3_neg_11_port, A4(10) => s_2A_3_neg_10_port, 
                           A4(9) => s_2A_3_neg_9_port, A4(8) => 
                           s_2A_3_neg_8_port, A4(7) => s_2A_3_neg_7_port, A4(6)
                           => s_2A_3_neg_6_port, A4(5) => s_2A_3_neg_5_port, 
                           A4(4) => s_2A_3_neg_4_port, A4(3) => 
                           s_2A_3_neg_3_port, A4(2) => s_2A_3_neg_2_port, A4(1)
                           => s_2A_3_neg_1_port, A4(0) => s_2A_3_neg_0_port, 
                           SEL(2) => enc_reg32_2_port, SEL(1) => 
                           enc_reg32_1_port, SEL(0) => enc_reg32_0_port, Y(31) 
                           => mux_3_out_31_port, Y(30) => mux_3_out_30_port, 
                           Y(29) => mux_3_out_29_port, Y(28) => 
                           mux_3_out_28_port, Y(27) => mux_3_out_27_port, Y(26)
                           => mux_3_out_26_port, Y(25) => mux_3_out_25_port, 
                           Y(24) => mux_3_out_24_port, Y(23) => 
                           mux_3_out_23_port, Y(22) => mux_3_out_22_port, Y(21)
                           => mux_3_out_21_port, Y(20) => mux_3_out_20_port, 
                           Y(19) => mux_3_out_19_port, Y(18) => 
                           mux_3_out_18_port, Y(17) => mux_3_out_17_port, Y(16)
                           => mux_3_out_16_port, Y(15) => mux_3_out_15_port, 
                           Y(14) => mux_3_out_14_port, Y(13) => 
                           mux_3_out_13_port, Y(12) => mux_3_out_12_port, Y(11)
                           => mux_3_out_11_port, Y(10) => mux_3_out_10_port, 
                           Y(9) => mux_3_out_9_port, Y(8) => mux_3_out_8_port, 
                           Y(7) => mux_3_out_7_port, Y(6) => mux_3_out_6_port, 
                           Y(5) => mux_3_out_5_port, Y(4) => mux_3_out_4_port, 
                           Y(3) => mux_3_out_3_port, Y(2) => mux_3_out_2_port, 
                           Y(1) => mux_3_out_1_port, Y(0) => mux_3_out_0_port);
   SUM2 : P4_ADDER_NBIT64_2 port map( A(63) => sum_reg2_63_port, A(62) => 
                           sum_reg2_62_port, A(61) => sum_reg2_61_port, A(60) 
                           => sum_reg2_60_port, A(59) => sum_reg2_59_port, 
                           A(58) => sum_reg2_58_port, A(57) => sum_reg2_57_port
                           , A(56) => sum_reg2_56_port, A(55) => 
                           sum_reg2_55_port, A(54) => sum_reg2_54_port, A(53) 
                           => sum_reg2_53_port, A(52) => sum_reg2_52_port, 
                           A(51) => sum_reg2_51_port, A(50) => sum_reg2_50_port
                           , A(49) => sum_reg2_49_port, A(48) => 
                           sum_reg2_48_port, A(47) => sum_reg2_47_port, A(46) 
                           => sum_reg2_46_port, A(45) => sum_reg2_45_port, 
                           A(44) => sum_reg2_44_port, A(43) => sum_reg2_43_port
                           , A(42) => sum_reg2_42_port, A(41) => 
                           sum_reg2_41_port, A(40) => sum_reg2_40_port, A(39) 
                           => sum_reg2_39_port, A(38) => sum_reg2_38_port, 
                           A(37) => sum_reg2_37_port, A(36) => sum_reg2_36_port
                           , A(35) => sum_reg2_35_port, A(34) => 
                           sum_reg2_34_port, A(33) => sum_reg2_33_port, A(32) 
                           => sum_reg2_32_port, A(31) => sum_reg2_31_port, 
                           A(30) => sum_reg2_30_port, A(29) => sum_reg2_29_port
                           , A(28) => sum_reg2_28_port, A(27) => 
                           sum_reg2_27_port, A(26) => sum_reg2_26_port, A(25) 
                           => sum_reg2_25_port, A(24) => sum_reg2_24_port, 
                           A(23) => sum_reg2_23_port, A(22) => sum_reg2_22_port
                           , A(21) => sum_reg2_21_port, A(20) => 
                           sum_reg2_20_port, A(19) => sum_reg2_19_port, A(18) 
                           => sum_reg2_18_port, A(17) => sum_reg2_17_port, 
                           A(16) => sum_reg2_16_port, A(15) => sum_reg2_15_port
                           , A(14) => sum_reg2_14_port, A(13) => 
                           sum_reg2_13_port, A(12) => sum_reg2_12_port, A(11) 
                           => sum_reg2_11_port, A(10) => sum_reg2_10_port, A(9)
                           => sum_reg2_9_port, A(8) => sum_reg2_8_port, A(7) =>
                           sum_reg2_7_port, A(6) => sum_reg2_6_port, A(5) => 
                           sum_reg2_5_port, A(4) => sum_reg2_4_port, A(3) => 
                           sum_reg2_3_port, A(2) => sum_reg2_2_port, A(1) => 
                           sum_reg2_1_port, A(0) => sum_reg2_0_port, B(63) => 
                           n6, B(62) => n6, B(61) => n6, B(60) => n6, B(59) => 
                           n6, B(58) => n6, B(57) => n6, B(56) => n6, B(55) => 
                           n6, B(54) => n6, B(53) => n6, B(52) => n5, B(51) => 
                           n5, B(50) => n5, B(49) => n5, B(48) => n5, B(47) => 
                           n5, B(46) => n5, B(45) => n5, B(44) => n5, B(43) => 
                           n5, B(42) => n5, B(41) => n4, B(40) => n4, B(39) => 
                           n4, B(38) => n4, B(37) => n4, B(36) => n4, B(35) => 
                           n4, B(34) => n4, B(33) => n4, B(32) => n4, B(31) => 
                           n4, B(30) => mux_reg2_30_port, B(29) => 
                           mux_reg2_29_port, B(28) => mux_reg2_28_port, B(27) 
                           => mux_reg2_27_port, B(26) => mux_reg2_26_port, 
                           B(25) => mux_reg2_25_port, B(24) => mux_reg2_24_port
                           , B(23) => mux_reg2_23_port, B(22) => 
                           mux_reg2_22_port, B(21) => mux_reg2_21_port, B(20) 
                           => mux_reg2_20_port, B(19) => mux_reg2_19_port, 
                           B(18) => mux_reg2_18_port, B(17) => mux_reg2_17_port
                           , B(16) => mux_reg2_16_port, B(15) => 
                           mux_reg2_15_port, B(14) => mux_reg2_14_port, B(13) 
                           => mux_reg2_13_port, B(12) => mux_reg2_12_port, 
                           B(11) => mux_reg2_11_port, B(10) => mux_reg2_10_port
                           , B(9) => mux_reg2_9_port, B(8) => mux_reg2_8_port, 
                           B(7) => mux_reg2_7_port, B(6) => mux_reg2_6_port, 
                           B(5) => mux_reg2_5_port, B(4) => mux_reg2_4_port, 
                           B(3) => mux_reg2_3_port, B(2) => mux_reg2_2_port, 
                           B(1) => mux_reg2_1_port, B(0) => mux_reg2_0_port, 
                           Cin => X_Logic0_port, S(63) => sum_3_out_63_port, 
                           S(62) => sum_3_out_62_port, S(61) => 
                           sum_3_out_61_port, S(60) => sum_3_out_60_port, S(59)
                           => sum_3_out_59_port, S(58) => sum_3_out_58_port, 
                           S(57) => sum_3_out_57_port, S(56) => 
                           sum_3_out_56_port, S(55) => sum_3_out_55_port, S(54)
                           => sum_3_out_54_port, S(53) => sum_3_out_53_port, 
                           S(52) => sum_3_out_52_port, S(51) => 
                           sum_3_out_51_port, S(50) => sum_3_out_50_port, S(49)
                           => sum_3_out_49_port, S(48) => sum_3_out_48_port, 
                           S(47) => sum_3_out_47_port, S(46) => 
                           sum_3_out_46_port, S(45) => sum_3_out_45_port, S(44)
                           => sum_3_out_44_port, S(43) => sum_3_out_43_port, 
                           S(42) => sum_3_out_42_port, S(41) => 
                           sum_3_out_41_port, S(40) => sum_3_out_40_port, S(39)
                           => sum_3_out_39_port, S(38) => sum_3_out_38_port, 
                           S(37) => sum_3_out_37_port, S(36) => 
                           sum_3_out_36_port, S(35) => sum_3_out_35_port, S(34)
                           => sum_3_out_34_port, S(33) => sum_3_out_33_port, 
                           S(32) => sum_3_out_32_port, S(31) => 
                           sum_3_out_31_port, S(30) => sum_3_out_30_port, S(29)
                           => sum_3_out_29_port, S(28) => sum_3_out_28_port, 
                           S(27) => sum_3_out_27_port, S(26) => 
                           sum_3_out_26_port, S(25) => sum_3_out_25_port, S(24)
                           => sum_3_out_24_port, S(23) => sum_3_out_23_port, 
                           S(22) => sum_3_out_22_port, S(21) => 
                           sum_3_out_21_port, S(20) => sum_3_out_20_port, S(19)
                           => sum_3_out_19_port, S(18) => sum_3_out_18_port, 
                           S(17) => sum_3_out_17_port, S(16) => 
                           sum_3_out_16_port, S(15) => sum_3_out_15_port, S(14)
                           => sum_3_out_14_port, S(13) => sum_3_out_13_port, 
                           S(12) => sum_3_out_12_port, S(11) => 
                           sum_3_out_11_port, S(10) => sum_3_out_10_port, S(9) 
                           => sum_3_out_9_port, S(8) => sum_3_out_8_port, S(7) 
                           => sum_3_out_7_port, S(6) => sum_3_out_6_port, S(5) 
                           => sum_3_out_5_port, S(4) => sum_3_out_4_port, S(3) 
                           => sum_3_out_3_port, S(2) => sum_3_out_2_port, S(1) 
                           => sum_3_out_1_port, S(0) => sum_3_out_0_port, Cout 
                           => n_1916, ovf => n_1917);
   SUM3 : P4_ADDER_NBIT64_1 port map( A(63) => sum_reg3_63_port, A(62) => 
                           sum_reg3_62_port, A(61) => sum_reg3_61_port, A(60) 
                           => sum_reg3_60_port, A(59) => sum_reg3_59_port, 
                           A(58) => sum_reg3_58_port, A(57) => sum_reg3_57_port
                           , A(56) => sum_reg3_56_port, A(55) => 
                           sum_reg3_55_port, A(54) => sum_reg3_54_port, A(53) 
                           => sum_reg3_53_port, A(52) => sum_reg3_52_port, 
                           A(51) => sum_reg3_51_port, A(50) => sum_reg3_50_port
                           , A(49) => sum_reg3_49_port, A(48) => 
                           sum_reg3_48_port, A(47) => sum_reg3_47_port, A(46) 
                           => sum_reg3_46_port, A(45) => sum_reg3_45_port, 
                           A(44) => sum_reg3_44_port, A(43) => sum_reg3_43_port
                           , A(42) => sum_reg3_42_port, A(41) => 
                           sum_reg3_41_port, A(40) => sum_reg3_40_port, A(39) 
                           => sum_reg3_39_port, A(38) => sum_reg3_38_port, 
                           A(37) => sum_reg3_37_port, A(36) => sum_reg3_36_port
                           , A(35) => sum_reg3_35_port, A(34) => 
                           sum_reg3_34_port, A(33) => sum_reg3_33_port, A(32) 
                           => sum_reg3_32_port, A(31) => sum_reg3_31_port, 
                           A(30) => sum_reg3_30_port, A(29) => sum_reg3_29_port
                           , A(28) => sum_reg3_28_port, A(27) => 
                           sum_reg3_27_port, A(26) => sum_reg3_26_port, A(25) 
                           => sum_reg3_25_port, A(24) => sum_reg3_24_port, 
                           A(23) => sum_reg3_23_port, A(22) => sum_reg3_22_port
                           , A(21) => sum_reg3_21_port, A(20) => 
                           sum_reg3_20_port, A(19) => sum_reg3_19_port, A(18) 
                           => sum_reg3_18_port, A(17) => sum_reg3_17_port, 
                           A(16) => sum_reg3_16_port, A(15) => sum_reg3_15_port
                           , A(14) => sum_reg3_14_port, A(13) => 
                           sum_reg3_13_port, A(12) => sum_reg3_12_port, A(11) 
                           => sum_reg3_11_port, A(10) => sum_reg3_10_port, A(9)
                           => sum_reg3_9_port, A(8) => sum_reg3_8_port, A(7) =>
                           sum_reg3_7_port, A(6) => sum_reg3_6_port, A(5) => 
                           sum_reg3_5_port, A(4) => sum_reg3_4_port, A(3) => 
                           sum_reg3_3_port, A(2) => sum_reg3_2_port, A(1) => 
                           sum_reg3_1_port, A(0) => sum_reg3_0_port, B(63) => 
                           n3, B(62) => n3, B(61) => n3, B(60) => n3, B(59) => 
                           n3, B(58) => n3, B(57) => n3, B(56) => n3, B(55) => 
                           n3, B(54) => n3, B(53) => n3, B(52) => n2, B(51) => 
                           n2, B(50) => n2, B(49) => n2, B(48) => n2, B(47) => 
                           n2, B(46) => n2, B(45) => n2, B(44) => n2, B(43) => 
                           n2, B(42) => n2, B(41) => n1, B(40) => n1, B(39) => 
                           n1, B(38) => n1, B(37) => n1, B(36) => n1, B(35) => 
                           n1, B(34) => n1, B(33) => n1, B(32) => n1, B(31) => 
                           n1, B(30) => mux_reg3_30_port, B(29) => 
                           mux_reg3_29_port, B(28) => mux_reg3_28_port, B(27) 
                           => mux_reg3_27_port, B(26) => mux_reg3_26_port, 
                           B(25) => mux_reg3_25_port, B(24) => mux_reg3_24_port
                           , B(23) => mux_reg3_23_port, B(22) => 
                           mux_reg3_22_port, B(21) => mux_reg3_21_port, B(20) 
                           => mux_reg3_20_port, B(19) => mux_reg3_19_port, 
                           B(18) => mux_reg3_18_port, B(17) => mux_reg3_17_port
                           , B(16) => mux_reg3_16_port, B(15) => 
                           mux_reg3_15_port, B(14) => mux_reg3_14_port, B(13) 
                           => mux_reg3_13_port, B(12) => mux_reg3_12_port, 
                           B(11) => mux_reg3_11_port, B(10) => mux_reg3_10_port
                           , B(9) => mux_reg3_9_port, B(8) => mux_reg3_8_port, 
                           B(7) => mux_reg3_7_port, B(6) => mux_reg3_6_port, 
                           B(5) => mux_reg3_5_port, B(4) => mux_reg3_4_port, 
                           B(3) => mux_reg3_3_port, B(2) => mux_reg3_2_port, 
                           B(1) => mux_reg3_1_port, B(0) => mux_reg3_0_port, 
                           Cin => X_Logic0_port, S(63) => P(63), S(62) => P(62)
                           , S(61) => P(61), S(60) => P(60), S(59) => P(59), 
                           S(58) => P(58), S(57) => P(57), S(56) => P(56), 
                           S(55) => P(55), S(54) => P(54), S(53) => P(53), 
                           S(52) => P(52), S(51) => P(51), S(50) => P(50), 
                           S(49) => P(49), S(48) => P(48), S(47) => P(47), 
                           S(46) => P(46), S(45) => P(45), S(44) => P(44), 
                           S(43) => P(43), S(42) => P(42), S(41) => P(41), 
                           S(40) => P(40), S(39) => P(39), S(38) => P(38), 
                           S(37) => P(37), S(36) => P(36), S(35) => P(35), 
                           S(34) => P(34), S(33) => P(33), S(32) => P(32), 
                           S(31) => P(31), S(30) => P(30), S(29) => P(29), 
                           S(28) => P(28), S(27) => P(27), S(26) => P(26), 
                           S(25) => P(25), S(24) => P(24), S(23) => P(23), 
                           S(22) => P(22), S(21) => P(21), S(20) => P(20), 
                           S(19) => P(19), S(18) => P(18), S(17) => P(17), 
                           S(16) => P(16), S(15) => P(15), S(14) => P(14), 
                           S(13) => P(13), S(12) => P(12), S(11) => P(11), 
                           S(10) => P(10), S(9) => P(9), S(8) => P(8), S(7) => 
                           P(7), S(6) => P(6), S(5) => P(5), S(4) => P(4), S(3)
                           => P(3), S(2) => P(2), S(1) => P(1), S(0) => P(0), 
                           Cout => n_1918, ovf => n_1919);
   U3 : BUF_X1 port map( A => n28, Z => n21);
   U4 : BUF_X1 port map( A => n28, Z => n22);
   U5 : BUF_X1 port map( A => n28, Z => n23);
   U6 : BUF_X1 port map( A => n27, Z => n24);
   U7 : BUF_X1 port map( A => n27, Z => n25);
   U8 : BUF_X1 port map( A => n29, Z => n19);
   U9 : BUF_X1 port map( A => n29, Z => n20);
   U10 : BUF_X1 port map( A => n27, Z => n26);
   U11 : BUF_X1 port map( A => RST, Z => n28);
   U12 : BUF_X1 port map( A => RST, Z => n27);
   U13 : BUF_X1 port map( A => RST, Z => n29);
   U14 : BUF_X2 port map( A => n11, Z => n15);
   U15 : BUF_X2 port map( A => n10, Z => n13);
   U16 : BUF_X2 port map( A => n11, Z => n16);
   U17 : BUF_X2 port map( A => n10, Z => n14);
   U18 : BUF_X2 port map( A => n10, Z => n12);
   U19 : BUF_X2 port map( A => n11, Z => n17);
   U20 : BUF_X1 port map( A => A(31), Z => n18);
   U21 : BUF_X1 port map( A => mux_reg2_31_port, Z => n5);
   U22 : BUF_X1 port map( A => mux_reg2_31_port, Z => n4);
   U23 : BUF_X1 port map( A => mux2_reg1_31_port, Z => n7);
   U24 : BUF_X1 port map( A => mux2_reg1_31_port, Z => n8);
   U25 : BUF_X1 port map( A => mux2_reg1_31_port, Z => n9);
   U26 : BUF_X1 port map( A => mux_reg2_31_port, Z => n6);
   U27 : BUF_X1 port map( A => mux1_reg1_31_port, Z => n11);
   U28 : BUF_X1 port map( A => mux1_reg1_31_port, Z => n10);
   U29 : BUF_X1 port map( A => mux_reg3_31_port, Z => n1);
   U30 : BUF_X1 port map( A => mux_reg3_31_port, Z => n2);
   U31 : BUF_X1 port map( A => mux_reg3_31_port, Z => n3);
   A4_reg1_2_port <= '0';
   A4_reg1_1_port <= '0';
   A4_reg1_0_port <= '0';
   A4_reg2_1_port <= '0';
   A4_reg2_0_port <= '0';
   U37 : CLKBUF_X1 port map( A => n19, Z => n30);
   U38 : CLKBUF_X1 port map( A => n19, Z => n31);
   U39 : CLKBUF_X1 port map( A => n19, Z => n32);
   U40 : CLKBUF_X1 port map( A => n19, Z => n33);
   U41 : CLKBUF_X1 port map( A => n20, Z => n34);
   U42 : CLKBUF_X1 port map( A => n20, Z => n35);
   U43 : CLKBUF_X1 port map( A => n20, Z => n36);
   U44 : CLKBUF_X1 port map( A => n20, Z => n37);
   U45 : CLKBUF_X1 port map( A => n21, Z => n38);
   U46 : CLKBUF_X1 port map( A => n21, Z => n39);
   U47 : CLKBUF_X1 port map( A => n21, Z => n40);
   U48 : CLKBUF_X1 port map( A => n21, Z => n41);
   U49 : CLKBUF_X1 port map( A => n22, Z => n42);
   U50 : CLKBUF_X1 port map( A => n22, Z => n43);
   U51 : CLKBUF_X1 port map( A => n22, Z => n44);
   U52 : CLKBUF_X1 port map( A => n22, Z => n45);
   U53 : CLKBUF_X1 port map( A => n23, Z => n46);
   U54 : CLKBUF_X1 port map( A => n23, Z => n47);
   U55 : CLKBUF_X1 port map( A => n23, Z => n48);
   U56 : CLKBUF_X1 port map( A => n23, Z => n49);
   U57 : CLKBUF_X1 port map( A => n24, Z => n50);
   U58 : CLKBUF_X1 port map( A => n24, Z => n51);
   U59 : CLKBUF_X1 port map( A => n24, Z => n52);
   U60 : CLKBUF_X1 port map( A => n24, Z => n53);
   U61 : CLKBUF_X1 port map( A => n25, Z => n54);
   U62 : CLKBUF_X1 port map( A => n25, Z => n55);
   U63 : CLKBUF_X1 port map( A => n25, Z => n56);
   U64 : CLKBUF_X1 port map( A => n25, Z => n57);
   U65 : CLKBUF_X1 port map( A => n26, Z => n58);
   U66 : CLKBUF_X1 port map( A => n26, Z => n59);
   U67 : CLKBUF_X1 port map( A => n26, Z => n60);
   s_2A_2_0_port <= '0';
   s_2A_2_1_port <= '0';
   s_2A_3_0_port <= '0';
   s_2A_3_1_port <= '0';
   s_A_2_0_port <= '0';
   s_A_3_0_port <= '0';
   s_8A_1_0_port <= '0';
   s_8A_1_1_port <= '0';
   s_8A_1_2_port <= '0';
   s_4A_1_0_port <= '0';
   s_4A_1_1_port <= '0';
   s_2A_1_0_port <= '0';

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity ALU_N32 is

   port( DATA1, DATA2 : in std_logic_vector (31 downto 0);  FUNC : in 
         std_logic_vector (3 downto 0);  SN : in std_logic;  OVF : out 
         std_logic;  OUTALU : out std_logic_vector (31 downto 0));

end ALU_N32;

architecture SYN_BEHAVIOR of ALU_N32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component comparator
      port( Z, cout : in std_logic;  eq, neq, gt, lt, ge, le : out std_logic);
   end component;
   
   component nor_generic_NBITS32
      port( input : in std_logic_vector (31 downto 0);  result : out std_logic
            );
   end component;
   
   component logicals_nbit32
      port( func : in std_logic_vector (3 downto 0);  SN : in std_logic;  in1, 
            in2 : in std_logic_vector (31 downto 0);  o : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component P4_ADDER_NBIT32_1
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  S :
            out std_logic_vector (31 downto 0);  Cout, ovf : out std_logic);
   end component;
   
   component shifter_NBITS32
      port( R1, R2 : in std_logic_vector (31 downto 0);  LnR, AnL, RnS : in 
            std_logic;  Rout : out std_logic_vector (31 downto 0));
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal s_LnR, s_AnL, s_RnS, shifter_out_31_port, shifter_out_30_port, 
      shifter_out_29_port, shifter_out_28_port, shifter_out_27_port, 
      shifter_out_26_port, shifter_out_25_port, shifter_out_24_port, 
      shifter_out_23_port, shifter_out_22_port, shifter_out_21_port, 
      shifter_out_20_port, shifter_out_19_port, shifter_out_18_port, 
      shifter_out_17_port, shifter_out_16_port, shifter_out_15_port, 
      shifter_out_14_port, shifter_out_13_port, shifter_out_12_port, 
      shifter_out_11_port, shifter_out_10_port, shifter_out_9_port, 
      shifter_out_8_port, shifter_out_7_port, shifter_out_6_port, 
      shifter_out_5_port, shifter_out_4_port, shifter_out_3_port, 
      shifter_out_2_port, shifter_out_1_port, shifter_out_0_port, p4_cin, 
      p4_sum_31_port, p4_sum_30_port, p4_sum_29_port, p4_sum_28_port, 
      p4_sum_27_port, p4_sum_26_port, p4_sum_25_port, p4_sum_24_port, 
      p4_sum_23_port, p4_sum_22_port, p4_sum_21_port, p4_sum_20_port, 
      p4_sum_19_port, p4_sum_18_port, p4_sum_17_port, p4_sum_16_port, 
      p4_sum_15_port, p4_sum_14_port, p4_sum_13_port, p4_sum_12_port, 
      p4_sum_11_port, p4_sum_10_port, p4_sum_9_port, p4_sum_8_port, 
      p4_sum_7_port, p4_sum_6_port, p4_sum_5_port, p4_sum_4_port, p4_sum_3_port
      , p4_sum_2_port, p4_sum_1_port, p4_sum_0_port, p4_cout, p4_ovf, 
      logic_func_3_port, logic_func_2_port, logic_func_1_port, 
      logic_func_0_port, logic_out_31_port, logic_out_30_port, 
      logic_out_29_port, logic_out_28_port, logic_out_27_port, 
      logic_out_26_port, logic_out_25_port, logic_out_24_port, 
      logic_out_23_port, logic_out_22_port, logic_out_21_port, 
      logic_out_20_port, logic_out_19_port, logic_out_18_port, 
      logic_out_17_port, logic_out_16_port, logic_out_15_port, 
      logic_out_14_port, logic_out_13_port, logic_out_12_port, 
      logic_out_11_port, logic_out_10_port, logic_out_9_port, logic_out_8_port,
      logic_out_7_port, logic_out_6_port, logic_out_5_port, logic_out_4_port, 
      logic_out_3_port, logic_out_2_port, logic_out_1_port, logic_out_0_port, 
      is_zero, s_eq, s_neq, s_gt, s_lt, N74, N75, N76, N77, N78, n44, n45, n46,
      n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61
      , n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74_port, 
      n75_port, n76_port, n77_port, n78_port, n79, n80, n81, n82, n83, n84, n85
      , n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, 
      n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n42, n43, n100, n101, n102, n103
      , n104, n105, n106, n107, n_1920, n_1921 : std_logic;

begin
   
   s_RnS_reg : DLH_X1 port map( G => n3, D => n97, Q => s_RnS);
   p4_cin_reg : DLH_X1 port map( G => N74, D => N75, Q => p4_cin);
   OVF_reg : DLH_X1 port map( G => n9, D => p4_ovf, Q => OVF);
   logic_func_reg_3_inst : DLH_X1 port map( G => n6, D => FUNC(3), Q => 
                           logic_func_3_port);
   logic_func_reg_2_inst : DLH_X1 port map( G => n6, D => FUNC(2), Q => 
                           logic_func_2_port);
   logic_func_reg_1_inst : DLH_X1 port map( G => n6, D => FUNC(1), Q => 
                           logic_func_1_port);
   logic_func_reg_0_inst : DLH_X1 port map( G => n6, D => FUNC(0), Q => 
                           logic_func_0_port);
   s_LnR_reg : DLH_X1 port map( G => n3, D => n98, Q => s_LnR);
   s_AnL_reg : DLH_X1 port map( G => n3, D => n99, Q => s_AnL);
   U102 : NAND3_X1 port map( A1 => n78_port, A2 => n79, A3 => n80, ZN => 
                           OUTALU(0));
   U103 : XOR2_X1 port map( A => DATA2(31), B => n10, Z => n94);
   U104 : NAND3_X1 port map( A1 => FUNC(1), A2 => n107, A3 => FUNC(2), ZN => 
                           n44);
   U105 : OAI33_X1 port map( A1 => n106, A2 => FUNC(3), A3 => FUNC(2), B1 => 
                           n46, B2 => FUNC(1), B3 => FUNC(0), ZN => N77);
   U106 : NAND3_X1 port map( A1 => FUNC(3), A2 => FUNC(2), A3 => n105, ZN => 
                           n88);
   alu_shifter : shifter_NBITS32 port map( R1(31) => n10, R1(30) => DATA1(30), 
                           R1(29) => DATA1(29), R1(28) => DATA1(28), R1(27) => 
                           DATA1(27), R1(26) => DATA1(26), R1(25) => DATA1(25),
                           R1(24) => DATA1(24), R1(23) => DATA1(23), R1(22) => 
                           DATA1(22), R1(21) => DATA1(21), R1(20) => DATA1(20),
                           R1(19) => DATA1(19), R1(18) => DATA1(18), R1(17) => 
                           DATA1(17), R1(16) => DATA1(16), R1(15) => DATA1(15),
                           R1(14) => DATA1(14), R1(13) => DATA1(13), R1(12) => 
                           DATA1(12), R1(11) => DATA1(11), R1(10) => DATA1(10),
                           R1(9) => DATA1(9), R1(8) => DATA1(8), R1(7) => 
                           DATA1(7), R1(6) => DATA1(6), R1(5) => DATA1(5), 
                           R1(4) => DATA1(4), R1(3) => DATA1(3), R1(2) => 
                           DATA1(2), R1(1) => DATA1(1), R1(0) => DATA1(0), 
                           R2(31) => DATA2(31), R2(30) => DATA2(30), R2(29) => 
                           DATA2(29), R2(28) => DATA2(28), R2(27) => DATA2(27),
                           R2(26) => DATA2(26), R2(25) => DATA2(25), R2(24) => 
                           DATA2(24), R2(23) => DATA2(23), R2(22) => DATA2(22),
                           R2(21) => DATA2(21), R2(20) => DATA2(20), R2(19) => 
                           DATA2(19), R2(18) => DATA2(18), R2(17) => DATA2(17),
                           R2(16) => DATA2(16), R2(15) => DATA2(15), R2(14) => 
                           DATA2(14), R2(13) => DATA2(13), R2(12) => DATA2(12),
                           R2(11) => DATA2(11), R2(10) => DATA2(10), R2(9) => 
                           DATA2(9), R2(8) => DATA2(8), R2(7) => DATA2(7), 
                           R2(6) => DATA2(6), R2(5) => DATA2(5), R2(4) => 
                           DATA2(4), R2(3) => DATA2(3), R2(2) => DATA2(2), 
                           R2(1) => DATA2(1), R2(0) => DATA2(0), LnR => s_LnR, 
                           AnL => s_AnL, RnS => s_RnS, Rout(31) => 
                           shifter_out_31_port, Rout(30) => shifter_out_30_port
                           , Rout(29) => shifter_out_29_port, Rout(28) => 
                           shifter_out_28_port, Rout(27) => shifter_out_27_port
                           , Rout(26) => shifter_out_26_port, Rout(25) => 
                           shifter_out_25_port, Rout(24) => shifter_out_24_port
                           , Rout(23) => shifter_out_23_port, Rout(22) => 
                           shifter_out_22_port, Rout(21) => shifter_out_21_port
                           , Rout(20) => shifter_out_20_port, Rout(19) => 
                           shifter_out_19_port, Rout(18) => shifter_out_18_port
                           , Rout(17) => shifter_out_17_port, Rout(16) => 
                           shifter_out_16_port, Rout(15) => shifter_out_15_port
                           , Rout(14) => shifter_out_14_port, Rout(13) => 
                           shifter_out_13_port, Rout(12) => shifter_out_12_port
                           , Rout(11) => shifter_out_11_port, Rout(10) => 
                           shifter_out_10_port, Rout(9) => shifter_out_9_port, 
                           Rout(8) => shifter_out_8_port, Rout(7) => 
                           shifter_out_7_port, Rout(6) => shifter_out_6_port, 
                           Rout(5) => shifter_out_5_port, Rout(4) => 
                           shifter_out_4_port, Rout(3) => shifter_out_3_port, 
                           Rout(2) => shifter_out_2_port, Rout(1) => 
                           shifter_out_1_port, Rout(0) => shifter_out_0_port);
   alu_adder : P4_ADDER_NBIT32_1 port map( A(31) => n10, A(30) => DATA1(30), 
                           A(29) => DATA1(29), A(28) => DATA1(28), A(27) => 
                           DATA1(27), A(26) => DATA1(26), A(25) => DATA1(25), 
                           A(24) => DATA1(24), A(23) => DATA1(23), A(22) => 
                           DATA1(22), A(21) => DATA1(21), A(20) => DATA1(20), 
                           A(19) => DATA1(19), A(18) => DATA1(18), A(17) => 
                           DATA1(17), A(16) => DATA1(16), A(15) => DATA1(15), 
                           A(14) => DATA1(14), A(13) => DATA1(13), A(12) => 
                           DATA1(12), A(11) => DATA1(11), A(10) => DATA1(10), 
                           A(9) => DATA1(9), A(8) => DATA1(8), A(7) => DATA1(7)
                           , A(6) => DATA1(6), A(5) => DATA1(5), A(4) => 
                           DATA1(4), A(3) => DATA1(3), A(2) => DATA1(2), A(1) 
                           => DATA1(1), A(0) => DATA1(0), B(31) => DATA2(31), 
                           B(30) => DATA2(30), B(29) => DATA2(29), B(28) => 
                           DATA2(28), B(27) => DATA2(27), B(26) => DATA2(26), 
                           B(25) => DATA2(25), B(24) => DATA2(24), B(23) => 
                           DATA2(23), B(22) => DATA2(22), B(21) => DATA2(21), 
                           B(20) => DATA2(20), B(19) => DATA2(19), B(18) => 
                           DATA2(18), B(17) => DATA2(17), B(16) => DATA2(16), 
                           B(15) => DATA2(15), B(14) => DATA2(14), B(13) => 
                           DATA2(13), B(12) => DATA2(12), B(11) => DATA2(11), 
                           B(10) => DATA2(10), B(9) => DATA2(9), B(8) => 
                           DATA2(8), B(7) => DATA2(7), B(6) => DATA2(6), B(5) 
                           => DATA2(5), B(4) => DATA2(4), B(3) => DATA2(3), 
                           B(2) => DATA2(2), B(1) => DATA2(1), B(0) => DATA2(0)
                           , Cin => p4_cin, S(31) => p4_sum_31_port, S(30) => 
                           p4_sum_30_port, S(29) => p4_sum_29_port, S(28) => 
                           p4_sum_28_port, S(27) => p4_sum_27_port, S(26) => 
                           p4_sum_26_port, S(25) => p4_sum_25_port, S(24) => 
                           p4_sum_24_port, S(23) => p4_sum_23_port, S(22) => 
                           p4_sum_22_port, S(21) => p4_sum_21_port, S(20) => 
                           p4_sum_20_port, S(19) => p4_sum_19_port, S(18) => 
                           p4_sum_18_port, S(17) => p4_sum_17_port, S(16) => 
                           p4_sum_16_port, S(15) => p4_sum_15_port, S(14) => 
                           p4_sum_14_port, S(13) => p4_sum_13_port, S(12) => 
                           p4_sum_12_port, S(11) => p4_sum_11_port, S(10) => 
                           p4_sum_10_port, S(9) => p4_sum_9_port, S(8) => 
                           p4_sum_8_port, S(7) => p4_sum_7_port, S(6) => 
                           p4_sum_6_port, S(5) => p4_sum_5_port, S(4) => 
                           p4_sum_4_port, S(3) => p4_sum_3_port, S(2) => 
                           p4_sum_2_port, S(1) => p4_sum_1_port, S(0) => 
                           p4_sum_0_port, Cout => p4_cout, ovf => p4_ovf);
   alu_logicals : logicals_nbit32 port map( func(3) => logic_func_3_port, 
                           func(2) => logic_func_2_port, func(1) => 
                           logic_func_1_port, func(0) => logic_func_0_port, SN 
                           => SN, in1(31) => n10, in1(30) => DATA1(30), in1(29)
                           => DATA1(29), in1(28) => DATA1(28), in1(27) => 
                           DATA1(27), in1(26) => DATA1(26), in1(25) => 
                           DATA1(25), in1(24) => DATA1(24), in1(23) => 
                           DATA1(23), in1(22) => DATA1(22), in1(21) => 
                           DATA1(21), in1(20) => DATA1(20), in1(19) => 
                           DATA1(19), in1(18) => DATA1(18), in1(17) => 
                           DATA1(17), in1(16) => DATA1(16), in1(15) => 
                           DATA1(15), in1(14) => DATA1(14), in1(13) => 
                           DATA1(13), in1(12) => DATA1(12), in1(11) => 
                           DATA1(11), in1(10) => DATA1(10), in1(9) => DATA1(9),
                           in1(8) => DATA1(8), in1(7) => DATA1(7), in1(6) => 
                           DATA1(6), in1(5) => DATA1(5), in1(4) => DATA1(4), 
                           in1(3) => DATA1(3), in1(2) => DATA1(2), in1(1) => 
                           DATA1(1), in1(0) => DATA1(0), in2(31) => DATA2(31), 
                           in2(30) => DATA2(30), in2(29) => DATA2(29), in2(28) 
                           => DATA2(28), in2(27) => DATA2(27), in2(26) => 
                           DATA2(26), in2(25) => DATA2(25), in2(24) => 
                           DATA2(24), in2(23) => DATA2(23), in2(22) => 
                           DATA2(22), in2(21) => DATA2(21), in2(20) => 
                           DATA2(20), in2(19) => DATA2(19), in2(18) => 
                           DATA2(18), in2(17) => DATA2(17), in2(16) => 
                           DATA2(16), in2(15) => DATA2(15), in2(14) => 
                           DATA2(14), in2(13) => DATA2(13), in2(12) => 
                           DATA2(12), in2(11) => DATA2(11), in2(10) => 
                           DATA2(10), in2(9) => DATA2(9), in2(8) => DATA2(8), 
                           in2(7) => DATA2(7), in2(6) => DATA2(6), in2(5) => 
                           DATA2(5), in2(4) => DATA2(4), in2(3) => DATA2(3), 
                           in2(2) => DATA2(2), in2(1) => DATA2(1), in2(0) => 
                           DATA2(0), o(31) => logic_out_31_port, o(30) => 
                           logic_out_30_port, o(29) => logic_out_29_port, o(28)
                           => logic_out_28_port, o(27) => logic_out_27_port, 
                           o(26) => logic_out_26_port, o(25) => 
                           logic_out_25_port, o(24) => logic_out_24_port, o(23)
                           => logic_out_23_port, o(22) => logic_out_22_port, 
                           o(21) => logic_out_21_port, o(20) => 
                           logic_out_20_port, o(19) => logic_out_19_port, o(18)
                           => logic_out_18_port, o(17) => logic_out_17_port, 
                           o(16) => logic_out_16_port, o(15) => 
                           logic_out_15_port, o(14) => logic_out_14_port, o(13)
                           => logic_out_13_port, o(12) => logic_out_12_port, 
                           o(11) => logic_out_11_port, o(10) => 
                           logic_out_10_port, o(9) => logic_out_9_port, o(8) =>
                           logic_out_8_port, o(7) => logic_out_7_port, o(6) => 
                           logic_out_6_port, o(5) => logic_out_5_port, o(4) => 
                           logic_out_4_port, o(3) => logic_out_3_port, o(2) => 
                           logic_out_2_port, o(1) => logic_out_1_port, o(0) => 
                           logic_out_0_port);
   nor_gen : nor_generic_NBITS32 port map( input(31) => p4_sum_31_port, 
                           input(30) => p4_sum_30_port, input(29) => 
                           p4_sum_29_port, input(28) => p4_sum_28_port, 
                           input(27) => p4_sum_27_port, input(26) => 
                           p4_sum_26_port, input(25) => p4_sum_25_port, 
                           input(24) => p4_sum_24_port, input(23) => 
                           p4_sum_23_port, input(22) => p4_sum_22_port, 
                           input(21) => p4_sum_21_port, input(20) => 
                           p4_sum_20_port, input(19) => p4_sum_19_port, 
                           input(18) => p4_sum_18_port, input(17) => 
                           p4_sum_17_port, input(16) => p4_sum_16_port, 
                           input(15) => p4_sum_15_port, input(14) => 
                           p4_sum_14_port, input(13) => p4_sum_13_port, 
                           input(12) => p4_sum_12_port, input(11) => 
                           p4_sum_11_port, input(10) => p4_sum_10_port, 
                           input(9) => p4_sum_9_port, input(8) => p4_sum_8_port
                           , input(7) => p4_sum_7_port, input(6) => 
                           p4_sum_6_port, input(5) => p4_sum_5_port, input(4) 
                           => p4_sum_4_port, input(3) => p4_sum_3_port, 
                           input(2) => p4_sum_2_port, input(1) => p4_sum_1_port
                           , input(0) => p4_sum_0_port, result => is_zero);
   comp : comparator port map( Z => is_zero, cout => p4_cout, eq => s_eq, neq 
                           => s_neq, gt => s_gt, lt => s_lt, ge => n_1920, le 
                           => n_1921);
   U2 : INV_X1 port map( A => n64, ZN => OUTALU(22));
   U3 : AOI222_X1 port map( A1 => shifter_out_22_port, A2 => n2, B1 => 
                           p4_sum_22_port, B2 => n8, C1 => logic_out_22_port, 
                           C2 => n5, ZN => n64);
   U4 : INV_X1 port map( A => n65, ZN => OUTALU(21));
   U5 : AOI222_X1 port map( A1 => shifter_out_21_port, A2 => n2, B1 => 
                           p4_sum_21_port, B2 => n8, C1 => logic_out_21_port, 
                           C2 => n5, ZN => n65);
   U6 : INV_X1 port map( A => n68, ZN => OUTALU(19));
   U7 : AOI222_X1 port map( A1 => shifter_out_19_port, A2 => n2, B1 => 
                           p4_sum_19_port, B2 => n8, C1 => logic_out_19_port, 
                           C2 => n5, ZN => n68);
   U8 : INV_X1 port map( A => n72, ZN => OUTALU(15));
   U9 : AOI222_X1 port map( A1 => shifter_out_15_port, A2 => n3, B1 => 
                           p4_sum_15_port, B2 => n9, C1 => logic_out_15_port, 
                           C2 => n6, ZN => n72);
   U10 : INV_X1 port map( A => n73, ZN => OUTALU(14));
   U11 : AOI222_X1 port map( A1 => shifter_out_14_port, A2 => n3, B1 => 
                           p4_sum_14_port, B2 => n9, C1 => logic_out_14_port, 
                           C2 => n6, ZN => n73);
   U12 : INV_X1 port map( A => n74_port, ZN => OUTALU(13));
   U13 : AOI222_X1 port map( A1 => shifter_out_13_port, A2 => n3, B1 => 
                           p4_sum_13_port, B2 => n9, C1 => logic_out_13_port, 
                           C2 => n6, ZN => n74_port);
   U14 : INV_X1 port map( A => n76_port, ZN => OUTALU(11));
   U15 : AOI222_X1 port map( A1 => shifter_out_11_port, A2 => n3, B1 => 
                           p4_sum_11_port, B2 => n9, C1 => logic_out_11_port, 
                           C2 => n6, ZN => n76_port);
   U16 : INV_X1 port map( A => n77_port, ZN => OUTALU(10));
   U17 : AOI222_X1 port map( A1 => shifter_out_10_port, A2 => n3, B1 => 
                           p4_sum_10_port, B2 => n9, C1 => logic_out_10_port, 
                           C2 => n6, ZN => n77_port);
   U18 : INV_X1 port map( A => n54, ZN => OUTALU(31));
   U19 : AOI222_X1 port map( A1 => shifter_out_31_port, A2 => n1, B1 => 
                           p4_sum_31_port, B2 => n7, C1 => logic_out_31_port, 
                           C2 => n4, ZN => n54);
   U20 : INV_X1 port map( A => n55, ZN => OUTALU(30));
   U21 : AOI222_X1 port map( A1 => shifter_out_30_port, A2 => n1, B1 => 
                           p4_sum_30_port, B2 => n7, C1 => logic_out_30_port, 
                           C2 => n4, ZN => n55);
   U22 : INV_X1 port map( A => n57, ZN => OUTALU(29));
   U23 : AOI222_X1 port map( A1 => shifter_out_29_port, A2 => n1, B1 => 
                           p4_sum_29_port, B2 => n7, C1 => logic_out_29_port, 
                           C2 => n4, ZN => n57);
   U24 : INV_X1 port map( A => n59, ZN => OUTALU(27));
   U25 : AOI222_X1 port map( A1 => shifter_out_27_port, A2 => n2, B1 => 
                           p4_sum_27_port, B2 => n8, C1 => logic_out_27_port, 
                           C2 => n5, ZN => n59);
   U26 : INV_X1 port map( A => n60, ZN => OUTALU(26));
   U27 : AOI222_X1 port map( A1 => shifter_out_26_port, A2 => n2, B1 => 
                           p4_sum_26_port, B2 => n8, C1 => logic_out_26_port, 
                           C2 => n5, ZN => n60);
   U28 : INV_X1 port map( A => n61, ZN => OUTALU(25));
   U29 : AOI222_X1 port map( A1 => shifter_out_25_port, A2 => n2, B1 => 
                           p4_sum_25_port, B2 => n8, C1 => logic_out_25_port, 
                           C2 => n5, ZN => n61);
   U30 : INV_X1 port map( A => n63, ZN => OUTALU(23));
   U31 : AOI222_X1 port map( A1 => shifter_out_23_port, A2 => n2, B1 => 
                           p4_sum_23_port, B2 => n8, C1 => logic_out_23_port, 
                           C2 => n5, ZN => n63);
   U32 : INV_X1 port map( A => n69, ZN => OUTALU(18));
   U33 : AOI222_X1 port map( A1 => shifter_out_18_port, A2 => n2, B1 => 
                           p4_sum_18_port, B2 => n8, C1 => logic_out_18_port, 
                           C2 => n5, ZN => n69);
   U34 : INV_X1 port map( A => n47, ZN => OUTALU(9));
   U35 : AOI222_X1 port map( A1 => shifter_out_9_port, A2 => n2, B1 => 
                           p4_sum_9_port, B2 => n8, C1 => logic_out_9_port, C2 
                           => n5, ZN => n47);
   U36 : INV_X1 port map( A => n49, ZN => OUTALU(7));
   U37 : AOI222_X1 port map( A1 => shifter_out_7_port, A2 => n1, B1 => 
                           p4_sum_7_port, B2 => n7, C1 => logic_out_7_port, C2 
                           => n4, ZN => n49);
   U38 : INV_X1 port map( A => n50, ZN => OUTALU(6));
   U39 : AOI222_X1 port map( A1 => shifter_out_6_port, A2 => n1, B1 => 
                           p4_sum_6_port, B2 => n7, C1 => logic_out_6_port, C2 
                           => n4, ZN => n50);
   U40 : INV_X1 port map( A => n51, ZN => OUTALU(5));
   U41 : AOI222_X1 port map( A1 => shifter_out_5_port, A2 => n1, B1 => 
                           p4_sum_5_port, B2 => n7, C1 => logic_out_5_port, C2 
                           => n4, ZN => n51);
   U42 : INV_X1 port map( A => n53, ZN => OUTALU(3));
   U43 : AOI222_X1 port map( A1 => shifter_out_3_port, A2 => n1, B1 => 
                           p4_sum_3_port, B2 => n7, C1 => logic_out_3_port, C2 
                           => n4, ZN => n53);
   U44 : INV_X1 port map( A => n56, ZN => OUTALU(2));
   U45 : AOI222_X1 port map( A1 => shifter_out_2_port, A2 => n1, B1 => 
                           p4_sum_2_port, B2 => n7, C1 => logic_out_2_port, C2 
                           => n4, ZN => n56);
   U46 : INV_X1 port map( A => n67, ZN => OUTALU(1));
   U47 : AOI222_X1 port map( A1 => shifter_out_1_port, A2 => n2, B1 => 
                           p4_sum_1_port, B2 => n8, C1 => logic_out_1_port, C2 
                           => n5, ZN => n67);
   U48 : INV_X1 port map( A => n70, ZN => OUTALU(17));
   U49 : AOI222_X1 port map( A1 => shifter_out_17_port, A2 => n3, B1 => 
                           p4_sum_17_port, B2 => n9, C1 => logic_out_17_port, 
                           C2 => n6, ZN => n70);
   U50 : BUF_X1 port map( A => N78, Z => n1);
   U51 : BUF_X1 port map( A => N78, Z => n2);
   U52 : BUF_X1 port map( A => N78, Z => n3);
   U53 : INV_X1 port map( A => n93, ZN => n100);
   U54 : OR2_X1 port map( A1 => n9, A2 => N75, ZN => N74);
   U55 : INV_X1 port map( A => n62, ZN => OUTALU(24));
   U56 : AOI222_X1 port map( A1 => shifter_out_24_port, A2 => n2, B1 => 
                           p4_sum_24_port, B2 => n8, C1 => logic_out_24_port, 
                           C2 => n5, ZN => n62);
   U57 : INV_X1 port map( A => n66, ZN => OUTALU(20));
   U58 : AOI222_X1 port map( A1 => shifter_out_20_port, A2 => n2, B1 => 
                           p4_sum_20_port, B2 => n8, C1 => logic_out_20_port, 
                           C2 => n5, ZN => n66);
   U59 : INV_X1 port map( A => n71, ZN => OUTALU(16));
   U60 : AOI222_X1 port map( A1 => shifter_out_16_port, A2 => n3, B1 => 
                           p4_sum_16_port, B2 => n9, C1 => logic_out_16_port, 
                           C2 => n6, ZN => n71);
   U61 : INV_X1 port map( A => n75_port, ZN => OUTALU(12));
   U62 : AOI222_X1 port map( A1 => shifter_out_12_port, A2 => n3, B1 => 
                           p4_sum_12_port, B2 => n9, C1 => logic_out_12_port, 
                           C2 => n6, ZN => n75_port);
   U63 : OAI222_X1 port map( A1 => s_lt, A2 => n88, B1 => s_eq, B2 => n90, C1 
                           => s_gt, C2 => n91, ZN => n81);
   U64 : AOI22_X1 port map( A1 => n92, A2 => s_gt, B1 => n93, B2 => s_lt, ZN =>
                           n90);
   U65 : BUF_X1 port map( A => DATA1(31), Z => n10);
   U66 : OAI21_X1 port map( B1 => n42, B2 => n84, A => n85, ZN => n83);
   U67 : OAI21_X1 port map( B1 => s_eq, B2 => n86, A => n87, ZN => n85);
   U68 : AOI22_X1 port map( A1 => s_lt, A2 => n103, B1 => s_gt, B2 => n102, ZN 
                           => n84);
   U69 : OAI22_X1 port map( A1 => n100, A2 => s_lt, B1 => n101, B2 => s_gt, ZN 
                           => n87);
   U70 : AOI22_X1 port map( A1 => logic_out_0_port, A2 => n4, B1 => 
                           shifter_out_0_port, B2 => n1, ZN => n78_port);
   U71 : AOI22_X1 port map( A1 => s_eq, A2 => n95, B1 => p4_sum_0_port, B2 => 
                           n7, ZN => n79);
   U72 : AOI221_X1 port map( B1 => n42, B2 => n81, C1 => n82, C2 => s_neq, A =>
                           n83, ZN => n80);
   U73 : INV_X1 port map( A => n58, ZN => OUTALU(28));
   U74 : AOI222_X1 port map( A1 => shifter_out_28_port, A2 => n1, B1 => 
                           p4_sum_28_port, B2 => n7, C1 => logic_out_28_port, 
                           C2 => n4, ZN => n58);
   U75 : INV_X1 port map( A => n48, ZN => OUTALU(8));
   U76 : AOI222_X1 port map( A1 => shifter_out_8_port, A2 => n1, B1 => 
                           p4_sum_8_port, B2 => n7, C1 => logic_out_8_port, C2 
                           => n4, ZN => n48);
   U77 : INV_X1 port map( A => n52, ZN => OUTALU(4));
   U78 : AOI222_X1 port map( A1 => shifter_out_4_port, A2 => n1, B1 => 
                           p4_sum_4_port, B2 => n7, C1 => logic_out_4_port, C2 
                           => n4, ZN => n52);
   U79 : INV_X1 port map( A => n86, ZN => n42);
   U80 : BUF_X1 port map( A => N76, Z => n7);
   U81 : BUF_X1 port map( A => N76, Z => n8);
   U82 : NOR3_X1 port map( A1 => n107, A2 => n106, A3 => n89, ZN => n93);
   U83 : BUF_X1 port map( A => N77, Z => n6);
   U84 : BUF_X1 port map( A => N76, Z => n9);
   U85 : BUF_X1 port map( A => N77, Z => n4);
   U86 : BUF_X1 port map( A => N77, Z => n5);
   U87 : OAI21_X1 port map( B1 => n107, B2 => n46, A => n44, ZN => N78);
   U88 : NOR2_X1 port map( A1 => n45, A2 => n89, ZN => n82);
   U89 : INV_X1 port map( A => n91, ZN => n102);
   U90 : INV_X1 port map( A => n88, ZN => n103);
   U91 : INV_X1 port map( A => n92, ZN => n101);
   U92 : INV_X1 port map( A => n45, ZN => n105);
   U93 : NOR3_X1 port map( A1 => n46, A2 => n106, A3 => n107, ZN => n99);
   U94 : NAND4_X1 port map( A1 => n100, A2 => n88, A3 => n101, A4 => n96, ZN =>
                           N75);
   U95 : AOI211_X1 port map( C1 => n105, C2 => n104, A => n102, B => n95, ZN =>
                           n96);
   U96 : NOR2_X1 port map( A1 => n44, A2 => n43, ZN => n97);
   U97 : NOR2_X1 port map( A1 => n45, A2 => n46, ZN => n98);
   U98 : NAND2_X1 port map( A1 => SN, A2 => n94, ZN => n86);
   U99 : NOR3_X1 port map( A1 => FUNC(0), A2 => FUNC(1), A3 => n89, ZN => n95);
   U100 : NOR3_X1 port map( A1 => n106, A2 => FUNC(0), A3 => n89, ZN => n92);
   U101 : NOR3_X1 port map( A1 => FUNC(2), A2 => FUNC(3), A3 => FUNC(1), ZN => 
                           N76);
   U107 : NAND4_X1 port map( A1 => FUNC(3), A2 => FUNC(2), A3 => n107, A4 => 
                           n106, ZN => n91);
   U108 : INV_X1 port map( A => FUNC(1), ZN => n106);
   U109 : NAND2_X1 port map( A1 => FUNC(2), A2 => n43, ZN => n46);
   U110 : NAND2_X1 port map( A1 => FUNC(3), A2 => n104, ZN => n89);
   U111 : NAND2_X1 port map( A1 => FUNC(0), A2 => n106, ZN => n45);
   U112 : INV_X1 port map( A => FUNC(0), ZN => n107);
   U113 : INV_X1 port map( A => FUNC(2), ZN => n104);
   U114 : INV_X1 port map( A => FUNC(3), ZN => n43);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_0 is

   port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  Y :
         out std_logic);

end MUX41_0;

architecture SYN_BEHAVIORAL_1 of MUX41_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X4
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n1, n2 : std_logic;

begin
   
   U8 : NAND3_X1 port map( A1 => n1, A2 => n2, A3 => A, ZN => n6);
   U1 : OAI211_X4 port map( C1 => n3, C2 => n4, A => n5, B => n6, ZN => Y);
   U2 : NOR2_X1 port map( A1 => S(0), A2 => n2, ZN => n7);
   U3 : NOR2_X1 port map( A1 => n1, A2 => S(1), ZN => n3);
   U4 : NAND2_X1 port map( A1 => B, A2 => n3, ZN => n5);
   U5 : AOI22_X1 port map( A1 => D, A2 => S(0), B1 => n7, B2 => C, ZN => n4);
   U6 : INV_X1 port map( A => S(0), ZN => n1);
   U7 : INV_X1 port map( A => S(1), ZN => n2);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity sum_generator_n_bit32_n_CSB8_0 is

   port( A, B : in std_logic_vector (31 downto 0);  C_in : in std_logic_vector 
         (7 downto 0);  S : out std_logic_vector (31 downto 0));

end sum_generator_n_bit32_n_CSB8_0;

architecture SYN_STRUCTURAL of sum_generator_n_bit32_n_CSB8_0 is

   component carry_select_block_n4_57
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_n4_58
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_n4_59
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_n4_60
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_n4_61
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_n4_62
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_n4_63
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_block_n4_0
      port( A, B : in std_logic_vector (3 downto 0);  C_sel : in std_logic;  S 
            : out std_logic_vector (3 downto 0));
   end component;

begin
   
   csb_0 : carry_select_block_n4_0 port map( A(3) => A(3), A(2) => A(2), A(1) 
                           => A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), 
                           B(1) => B(1), B(0) => B(0), C_sel => C_in(0), S(3) 
                           => S(3), S(2) => S(2), S(1) => S(1), S(0) => S(0));
   csb_1 : carry_select_block_n4_63 port map( A(3) => A(7), A(2) => A(6), A(1) 
                           => A(5), A(0) => A(4), B(3) => B(7), B(2) => B(6), 
                           B(1) => B(5), B(0) => B(4), C_sel => C_in(1), S(3) 
                           => S(7), S(2) => S(6), S(1) => S(5), S(0) => S(4));
   csb_2 : carry_select_block_n4_62 port map( A(3) => A(11), A(2) => A(10), 
                           A(1) => A(9), A(0) => A(8), B(3) => B(11), B(2) => 
                           B(10), B(1) => B(9), B(0) => B(8), C_sel => C_in(2),
                           S(3) => S(11), S(2) => S(10), S(1) => S(9), S(0) => 
                           S(8));
   csb_3 : carry_select_block_n4_61 port map( A(3) => A(15), A(2) => A(14), 
                           A(1) => A(13), A(0) => A(12), B(3) => B(15), B(2) =>
                           B(14), B(1) => B(13), B(0) => B(12), C_sel => 
                           C_in(3), S(3) => S(15), S(2) => S(14), S(1) => S(13)
                           , S(0) => S(12));
   csb_4 : carry_select_block_n4_60 port map( A(3) => A(19), A(2) => A(18), 
                           A(1) => A(17), A(0) => A(16), B(3) => B(19), B(2) =>
                           B(18), B(1) => B(17), B(0) => B(16), C_sel => 
                           C_in(4), S(3) => S(19), S(2) => S(18), S(1) => S(17)
                           , S(0) => S(16));
   csb_5 : carry_select_block_n4_59 port map( A(3) => A(23), A(2) => A(22), 
                           A(1) => A(21), A(0) => A(20), B(3) => B(23), B(2) =>
                           B(22), B(1) => B(21), B(0) => B(20), C_sel => 
                           C_in(5), S(3) => S(23), S(2) => S(22), S(1) => S(21)
                           , S(0) => S(20));
   csb_6 : carry_select_block_n4_58 port map( A(3) => A(27), A(2) => A(26), 
                           A(1) => A(25), A(0) => A(24), B(3) => B(27), B(2) =>
                           B(26), B(1) => B(25), B(0) => B(24), C_sel => 
                           C_in(6), S(3) => S(27), S(2) => S(26), S(1) => S(25)
                           , S(0) => S(24));
   csb_7 : carry_select_block_n4_57 port map( A(3) => A(31), A(2) => A(30), 
                           A(1) => A(29), A(0) => A(28), B(3) => B(31), B(2) =>
                           B(30), B(1) => B(29), B(0) => B(28), C_sel => 
                           C_in(7), S(3) => S(31), S(2) => S(30), S(1) => S(29)
                           , S(0) => S(28));

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_0 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co : 
         out std_logic_vector (7 downto 0));

end CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_0;

architecture SYN_structural of CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component G_BLOCK_61
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component G_BLOCK_62
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component G_BLOCK_63
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component G_BLOCK_64
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component G_BLOCK_65
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component G_BLOCK_66
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component PG_BLOCK_217
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_218
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component G_BLOCK_67
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component PG_BLOCK_219
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_220
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_221
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component G_BLOCK_68
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component PG_BLOCK_222
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_223
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_224
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_225
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_226
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_227
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_228
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component G_BLOCK_0
      port( p2, g2, g1 : in std_logic;  G : out std_logic);
   end component;
   
   component PG_BLOCK_229
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_230
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_231
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_232
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_233
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_234
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_235
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_236
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_237
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_238
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_239
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_240
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_241
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_242
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component PG_BLOCK_0
      port( p2, g2, p1, g1 : in std_logic;  PG_P, PG_G : out std_logic);
   end component;
   
   component pg_net_221
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_222
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_223
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_224
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_225
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_226
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_227
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_228
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_229
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_230
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_231
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_232
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_233
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_234
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_235
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_236
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_237
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_238
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_239
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_240
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_241
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_242
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_243
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_244
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_245
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_246
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_247
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_248
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_249
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_250
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   component pg_net_0
      port( a, b : in std_logic;  p, g : out std_logic);
   end component;
   
   signal Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, Co_2_port, 
      Co_1_port, Co_0_port, g_vector_4_31_port, g_vector_4_27_port, 
      g_vector_3_31_port, g_vector_3_23_port, g_vector_3_15_port, 
      g_vector_2_31_port, g_vector_2_27_port, g_vector_2_23_port, 
      g_vector_2_19_port, g_vector_2_15_port, g_vector_2_11_port, 
      g_vector_2_7_port, g_vector_1_31_port, g_vector_1_29_port, 
      g_vector_1_27_port, g_vector_1_25_port, g_vector_1_23_port, 
      g_vector_1_21_port, g_vector_1_19_port, g_vector_1_17_port, 
      g_vector_1_15_port, g_vector_1_13_port, g_vector_1_11_port, 
      g_vector_1_9_port, g_vector_1_7_port, g_vector_1_5_port, 
      g_vector_1_3_port, g_vector_1_1_port, g_vector_0_31_port, 
      g_vector_0_30_port, g_vector_0_29_port, g_vector_0_28_port, 
      g_vector_0_27_port, g_vector_0_26_port, g_vector_0_25_port, 
      g_vector_0_24_port, g_vector_0_23_port, g_vector_0_22_port, 
      g_vector_0_21_port, g_vector_0_20_port, g_vector_0_19_port, 
      g_vector_0_18_port, g_vector_0_17_port, g_vector_0_16_port, 
      g_vector_0_15_port, g_vector_0_14_port, g_vector_0_13_port, 
      g_vector_0_12_port, g_vector_0_11_port, g_vector_0_10_port, 
      g_vector_0_9_port, g_vector_0_8_port, g_vector_0_7_port, 
      g_vector_0_6_port, g_vector_0_5_port, g_vector_0_4_port, 
      g_vector_0_3_port, g_vector_0_2_port, g_vector_0_1_port, 
      g_vector_0_0_port, p_vector_4_31_port, p_vector_4_27_port, 
      p_vector_3_31_port, p_vector_3_23_port, p_vector_3_15_port, 
      p_vector_2_31_port, p_vector_2_27_port, p_vector_2_23_port, 
      p_vector_2_19_port, p_vector_2_15_port, p_vector_2_11_port, 
      p_vector_2_7_port, p_vector_1_31_port, p_vector_1_29_port, 
      p_vector_1_27_port, p_vector_1_25_port, p_vector_1_23_port, 
      p_vector_1_21_port, p_vector_1_19_port, p_vector_1_17_port, 
      p_vector_1_15_port, p_vector_1_13_port, p_vector_1_11_port, 
      p_vector_1_9_port, p_vector_1_7_port, p_vector_1_5_port, 
      p_vector_1_3_port, p_vector_0_31_port, p_vector_0_30_port, 
      p_vector_0_29_port, p_vector_0_28_port, p_vector_0_27_port, 
      p_vector_0_26_port, p_vector_0_25_port, p_vector_0_24_port, 
      p_vector_0_23_port, p_vector_0_22_port, p_vector_0_21_port, 
      p_vector_0_20_port, p_vector_0_19_port, p_vector_0_18_port, 
      p_vector_0_17_port, p_vector_0_16_port, p_vector_0_15_port, 
      p_vector_0_14_port, p_vector_0_13_port, p_vector_0_12_port, 
      p_vector_0_11_port, p_vector_0_10_port, p_vector_0_9_port, 
      p_vector_0_8_port, p_vector_0_7_port, p_vector_0_6_port, 
      p_vector_0_5_port, p_vector_0_4_port, p_vector_0_3_port, 
      p_vector_0_2_port, p_vector_0_1_port, n3, n1, n2 : std_logic;

begin
   Co <= ( Co_7_port, Co_6_port, Co_5_port, Co_4_port, Co_3_port, Co_2_port, 
      Co_1_port, Co_0_port );
   
   pg_network_31 : pg_net_0 port map( a => A(31), b => B(31), p => 
                           p_vector_0_31_port, g => g_vector_0_31_port);
   pg_network_30 : pg_net_250 port map( a => A(30), b => B(30), p => 
                           p_vector_0_30_port, g => g_vector_0_30_port);
   pg_network_29 : pg_net_249 port map( a => A(29), b => B(29), p => 
                           p_vector_0_29_port, g => g_vector_0_29_port);
   pg_network_28 : pg_net_248 port map( a => A(28), b => B(28), p => 
                           p_vector_0_28_port, g => g_vector_0_28_port);
   pg_network_27 : pg_net_247 port map( a => A(27), b => B(27), p => 
                           p_vector_0_27_port, g => g_vector_0_27_port);
   pg_network_26 : pg_net_246 port map( a => A(26), b => B(26), p => 
                           p_vector_0_26_port, g => g_vector_0_26_port);
   pg_network_25 : pg_net_245 port map( a => A(25), b => B(25), p => 
                           p_vector_0_25_port, g => g_vector_0_25_port);
   pg_network_24 : pg_net_244 port map( a => A(24), b => B(24), p => 
                           p_vector_0_24_port, g => g_vector_0_24_port);
   pg_network_23 : pg_net_243 port map( a => A(23), b => B(23), p => 
                           p_vector_0_23_port, g => g_vector_0_23_port);
   pg_network_22 : pg_net_242 port map( a => A(22), b => B(22), p => 
                           p_vector_0_22_port, g => g_vector_0_22_port);
   pg_network_21 : pg_net_241 port map( a => A(21), b => B(21), p => 
                           p_vector_0_21_port, g => g_vector_0_21_port);
   pg_network_20 : pg_net_240 port map( a => A(20), b => B(20), p => 
                           p_vector_0_20_port, g => g_vector_0_20_port);
   pg_network_19 : pg_net_239 port map( a => A(19), b => B(19), p => 
                           p_vector_0_19_port, g => g_vector_0_19_port);
   pg_network_18 : pg_net_238 port map( a => A(18), b => B(18), p => 
                           p_vector_0_18_port, g => g_vector_0_18_port);
   pg_network_17 : pg_net_237 port map( a => A(17), b => B(17), p => 
                           p_vector_0_17_port, g => g_vector_0_17_port);
   pg_network_16 : pg_net_236 port map( a => A(16), b => B(16), p => 
                           p_vector_0_16_port, g => g_vector_0_16_port);
   pg_network_15 : pg_net_235 port map( a => A(15), b => B(15), p => 
                           p_vector_0_15_port, g => g_vector_0_15_port);
   pg_network_14 : pg_net_234 port map( a => A(14), b => B(14), p => 
                           p_vector_0_14_port, g => g_vector_0_14_port);
   pg_network_13 : pg_net_233 port map( a => A(13), b => B(13), p => 
                           p_vector_0_13_port, g => g_vector_0_13_port);
   pg_network_12 : pg_net_232 port map( a => A(12), b => B(12), p => 
                           p_vector_0_12_port, g => g_vector_0_12_port);
   pg_network_11 : pg_net_231 port map( a => A(11), b => B(11), p => 
                           p_vector_0_11_port, g => g_vector_0_11_port);
   pg_network_10 : pg_net_230 port map( a => A(10), b => B(10), p => 
                           p_vector_0_10_port, g => g_vector_0_10_port);
   pg_network_9 : pg_net_229 port map( a => A(9), b => B(9), p => 
                           p_vector_0_9_port, g => g_vector_0_9_port);
   pg_network_8 : pg_net_228 port map( a => A(8), b => B(8), p => 
                           p_vector_0_8_port, g => g_vector_0_8_port);
   pg_network_7 : pg_net_227 port map( a => A(7), b => B(7), p => 
                           p_vector_0_7_port, g => g_vector_0_7_port);
   pg_network_6 : pg_net_226 port map( a => A(6), b => B(6), p => 
                           p_vector_0_6_port, g => g_vector_0_6_port);
   pg_network_5 : pg_net_225 port map( a => A(5), b => B(5), p => 
                           p_vector_0_5_port, g => g_vector_0_5_port);
   pg_network_4 : pg_net_224 port map( a => A(4), b => B(4), p => 
                           p_vector_0_4_port, g => g_vector_0_4_port);
   pg_network_3 : pg_net_223 port map( a => A(3), b => B(3), p => 
                           p_vector_0_3_port, g => g_vector_0_3_port);
   pg_network_2 : pg_net_222 port map( a => A(2), b => B(2), p => 
                           p_vector_0_2_port, g => g_vector_0_2_port);
   pg_network_1 : pg_net_221 port map( a => A(1), b => B(1), p => 
                           p_vector_0_1_port, g => g_vector_0_1_port);
   std_PG_1_31 : PG_BLOCK_0 port map( p2 => p_vector_0_31_port, g2 => 
                           g_vector_0_31_port, p1 => p_vector_0_30_port, g1 => 
                           g_vector_0_30_port, PG_P => p_vector_1_31_port, PG_G
                           => g_vector_1_31_port);
   std_PG_1_29 : PG_BLOCK_242 port map( p2 => p_vector_0_29_port, g2 => 
                           g_vector_0_29_port, p1 => p_vector_0_28_port, g1 => 
                           g_vector_0_28_port, PG_P => p_vector_1_29_port, PG_G
                           => g_vector_1_29_port);
   std_PG_1_27 : PG_BLOCK_241 port map( p2 => p_vector_0_27_port, g2 => 
                           g_vector_0_27_port, p1 => p_vector_0_26_port, g1 => 
                           g_vector_0_26_port, PG_P => p_vector_1_27_port, PG_G
                           => g_vector_1_27_port);
   std_PG_1_25 : PG_BLOCK_240 port map( p2 => p_vector_0_25_port, g2 => 
                           g_vector_0_25_port, p1 => p_vector_0_24_port, g1 => 
                           g_vector_0_24_port, PG_P => p_vector_1_25_port, PG_G
                           => g_vector_1_25_port);
   std_PG_1_23 : PG_BLOCK_239 port map( p2 => p_vector_0_23_port, g2 => 
                           g_vector_0_23_port, p1 => p_vector_0_22_port, g1 => 
                           g_vector_0_22_port, PG_P => p_vector_1_23_port, PG_G
                           => g_vector_1_23_port);
   std_PG_1_21 : PG_BLOCK_238 port map( p2 => p_vector_0_21_port, g2 => 
                           g_vector_0_21_port, p1 => p_vector_0_20_port, g1 => 
                           g_vector_0_20_port, PG_P => p_vector_1_21_port, PG_G
                           => g_vector_1_21_port);
   std_PG_1_19 : PG_BLOCK_237 port map( p2 => p_vector_0_19_port, g2 => 
                           g_vector_0_19_port, p1 => p_vector_0_18_port, g1 => 
                           g_vector_0_18_port, PG_P => p_vector_1_19_port, PG_G
                           => g_vector_1_19_port);
   std_PG_1_17 : PG_BLOCK_236 port map( p2 => p_vector_0_17_port, g2 => 
                           g_vector_0_17_port, p1 => p_vector_0_16_port, g1 => 
                           g_vector_0_16_port, PG_P => p_vector_1_17_port, PG_G
                           => g_vector_1_17_port);
   std_PG_1_15 : PG_BLOCK_235 port map( p2 => p_vector_0_15_port, g2 => 
                           g_vector_0_15_port, p1 => p_vector_0_14_port, g1 => 
                           g_vector_0_14_port, PG_P => p_vector_1_15_port, PG_G
                           => g_vector_1_15_port);
   std_PG_1_13 : PG_BLOCK_234 port map( p2 => p_vector_0_13_port, g2 => 
                           g_vector_0_13_port, p1 => p_vector_0_12_port, g1 => 
                           g_vector_0_12_port, PG_P => p_vector_1_13_port, PG_G
                           => g_vector_1_13_port);
   std_PG_1_11 : PG_BLOCK_233 port map( p2 => p_vector_0_11_port, g2 => 
                           g_vector_0_11_port, p1 => p_vector_0_10_port, g1 => 
                           g_vector_0_10_port, PG_P => p_vector_1_11_port, PG_G
                           => g_vector_1_11_port);
   std_PG_1_9 : PG_BLOCK_232 port map( p2 => p_vector_0_9_port, g2 => 
                           g_vector_0_9_port, p1 => p_vector_0_8_port, g1 => 
                           g_vector_0_8_port, PG_P => p_vector_1_9_port, PG_G 
                           => g_vector_1_9_port);
   std_PG_1_7 : PG_BLOCK_231 port map( p2 => p_vector_0_7_port, g2 => 
                           g_vector_0_7_port, p1 => p_vector_0_6_port, g1 => 
                           g_vector_0_6_port, PG_P => p_vector_1_7_port, PG_G 
                           => g_vector_1_7_port);
   std_PG_1_5 : PG_BLOCK_230 port map( p2 => p_vector_0_5_port, g2 => 
                           g_vector_0_5_port, p1 => p_vector_0_4_port, g1 => 
                           g_vector_0_4_port, PG_P => p_vector_1_5_port, PG_G 
                           => g_vector_1_5_port);
   std_PG_1_3 : PG_BLOCK_229 port map( p2 => p_vector_0_3_port, g2 => 
                           g_vector_0_3_port, p1 => p_vector_0_2_port, g1 => 
                           g_vector_0_2_port, PG_P => p_vector_1_3_port, PG_G 
                           => g_vector_1_3_port);
   std_G_1_1 : G_BLOCK_0 port map( p2 => p_vector_0_1_port, g2 => 
                           g_vector_0_1_port, g1 => g_vector_0_0_port, G => 
                           g_vector_1_1_port);
   std_PG_2_31 : PG_BLOCK_228 port map( p2 => p_vector_1_31_port, g2 => 
                           g_vector_1_31_port, p1 => p_vector_1_29_port, g1 => 
                           g_vector_1_29_port, PG_P => p_vector_2_31_port, PG_G
                           => g_vector_2_31_port);
   std_PG_2_27 : PG_BLOCK_227 port map( p2 => p_vector_1_27_port, g2 => 
                           g_vector_1_27_port, p1 => p_vector_1_25_port, g1 => 
                           g_vector_1_25_port, PG_P => p_vector_2_27_port, PG_G
                           => g_vector_2_27_port);
   std_PG_2_23 : PG_BLOCK_226 port map( p2 => p_vector_1_23_port, g2 => 
                           g_vector_1_23_port, p1 => p_vector_1_21_port, g1 => 
                           g_vector_1_21_port, PG_P => p_vector_2_23_port, PG_G
                           => g_vector_2_23_port);
   std_PG_2_19 : PG_BLOCK_225 port map( p2 => p_vector_1_19_port, g2 => 
                           g_vector_1_19_port, p1 => p_vector_1_17_port, g1 => 
                           g_vector_1_17_port, PG_P => p_vector_2_19_port, PG_G
                           => g_vector_2_19_port);
   std_PG_2_15 : PG_BLOCK_224 port map( p2 => p_vector_1_15_port, g2 => 
                           g_vector_1_15_port, p1 => p_vector_1_13_port, g1 => 
                           g_vector_1_13_port, PG_P => p_vector_2_15_port, PG_G
                           => g_vector_2_15_port);
   std_PG_2_11 : PG_BLOCK_223 port map( p2 => p_vector_1_11_port, g2 => 
                           g_vector_1_11_port, p1 => p_vector_1_9_port, g1 => 
                           g_vector_1_9_port, PG_P => p_vector_2_11_port, PG_G 
                           => g_vector_2_11_port);
   std_PG_2_7 : PG_BLOCK_222 port map( p2 => p_vector_1_7_port, g2 => 
                           g_vector_1_7_port, p1 => p_vector_1_5_port, g1 => 
                           g_vector_1_5_port, PG_P => p_vector_2_7_port, PG_G 
                           => g_vector_2_7_port);
   std_G_2_3 : G_BLOCK_68 port map( p2 => p_vector_1_3_port, g2 => 
                           g_vector_1_3_port, g1 => g_vector_1_1_port, G => 
                           Co_0_port);
   std_PG_3_31 : PG_BLOCK_221 port map( p2 => p_vector_2_31_port, g2 => 
                           g_vector_2_31_port, p1 => p_vector_2_27_port, g1 => 
                           g_vector_2_27_port, PG_P => p_vector_3_31_port, PG_G
                           => g_vector_3_31_port);
   std_PG_3_23 : PG_BLOCK_220 port map( p2 => p_vector_2_23_port, g2 => 
                           g_vector_2_23_port, p1 => p_vector_2_19_port, g1 => 
                           g_vector_2_19_port, PG_P => p_vector_3_23_port, PG_G
                           => g_vector_3_23_port);
   std_PG_3_15 : PG_BLOCK_219 port map( p2 => p_vector_2_15_port, g2 => 
                           g_vector_2_15_port, p1 => p_vector_2_11_port, g1 => 
                           g_vector_2_11_port, PG_P => p_vector_3_15_port, PG_G
                           => g_vector_3_15_port);
   std_G_3_7 : G_BLOCK_67 port map( p2 => p_vector_2_7_port, g2 => 
                           g_vector_2_7_port, g1 => Co_0_port, G => Co_1_port);
   std_PG_4_31 : PG_BLOCK_218 port map( p2 => p_vector_3_31_port, g2 => 
                           g_vector_3_31_port, p1 => p_vector_3_23_port, g1 => 
                           g_vector_3_23_port, PG_P => p_vector_4_31_port, PG_G
                           => g_vector_4_31_port);
   add_PG_4_31_1 : PG_BLOCK_217 port map( p2 => p_vector_2_27_port, g2 => 
                           g_vector_2_27_port, p1 => p_vector_3_23_port, g1 => 
                           g_vector_3_23_port, PG_P => p_vector_4_27_port, PG_G
                           => g_vector_4_27_port);
   std_G_4_15 : G_BLOCK_66 port map( p2 => p_vector_3_15_port, g2 => 
                           g_vector_3_15_port, g1 => Co_1_port, G => Co_3_port)
                           ;
   add_G_4_15_1 : G_BLOCK_65 port map( p2 => p_vector_2_11_port, g2 => 
                           g_vector_2_11_port, g1 => Co_1_port, G => Co_2_port)
                           ;
   std_G_5_31 : G_BLOCK_64 port map( p2 => p_vector_4_31_port, g2 => 
                           g_vector_4_31_port, g1 => Co_3_port, G => Co_7_port)
                           ;
   add_G_5_31_1 : G_BLOCK_63 port map( p2 => p_vector_4_27_port, g2 => 
                           g_vector_4_27_port, g1 => Co_3_port, G => Co_6_port)
                           ;
   add_G_5_31_2 : G_BLOCK_62 port map( p2 => p_vector_3_23_port, g2 => 
                           g_vector_3_23_port, g1 => Co_3_port, G => Co_5_port)
                           ;
   add_G_5_31_3 : G_BLOCK_61 port map( p2 => p_vector_2_19_port, g2 => 
                           g_vector_2_19_port, g1 => Co_3_port, G => Co_4_port)
                           ;
   U1 : INV_X1 port map( A => B(0), ZN => n2);
   U2 : OAI21_X1 port map( B1 => n1, B2 => n2, A => n3, ZN => g_vector_0_0_port
                           );
   U3 : OAI21_X1 port map( B1 => A(0), B2 => B(0), A => Cin, ZN => n3);
   U4 : INV_X1 port map( A => A(0), ZN => n1);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity my_xor_0 is

   port( A, B : in std_logic;  xor_out : out std_logic);

end my_xor_0;

architecture SYN_behavioral of my_xor_0 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => xor_out);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX51_GENERIC_NBIT32 is

   port( A, B, C, D, E : in std_logic_vector (31 downto 0);  SEL : in 
         std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end MUX51_GENERIC_NBIT32;

architecture SYN_structural of MUX51_GENERIC_NBIT32 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX51_1
      port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0)
            ;  Y : out std_logic);
   end component;
   
   component MUX51_2
      port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0)
            ;  Y : out std_logic);
   end component;
   
   component MUX51_3
      port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0)
            ;  Y : out std_logic);
   end component;
   
   component MUX51_4
      port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0)
            ;  Y : out std_logic);
   end component;
   
   component MUX51_5
      port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0)
            ;  Y : out std_logic);
   end component;
   
   component MUX51_6
      port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0)
            ;  Y : out std_logic);
   end component;
   
   component MUX51_7
      port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0)
            ;  Y : out std_logic);
   end component;
   
   component MUX51_8
      port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0)
            ;  Y : out std_logic);
   end component;
   
   component MUX51_9
      port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0)
            ;  Y : out std_logic);
   end component;
   
   component MUX51_10
      port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0)
            ;  Y : out std_logic);
   end component;
   
   component MUX51_11
      port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0)
            ;  Y : out std_logic);
   end component;
   
   component MUX51_12
      port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0)
            ;  Y : out std_logic);
   end component;
   
   component MUX51_13
      port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0)
            ;  Y : out std_logic);
   end component;
   
   component MUX51_14
      port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0)
            ;  Y : out std_logic);
   end component;
   
   component MUX51_15
      port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0)
            ;  Y : out std_logic);
   end component;
   
   component MUX51_16
      port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0)
            ;  Y : out std_logic);
   end component;
   
   component MUX51_17
      port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0)
            ;  Y : out std_logic);
   end component;
   
   component MUX51_18
      port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0)
            ;  Y : out std_logic);
   end component;
   
   component MUX51_19
      port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0)
            ;  Y : out std_logic);
   end component;
   
   component MUX51_20
      port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0)
            ;  Y : out std_logic);
   end component;
   
   component MUX51_21
      port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0)
            ;  Y : out std_logic);
   end component;
   
   component MUX51_22
      port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0)
            ;  Y : out std_logic);
   end component;
   
   component MUX51_23
      port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0)
            ;  Y : out std_logic);
   end component;
   
   component MUX51_24
      port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0)
            ;  Y : out std_logic);
   end component;
   
   component MUX51_25
      port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0)
            ;  Y : out std_logic);
   end component;
   
   component MUX51_26
      port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0)
            ;  Y : out std_logic);
   end component;
   
   component MUX51_27
      port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0)
            ;  Y : out std_logic);
   end component;
   
   component MUX51_28
      port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0)
            ;  Y : out std_logic);
   end component;
   
   component MUX51_29
      port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0)
            ;  Y : out std_logic);
   end component;
   
   component MUX51_30
      port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0)
            ;  Y : out std_logic);
   end component;
   
   component MUX51_31
      port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0)
            ;  Y : out std_logic);
   end component;
   
   component MUX51_0
      port( A, B, C, D, E : in std_logic;  S : in std_logic_vector (2 downto 0)
            ;  Y : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9 : std_logic;

begin
   
   MUXES_0 : MUX51_0 port map( A => A(0), B => B(0), C => C(0), D => D(0), E =>
                           E(0), S(2) => n9, S(1) => n6, S(0) => n3, Y => Y(0))
                           ;
   MUXES_1 : MUX51_31 port map( A => A(1), B => B(1), C => C(1), D => D(1), E 
                           => E(1), S(2) => n7, S(1) => n4, S(0) => n1, Y => 
                           Y(1));
   MUXES_2 : MUX51_30 port map( A => A(2), B => B(2), C => C(2), D => D(2), E 
                           => E(2), S(2) => n7, S(1) => n4, S(0) => n1, Y => 
                           Y(2));
   MUXES_3 : MUX51_29 port map( A => A(3), B => B(3), C => C(3), D => D(3), E 
                           => E(3), S(2) => n7, S(1) => n4, S(0) => n1, Y => 
                           Y(3));
   MUXES_4 : MUX51_28 port map( A => A(4), B => B(4), C => C(4), D => D(4), E 
                           => E(4), S(2) => n7, S(1) => n4, S(0) => n1, Y => 
                           Y(4));
   MUXES_5 : MUX51_27 port map( A => A(5), B => B(5), C => C(5), D => D(5), E 
                           => E(5), S(2) => n7, S(1) => n4, S(0) => n1, Y => 
                           Y(5));
   MUXES_6 : MUX51_26 port map( A => A(6), B => B(6), C => C(6), D => D(6), E 
                           => E(6), S(2) => n7, S(1) => n4, S(0) => n1, Y => 
                           Y(6));
   MUXES_7 : MUX51_25 port map( A => A(7), B => B(7), C => C(7), D => D(7), E 
                           => E(7), S(2) => n7, S(1) => n4, S(0) => n1, Y => 
                           Y(7));
   MUXES_8 : MUX51_24 port map( A => A(8), B => B(8), C => C(8), D => D(8), E 
                           => E(8), S(2) => n7, S(1) => n4, S(0) => n1, Y => 
                           Y(8));
   MUXES_9 : MUX51_23 port map( A => A(9), B => B(9), C => C(9), D => D(9), E 
                           => E(9), S(2) => n7, S(1) => n4, S(0) => n1, Y => 
                           Y(9));
   MUXES_10 : MUX51_22 port map( A => A(10), B => B(10), C => C(10), D => D(10)
                           , E => E(10), S(2) => n7, S(1) => n4, S(0) => n1, Y 
                           => Y(10));
   MUXES_11 : MUX51_21 port map( A => A(11), B => B(11), C => C(11), D => D(11)
                           , E => E(11), S(2) => n7, S(1) => n4, S(0) => n1, Y 
                           => Y(11));
   MUXES_12 : MUX51_20 port map( A => A(12), B => B(12), C => C(12), D => D(12)
                           , E => E(12), S(2) => n7, S(1) => n4, S(0) => n1, Y 
                           => Y(12));
   MUXES_13 : MUX51_19 port map( A => A(13), B => B(13), C => C(13), D => D(13)
                           , E => E(13), S(2) => n8, S(1) => n5, S(0) => n2, Y 
                           => Y(13));
   MUXES_14 : MUX51_18 port map( A => A(14), B => B(14), C => C(14), D => D(14)
                           , E => E(14), S(2) => n8, S(1) => n5, S(0) => n2, Y 
                           => Y(14));
   MUXES_15 : MUX51_17 port map( A => A(15), B => B(15), C => C(15), D => D(15)
                           , E => E(15), S(2) => n8, S(1) => n5, S(0) => n2, Y 
                           => Y(15));
   MUXES_16 : MUX51_16 port map( A => A(16), B => B(16), C => C(16), D => D(16)
                           , E => E(16), S(2) => n8, S(1) => n5, S(0) => n2, Y 
                           => Y(16));
   MUXES_17 : MUX51_15 port map( A => A(17), B => B(17), C => C(17), D => D(17)
                           , E => E(17), S(2) => n8, S(1) => n5, S(0) => n2, Y 
                           => Y(17));
   MUXES_18 : MUX51_14 port map( A => A(18), B => B(18), C => C(18), D => D(18)
                           , E => E(18), S(2) => n8, S(1) => n5, S(0) => n2, Y 
                           => Y(18));
   MUXES_19 : MUX51_13 port map( A => A(19), B => B(19), C => C(19), D => D(19)
                           , E => E(19), S(2) => n8, S(1) => n5, S(0) => n2, Y 
                           => Y(19));
   MUXES_20 : MUX51_12 port map( A => A(20), B => B(20), C => C(20), D => D(20)
                           , E => E(20), S(2) => n8, S(1) => n5, S(0) => n2, Y 
                           => Y(20));
   MUXES_21 : MUX51_11 port map( A => A(21), B => B(21), C => C(21), D => D(21)
                           , E => E(21), S(2) => n8, S(1) => n5, S(0) => n2, Y 
                           => Y(21));
   MUXES_22 : MUX51_10 port map( A => A(22), B => B(22), C => C(22), D => D(22)
                           , E => E(22), S(2) => n8, S(1) => n5, S(0) => n2, Y 
                           => Y(22));
   MUXES_23 : MUX51_9 port map( A => A(23), B => B(23), C => C(23), D => D(23),
                           E => E(23), S(2) => n8, S(1) => n5, S(0) => n2, Y =>
                           Y(23));
   MUXES_24 : MUX51_8 port map( A => A(24), B => B(24), C => C(24), D => D(24),
                           E => E(24), S(2) => n8, S(1) => n5, S(0) => n2, Y =>
                           Y(24));
   MUXES_25 : MUX51_7 port map( A => A(25), B => B(25), C => C(25), D => D(25),
                           E => E(25), S(2) => n9, S(1) => n6, S(0) => n3, Y =>
                           Y(25));
   MUXES_26 : MUX51_6 port map( A => A(26), B => B(26), C => C(26), D => D(26),
                           E => E(26), S(2) => n9, S(1) => n6, S(0) => n3, Y =>
                           Y(26));
   MUXES_27 : MUX51_5 port map( A => A(27), B => B(27), C => C(27), D => D(27),
                           E => E(27), S(2) => n9, S(1) => n6, S(0) => n3, Y =>
                           Y(27));
   MUXES_28 : MUX51_4 port map( A => A(28), B => B(28), C => C(28), D => D(28),
                           E => E(28), S(2) => n9, S(1) => n6, S(0) => n3, Y =>
                           Y(28));
   MUXES_29 : MUX51_3 port map( A => A(29), B => B(29), C => C(29), D => D(29),
                           E => E(29), S(2) => n9, S(1) => n6, S(0) => n3, Y =>
                           Y(29));
   MUXES_30 : MUX51_2 port map( A => A(30), B => B(30), C => C(30), D => D(30),
                           E => E(30), S(2) => n9, S(1) => n6, S(0) => n3, Y =>
                           Y(30));
   MUXES_31 : MUX51_1 port map( A => A(31), B => B(31), C => C(31), D => D(31),
                           E => E(31), S(2) => n9, S(1) => n6, S(0) => n3, Y =>
                           Y(31));
   U1 : BUF_X1 port map( A => SEL(0), Z => n3);
   U2 : BUF_X2 port map( A => SEL(0), Z => n2);
   U3 : BUF_X2 port map( A => SEL(0), Z => n1);
   U4 : BUF_X1 port map( A => SEL(1), Z => n5);
   U5 : BUF_X1 port map( A => SEL(1), Z => n4);
   U6 : BUF_X1 port map( A => SEL(2), Z => n8);
   U7 : BUF_X1 port map( A => SEL(2), Z => n7);
   U8 : BUF_X1 port map( A => SEL(1), Z => n6);
   U9 : BUF_X1 port map( A => SEL(2), Z => n9);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MMU_WORD_size32 is

   port( Wrd, BHU0 : in std_logic;  wdata_size : out std_logic_vector (1 downto
         0));

end MMU_WORD_size32;

architecture SYN_Behavioral of MMU_WORD_size32 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal N3 : std_logic;

begin
   wdata_size <= ( Wrd, N3 );
   
   U2 : OR2_X1 port map( A1 => BHU0, A2 => Wrd, ZN => N3);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity EXU_N32 is

   port( DATA1, DATA2 : in std_logic_vector (31 downto 0);  FUNC : in 
         std_logic_vector (3 downto 0);  RD_in : in std_logic_vector (4 downto 
         0);  SN, CLK, RST : in std_logic;  OVF, stall_flag, RD_sel_flag : out 
         std_logic;  OUTPUT : out std_logic_vector (31 downto 0);  RD_stall, 
         RD_out : out std_logic_vector (4 downto 0);  H_MULOUT : out 
         std_logic_vector (31 downto 0));

end EXU_N32;

architecture SYN_structural of EXU_N32 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX21_GENERIC_NBIT32_1
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component boothmul_NBIT_in32
      port( A, B : in std_logic_vector (31 downto 0);  mulin_flag, CLK, RST : 
            in std_logic;  MULready : out std_logic;  P : out std_logic_vector 
            (63 downto 0));
   end component;
   
   component ALU_N32
      port( DATA1, DATA2 : in std_logic_vector (31 downto 0);  FUNC : in 
            std_logic_vector (3 downto 0);  SN : in std_logic;  OVF : out 
            std_logic;  OUTALU : out std_logic_vector (31 downto 0));
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal RD_sel_flag_port, RD_stall_4_port, RD_stall_3_port, RD_stall_2_port, 
      RD_stall_1_port, RD_stall_0_port, RD_reg2_4_port, RD_reg2_3_port, 
      RD_reg2_2_port, RD_reg2_1_port, RD_reg2_0_port, mul_flag_reg1, 
      s_RD_in_4_port, s_RD_in_3_port, s_RD_in_2_port, s_RD_in_1_port, 
      s_RD_in_0_port, N3, s_ALUout_31_port, s_ALUout_30_port, s_ALUout_29_port,
      s_ALUout_28_port, s_ALUout_27_port, s_ALUout_26_port, s_ALUout_25_port, 
      s_ALUout_24_port, s_ALUout_23_port, s_ALUout_22_port, s_ALUout_21_port, 
      s_ALUout_20_port, s_ALUout_19_port, s_ALUout_18_port, s_ALUout_17_port, 
      s_ALUout_16_port, s_ALUout_15_port, s_ALUout_14_port, s_ALUout_13_port, 
      s_ALUout_12_port, s_ALUout_11_port, s_ALUout_10_port, s_ALUout_9_port, 
      s_ALUout_8_port, s_ALUout_7_port, s_ALUout_6_port, s_ALUout_5_port, 
      s_ALUout_4_port, s_ALUout_3_port, s_ALUout_2_port, s_ALUout_1_port, 
      s_ALUout_0_port, s_mul_out_31_port, s_mul_out_30_port, s_mul_out_29_port,
      s_mul_out_28_port, s_mul_out_27_port, s_mul_out_26_port, 
      s_mul_out_25_port, s_mul_out_24_port, s_mul_out_23_port, 
      s_mul_out_22_port, s_mul_out_21_port, s_mul_out_20_port, 
      s_mul_out_19_port, s_mul_out_18_port, s_mul_out_17_port, 
      s_mul_out_16_port, s_mul_out_15_port, s_mul_out_14_port, 
      s_mul_out_13_port, s_mul_out_12_port, s_mul_out_11_port, 
      s_mul_out_10_port, s_mul_out_9_port, s_mul_out_8_port, s_mul_out_7_port, 
      s_mul_out_6_port, s_mul_out_5_port, s_mul_out_4_port, s_mul_out_3_port, 
      s_mul_out_2_port, s_mul_out_1_port, s_mul_out_0_port, n1, n_1922, n_1923,
      n_1924, n_1925, n_1926, n_1927, n_1928, n_1929, n_1930, n_1931, n_1932, 
      n_1933, n_1934, n_1935, n_1936, n_1937, n_1938 : std_logic;

begin
   RD_sel_flag <= RD_sel_flag_port;
   RD_stall <= ( RD_stall_4_port, RD_stall_3_port, RD_stall_2_port, 
      RD_stall_1_port, RD_stall_0_port );
   
   RD_reg1_reg_4_inst : DFFR_X1 port map( D => s_RD_in_4_port, CK => CLK, RN =>
                           n1, Q => RD_stall_4_port, QN => n_1922);
   RD_reg1_reg_3_inst : DFFR_X1 port map( D => s_RD_in_3_port, CK => CLK, RN =>
                           n1, Q => RD_stall_3_port, QN => n_1923);
   RD_reg1_reg_2_inst : DFFR_X1 port map( D => s_RD_in_2_port, CK => CLK, RN =>
                           n1, Q => RD_stall_2_port, QN => n_1924);
   RD_reg1_reg_1_inst : DFFR_X1 port map( D => s_RD_in_1_port, CK => CLK, RN =>
                           n1, Q => RD_stall_1_port, QN => n_1925);
   RD_reg1_reg_0_inst : DFFR_X1 port map( D => s_RD_in_0_port, CK => CLK, RN =>
                           n1, Q => RD_stall_0_port, QN => n_1926);
   RD_reg2_reg_4_inst : DFFR_X1 port map( D => RD_stall_4_port, CK => CLK, RN 
                           => n1, Q => RD_reg2_4_port, QN => n_1927);
   RD_reg2_reg_3_inst : DFFR_X1 port map( D => RD_stall_3_port, CK => CLK, RN 
                           => n1, Q => RD_reg2_3_port, QN => n_1928);
   RD_reg2_reg_2_inst : DFFR_X1 port map( D => RD_stall_2_port, CK => CLK, RN 
                           => n1, Q => RD_reg2_2_port, QN => n_1929);
   RD_reg2_reg_1_inst : DFFR_X1 port map( D => RD_stall_1_port, CK => CLK, RN 
                           => n1, Q => RD_reg2_1_port, QN => n_1930);
   RD_reg2_reg_0_inst : DFFR_X1 port map( D => RD_stall_0_port, CK => CLK, RN 
                           => n1, Q => RD_reg2_0_port, QN => n_1931);
   RD_reg3_reg_4_inst : DFFR_X1 port map( D => RD_reg2_4_port, CK => CLK, RN =>
                           n1, Q => RD_out(4), QN => n_1932);
   RD_reg3_reg_3_inst : DFFR_X1 port map( D => RD_reg2_3_port, CK => CLK, RN =>
                           n1, Q => RD_out(3), QN => n_1933);
   RD_reg3_reg_2_inst : DFFR_X1 port map( D => RD_reg2_2_port, CK => CLK, RN =>
                           n1, Q => RD_out(2), QN => n_1934);
   RD_reg3_reg_1_inst : DFFR_X1 port map( D => RD_reg2_1_port, CK => CLK, RN =>
                           n1, Q => RD_out(1), QN => n_1935);
   RD_reg3_reg_0_inst : DFFR_X1 port map( D => RD_reg2_0_port, CK => CLK, RN =>
                           n1, Q => RD_out(0), QN => n_1936);
   mul_flag_reg1_reg : DFFR_X1 port map( D => N3, CK => CLK, RN => n1, Q => 
                           mul_flag_reg1, QN => n_1937);
   mul_flag_reg2_reg : DFFR_X1 port map( D => mul_flag_reg1, CK => CLK, RN => 
                           n1, Q => stall_flag, QN => n_1938);
   ALU1 : ALU_N32 port map( DATA1(31) => DATA1(31), DATA1(30) => DATA1(30), 
                           DATA1(29) => DATA1(29), DATA1(28) => DATA1(28), 
                           DATA1(27) => DATA1(27), DATA1(26) => DATA1(26), 
                           DATA1(25) => DATA1(25), DATA1(24) => DATA1(24), 
                           DATA1(23) => DATA1(23), DATA1(22) => DATA1(22), 
                           DATA1(21) => DATA1(21), DATA1(20) => DATA1(20), 
                           DATA1(19) => DATA1(19), DATA1(18) => DATA1(18), 
                           DATA1(17) => DATA1(17), DATA1(16) => DATA1(16), 
                           DATA1(15) => DATA1(15), DATA1(14) => DATA1(14), 
                           DATA1(13) => DATA1(13), DATA1(12) => DATA1(12), 
                           DATA1(11) => DATA1(11), DATA1(10) => DATA1(10), 
                           DATA1(9) => DATA1(9), DATA1(8) => DATA1(8), DATA1(7)
                           => DATA1(7), DATA1(6) => DATA1(6), DATA1(5) => 
                           DATA1(5), DATA1(4) => DATA1(4), DATA1(3) => DATA1(3)
                           , DATA1(2) => DATA1(2), DATA1(1) => DATA1(1), 
                           DATA1(0) => DATA1(0), DATA2(31) => DATA2(31), 
                           DATA2(30) => DATA2(30), DATA2(29) => DATA2(29), 
                           DATA2(28) => DATA2(28), DATA2(27) => DATA2(27), 
                           DATA2(26) => DATA2(26), DATA2(25) => DATA2(25), 
                           DATA2(24) => DATA2(24), DATA2(23) => DATA2(23), 
                           DATA2(22) => DATA2(22), DATA2(21) => DATA2(21), 
                           DATA2(20) => DATA2(20), DATA2(19) => DATA2(19), 
                           DATA2(18) => DATA2(18), DATA2(17) => DATA2(17), 
                           DATA2(16) => DATA2(16), DATA2(15) => DATA2(15), 
                           DATA2(14) => DATA2(14), DATA2(13) => DATA2(13), 
                           DATA2(12) => DATA2(12), DATA2(11) => DATA2(11), 
                           DATA2(10) => DATA2(10), DATA2(9) => DATA2(9), 
                           DATA2(8) => DATA2(8), DATA2(7) => DATA2(7), DATA2(6)
                           => DATA2(6), DATA2(5) => DATA2(5), DATA2(4) => 
                           DATA2(4), DATA2(3) => DATA2(3), DATA2(2) => DATA2(2)
                           , DATA2(1) => DATA2(1), DATA2(0) => DATA2(0), 
                           FUNC(3) => FUNC(3), FUNC(2) => FUNC(2), FUNC(1) => 
                           FUNC(1), FUNC(0) => FUNC(0), SN => SN, OVF => OVF, 
                           OUTALU(31) => s_ALUout_31_port, OUTALU(30) => 
                           s_ALUout_30_port, OUTALU(29) => s_ALUout_29_port, 
                           OUTALU(28) => s_ALUout_28_port, OUTALU(27) => 
                           s_ALUout_27_port, OUTALU(26) => s_ALUout_26_port, 
                           OUTALU(25) => s_ALUout_25_port, OUTALU(24) => 
                           s_ALUout_24_port, OUTALU(23) => s_ALUout_23_port, 
                           OUTALU(22) => s_ALUout_22_port, OUTALU(21) => 
                           s_ALUout_21_port, OUTALU(20) => s_ALUout_20_port, 
                           OUTALU(19) => s_ALUout_19_port, OUTALU(18) => 
                           s_ALUout_18_port, OUTALU(17) => s_ALUout_17_port, 
                           OUTALU(16) => s_ALUout_16_port, OUTALU(15) => 
                           s_ALUout_15_port, OUTALU(14) => s_ALUout_14_port, 
                           OUTALU(13) => s_ALUout_13_port, OUTALU(12) => 
                           s_ALUout_12_port, OUTALU(11) => s_ALUout_11_port, 
                           OUTALU(10) => s_ALUout_10_port, OUTALU(9) => 
                           s_ALUout_9_port, OUTALU(8) => s_ALUout_8_port, 
                           OUTALU(7) => s_ALUout_7_port, OUTALU(6) => 
                           s_ALUout_6_port, OUTALU(5) => s_ALUout_5_port, 
                           OUTALU(4) => s_ALUout_4_port, OUTALU(3) => 
                           s_ALUout_3_port, OUTALU(2) => s_ALUout_2_port, 
                           OUTALU(1) => s_ALUout_1_port, OUTALU(0) => 
                           s_ALUout_0_port);
   MUL : boothmul_NBIT_in32 port map( A(31) => DATA1(31), A(30) => DATA1(30), 
                           A(29) => DATA1(29), A(28) => DATA1(28), A(27) => 
                           DATA1(27), A(26) => DATA1(26), A(25) => DATA1(25), 
                           A(24) => DATA1(24), A(23) => DATA1(23), A(22) => 
                           DATA1(22), A(21) => DATA1(21), A(20) => DATA1(20), 
                           A(19) => DATA1(19), A(18) => DATA1(18), A(17) => 
                           DATA1(17), A(16) => DATA1(16), A(15) => DATA1(15), 
                           A(14) => DATA1(14), A(13) => DATA1(13), A(12) => 
                           DATA1(12), A(11) => DATA1(11), A(10) => DATA1(10), 
                           A(9) => DATA1(9), A(8) => DATA1(8), A(7) => DATA1(7)
                           , A(6) => DATA1(6), A(5) => DATA1(5), A(4) => 
                           DATA1(4), A(3) => DATA1(3), A(2) => DATA1(2), A(1) 
                           => DATA1(1), A(0) => DATA1(0), B(31) => DATA2(31), 
                           B(30) => DATA2(30), B(29) => DATA2(29), B(28) => 
                           DATA2(28), B(27) => DATA2(27), B(26) => DATA2(26), 
                           B(25) => DATA2(25), B(24) => DATA2(24), B(23) => 
                           DATA2(23), B(22) => DATA2(22), B(21) => DATA2(21), 
                           B(20) => DATA2(20), B(19) => DATA2(19), B(18) => 
                           DATA2(18), B(17) => DATA2(17), B(16) => DATA2(16), 
                           B(15) => DATA2(15), B(14) => DATA2(14), B(13) => 
                           DATA2(13), B(12) => DATA2(12), B(11) => DATA2(11), 
                           B(10) => DATA2(10), B(9) => DATA2(9), B(8) => 
                           DATA2(8), B(7) => DATA2(7), B(6) => DATA2(6), B(5) 
                           => DATA2(5), B(4) => DATA2(4), B(3) => DATA2(3), 
                           B(2) => DATA2(2), B(1) => DATA2(1), B(0) => DATA2(0)
                           , mulin_flag => N3, CLK => CLK, RST => n1, MULready 
                           => RD_sel_flag_port, P(63) => H_MULOUT(31), P(62) =>
                           H_MULOUT(30), P(61) => H_MULOUT(29), P(60) => 
                           H_MULOUT(28), P(59) => H_MULOUT(27), P(58) => 
                           H_MULOUT(26), P(57) => H_MULOUT(25), P(56) => 
                           H_MULOUT(24), P(55) => H_MULOUT(23), P(54) => 
                           H_MULOUT(22), P(53) => H_MULOUT(21), P(52) => 
                           H_MULOUT(20), P(51) => H_MULOUT(19), P(50) => 
                           H_MULOUT(18), P(49) => H_MULOUT(17), P(48) => 
                           H_MULOUT(16), P(47) => H_MULOUT(15), P(46) => 
                           H_MULOUT(14), P(45) => H_MULOUT(13), P(44) => 
                           H_MULOUT(12), P(43) => H_MULOUT(11), P(42) => 
                           H_MULOUT(10), P(41) => H_MULOUT(9), P(40) => 
                           H_MULOUT(8), P(39) => H_MULOUT(7), P(38) => 
                           H_MULOUT(6), P(37) => H_MULOUT(5), P(36) => 
                           H_MULOUT(4), P(35) => H_MULOUT(3), P(34) => 
                           H_MULOUT(2), P(33) => H_MULOUT(1), P(32) => 
                           H_MULOUT(0), P(31) => s_mul_out_31_port, P(30) => 
                           s_mul_out_30_port, P(29) => s_mul_out_29_port, P(28)
                           => s_mul_out_28_port, P(27) => s_mul_out_27_port, 
                           P(26) => s_mul_out_26_port, P(25) => 
                           s_mul_out_25_port, P(24) => s_mul_out_24_port, P(23)
                           => s_mul_out_23_port, P(22) => s_mul_out_22_port, 
                           P(21) => s_mul_out_21_port, P(20) => 
                           s_mul_out_20_port, P(19) => s_mul_out_19_port, P(18)
                           => s_mul_out_18_port, P(17) => s_mul_out_17_port, 
                           P(16) => s_mul_out_16_port, P(15) => 
                           s_mul_out_15_port, P(14) => s_mul_out_14_port, P(13)
                           => s_mul_out_13_port, P(12) => s_mul_out_12_port, 
                           P(11) => s_mul_out_11_port, P(10) => 
                           s_mul_out_10_port, P(9) => s_mul_out_9_port, P(8) =>
                           s_mul_out_8_port, P(7) => s_mul_out_7_port, P(6) => 
                           s_mul_out_6_port, P(5) => s_mul_out_5_port, P(4) => 
                           s_mul_out_4_port, P(3) => s_mul_out_3_port, P(2) => 
                           s_mul_out_2_port, P(1) => s_mul_out_1_port, P(0) => 
                           s_mul_out_0_port);
   OUTPUT_MUX : MUX21_GENERIC_NBIT32_1 port map( A(31) => s_ALUout_31_port, 
                           A(30) => s_ALUout_30_port, A(29) => s_ALUout_29_port
                           , A(28) => s_ALUout_28_port, A(27) => 
                           s_ALUout_27_port, A(26) => s_ALUout_26_port, A(25) 
                           => s_ALUout_25_port, A(24) => s_ALUout_24_port, 
                           A(23) => s_ALUout_23_port, A(22) => s_ALUout_22_port
                           , A(21) => s_ALUout_21_port, A(20) => 
                           s_ALUout_20_port, A(19) => s_ALUout_19_port, A(18) 
                           => s_ALUout_18_port, A(17) => s_ALUout_17_port, 
                           A(16) => s_ALUout_16_port, A(15) => s_ALUout_15_port
                           , A(14) => s_ALUout_14_port, A(13) => 
                           s_ALUout_13_port, A(12) => s_ALUout_12_port, A(11) 
                           => s_ALUout_11_port, A(10) => s_ALUout_10_port, A(9)
                           => s_ALUout_9_port, A(8) => s_ALUout_8_port, A(7) =>
                           s_ALUout_7_port, A(6) => s_ALUout_6_port, A(5) => 
                           s_ALUout_5_port, A(4) => s_ALUout_4_port, A(3) => 
                           s_ALUout_3_port, A(2) => s_ALUout_2_port, A(1) => 
                           s_ALUout_1_port, A(0) => s_ALUout_0_port, B(31) => 
                           s_mul_out_31_port, B(30) => s_mul_out_30_port, B(29)
                           => s_mul_out_29_port, B(28) => s_mul_out_28_port, 
                           B(27) => s_mul_out_27_port, B(26) => 
                           s_mul_out_26_port, B(25) => s_mul_out_25_port, B(24)
                           => s_mul_out_24_port, B(23) => s_mul_out_23_port, 
                           B(22) => s_mul_out_22_port, B(21) => 
                           s_mul_out_21_port, B(20) => s_mul_out_20_port, B(19)
                           => s_mul_out_19_port, B(18) => s_mul_out_18_port, 
                           B(17) => s_mul_out_17_port, B(16) => 
                           s_mul_out_16_port, B(15) => s_mul_out_15_port, B(14)
                           => s_mul_out_14_port, B(13) => s_mul_out_13_port, 
                           B(12) => s_mul_out_12_port, B(11) => 
                           s_mul_out_11_port, B(10) => s_mul_out_10_port, B(9) 
                           => s_mul_out_9_port, B(8) => s_mul_out_8_port, B(7) 
                           => s_mul_out_7_port, B(6) => s_mul_out_6_port, B(5) 
                           => s_mul_out_5_port, B(4) => s_mul_out_4_port, B(3) 
                           => s_mul_out_3_port, B(2) => s_mul_out_2_port, B(1) 
                           => s_mul_out_1_port, B(0) => s_mul_out_0_port, SEL 
                           => RD_sel_flag_port, Y(31) => OUTPUT(31), Y(30) => 
                           OUTPUT(30), Y(29) => OUTPUT(29), Y(28) => OUTPUT(28)
                           , Y(27) => OUTPUT(27), Y(26) => OUTPUT(26), Y(25) =>
                           OUTPUT(25), Y(24) => OUTPUT(24), Y(23) => OUTPUT(23)
                           , Y(22) => OUTPUT(22), Y(21) => OUTPUT(21), Y(20) =>
                           OUTPUT(20), Y(19) => OUTPUT(19), Y(18) => OUTPUT(18)
                           , Y(17) => OUTPUT(17), Y(16) => OUTPUT(16), Y(15) =>
                           OUTPUT(15), Y(14) => OUTPUT(14), Y(13) => OUTPUT(13)
                           , Y(12) => OUTPUT(12), Y(11) => OUTPUT(11), Y(10) =>
                           OUTPUT(10), Y(9) => OUTPUT(9), Y(8) => OUTPUT(8), 
                           Y(7) => OUTPUT(7), Y(6) => OUTPUT(6), Y(5) => 
                           OUTPUT(5), Y(4) => OUTPUT(4), Y(3) => OUTPUT(3), 
                           Y(2) => OUTPUT(2), Y(1) => OUTPUT(1), Y(0) => 
                           OUTPUT(0));
   U3 : BUF_X1 port map( A => RST, Z => n1);
   U4 : AND4_X1 port map( A1 => FUNC(3), A2 => FUNC(2), A3 => FUNC(1), A4 => 
                           FUNC(0), ZN => N3);
   U5 : AND2_X1 port map( A1 => RD_in(4), A2 => N3, ZN => s_RD_in_4_port);
   U6 : AND2_X1 port map( A1 => RD_in(2), A2 => N3, ZN => s_RD_in_2_port);
   U7 : AND2_X1 port map( A1 => RD_in(0), A2 => N3, ZN => s_RD_in_0_port);
   U8 : AND2_X1 port map( A1 => RD_in(1), A2 => N3, ZN => s_RD_in_1_port);
   U9 : AND2_X1 port map( A1 => RD_in(3), A2 => N3, ZN => s_RD_in_3_port);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT5_0 is

   port( A, B : in std_logic_vector (4 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (4 downto 0));

end MUX21_GENERIC_NBIT5_0;

architecture SYN_structural of MUX21_GENERIC_NBIT5_0 is

   component MUX21_462
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_463
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_464
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_465
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_466
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;

begin
   
   MUXES_0 : MUX21_466 port map( A => A(0), B => B(0), S => SEL, Y => Y(0));
   MUXES_1 : MUX21_465 port map( A => A(1), B => B(1), S => SEL, Y => Y(1));
   MUXES_2 : MUX21_464 port map( A => A(2), B => B(2), S => SEL, Y => Y(2));
   MUXES_3 : MUX21_463 port map( A => A(3), B => B(3), S => SEL, Y => Y(3));
   MUXES_4 : MUX21_462 port map( A => A(4), B => B(4), S => SEL, Y => Y(4));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX41_GENERIC_NBIT32_0 is

   port( A, B, C, D : in std_logic_vector (31 downto 0);  SEL : in 
         std_logic_vector (1 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end MUX41_GENERIC_NBIT32_0;

architecture SYN_structural of MUX41_GENERIC_NBIT32_0 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX41_137
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_138
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_139
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_140
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_141
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_142
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_143
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_144
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_145
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_146
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_147
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_148
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_149
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_150
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_151
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_152
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_153
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_154
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_155
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_156
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_157
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_158
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_159
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_160
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_161
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_162
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_163
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_164
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_165
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_166
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_167
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   component MUX41_0
      port( A, B, C, D : in std_logic;  S : in std_logic_vector (1 downto 0);  
            Y : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6 : std_logic;

begin
   
   MUXES_0 : MUX41_0 port map( A => A(0), B => B(0), C => C(0), D => D(0), S(1)
                           => n6, S(0) => n3, Y => Y(0));
   MUXES_1 : MUX41_167 port map( A => A(1), B => B(1), C => C(1), D => D(1), 
                           S(1) => n4, S(0) => n1, Y => Y(1));
   MUXES_2 : MUX41_166 port map( A => A(2), B => B(2), C => C(2), D => D(2), 
                           S(1) => n4, S(0) => n1, Y => Y(2));
   MUXES_3 : MUX41_165 port map( A => A(3), B => B(3), C => C(3), D => D(3), 
                           S(1) => n4, S(0) => n1, Y => Y(3));
   MUXES_4 : MUX41_164 port map( A => A(4), B => B(4), C => C(4), D => D(4), 
                           S(1) => n4, S(0) => n1, Y => Y(4));
   MUXES_5 : MUX41_163 port map( A => A(5), B => B(5), C => C(5), D => D(5), 
                           S(1) => n4, S(0) => n1, Y => Y(5));
   MUXES_6 : MUX41_162 port map( A => A(6), B => B(6), C => C(6), D => D(6), 
                           S(1) => n4, S(0) => n1, Y => Y(6));
   MUXES_7 : MUX41_161 port map( A => A(7), B => B(7), C => C(7), D => D(7), 
                           S(1) => n4, S(0) => n1, Y => Y(7));
   MUXES_8 : MUX41_160 port map( A => A(8), B => B(8), C => C(8), D => D(8), 
                           S(1) => n4, S(0) => n1, Y => Y(8));
   MUXES_9 : MUX41_159 port map( A => A(9), B => B(9), C => C(9), D => D(9), 
                           S(1) => n4, S(0) => n1, Y => Y(9));
   MUXES_10 : MUX41_158 port map( A => A(10), B => B(10), C => C(10), D => 
                           D(10), S(1) => n4, S(0) => n1, Y => Y(10));
   MUXES_11 : MUX41_157 port map( A => A(11), B => B(11), C => C(11), D => 
                           D(11), S(1) => n4, S(0) => n1, Y => Y(11));
   MUXES_12 : MUX41_156 port map( A => A(12), B => B(12), C => C(12), D => 
                           D(12), S(1) => n4, S(0) => n2, Y => Y(12));
   MUXES_13 : MUX41_155 port map( A => A(13), B => B(13), C => C(13), D => 
                           D(13), S(1) => n5, S(0) => n2, Y => Y(13));
   MUXES_14 : MUX41_154 port map( A => A(14), B => B(14), C => C(14), D => 
                           D(14), S(1) => n5, S(0) => n2, Y => Y(14));
   MUXES_15 : MUX41_153 port map( A => A(15), B => B(15), C => C(15), D => 
                           D(15), S(1) => n5, S(0) => n2, Y => Y(15));
   MUXES_16 : MUX41_152 port map( A => A(16), B => B(16), C => C(16), D => 
                           D(16), S(1) => n5, S(0) => n2, Y => Y(16));
   MUXES_17 : MUX41_151 port map( A => A(17), B => B(17), C => C(17), D => 
                           D(17), S(1) => n5, S(0) => n2, Y => Y(17));
   MUXES_18 : MUX41_150 port map( A => A(18), B => B(18), C => C(18), D => 
                           D(18), S(1) => n5, S(0) => n2, Y => Y(18));
   MUXES_19 : MUX41_149 port map( A => A(19), B => B(19), C => C(19), D => 
                           D(19), S(1) => n5, S(0) => n2, Y => Y(19));
   MUXES_20 : MUX41_148 port map( A => A(20), B => B(20), C => C(20), D => 
                           D(20), S(1) => n5, S(0) => n2, Y => Y(20));
   MUXES_21 : MUX41_147 port map( A => A(21), B => B(21), C => C(21), D => 
                           D(21), S(1) => n5, S(0) => n2, Y => Y(21));
   MUXES_22 : MUX41_146 port map( A => A(22), B => B(22), C => C(22), D => 
                           D(22), S(1) => n5, S(0) => n2, Y => Y(22));
   MUXES_23 : MUX41_145 port map( A => A(23), B => B(23), C => C(23), D => 
                           D(23), S(1) => n5, S(0) => n3, Y => Y(23));
   MUXES_24 : MUX41_144 port map( A => A(24), B => B(24), C => C(24), D => 
                           D(24), S(1) => n5, S(0) => n3, Y => Y(24));
   MUXES_25 : MUX41_143 port map( A => A(25), B => B(25), C => C(25), D => 
                           D(25), S(1) => n6, S(0) => n3, Y => Y(25));
   MUXES_26 : MUX41_142 port map( A => A(26), B => B(26), C => C(26), D => 
                           D(26), S(1) => n6, S(0) => n3, Y => Y(26));
   MUXES_27 : MUX41_141 port map( A => A(27), B => B(27), C => C(27), D => 
                           D(27), S(1) => n6, S(0) => n3, Y => Y(27));
   MUXES_28 : MUX41_140 port map( A => A(28), B => B(28), C => C(28), D => 
                           D(28), S(1) => n6, S(0) => n3, Y => Y(28));
   MUXES_29 : MUX41_139 port map( A => A(29), B => B(29), C => C(29), D => 
                           D(29), S(1) => n6, S(0) => n3, Y => Y(29));
   MUXES_30 : MUX41_138 port map( A => A(30), B => B(30), C => C(30), D => 
                           D(30), S(1) => n6, S(0) => n3, Y => Y(30));
   MUXES_31 : MUX41_137 port map( A => A(31), B => B(31), C => C(31), D => 
                           D(31), S(1) => n6, S(0) => n3, Y => Y(31));
   U1 : BUF_X1 port map( A => SEL(1), Z => n4);
   U2 : BUF_X1 port map( A => SEL(1), Z => n5);
   U3 : BUF_X1 port map( A => SEL(1), Z => n6);
   U4 : BUF_X1 port map( A => SEL(0), Z => n1);
   U5 : BUF_X1 port map( A => SEL(0), Z => n2);
   U6 : BUF_X1 port map( A => SEL(0), Z => n3);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity forwarding_unit_WORD_size32_NREG32 is

   port( RSA, RSB : in std_logic_vector (4 downto 0);  ALU_outmem, WB_out : in 
         std_logic_vector (31 downto 0);  MEM_RD, WB_RD : in std_logic_vector 
         (4 downto 0);  LD_EN, WB_EN, S1, S2 : in std_logic;  SEL1, SEL2, SEL3 
         : out std_logic_vector (1 downto 0));

end forwarding_unit_WORD_size32_NREG32;

architecture SYN_Structural of forwarding_unit_WORD_size32_NREG32 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal SEL3_1_port, SEL3_0_port, N30, N31, N32, N49, N50, N51, n1, n2, n3, 
      n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
      n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30_port, n31_port, 
      n32_port, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44 : 
      std_logic;

begin
   SEL3 <= ( SEL3_1_port, SEL3_0_port );
   
   SEL1_reg_1_inst : DLH_X1 port map( G => N30, D => N32, Q => SEL1(1));
   SEL1_reg_0_inst : DLH_X1 port map( G => N30, D => N31, Q => SEL1(0));
   SEL2_reg_1_inst : DLH_X1 port map( G => N49, D => N51, Q => SEL2(1));
   SEL2_reg_0_inst : DLH_X1 port map( G => N49, D => N50, Q => SEL2(0));
   U3 : NAND2_X1 port map( A1 => SEL3_0_port, A2 => n1, ZN => SEL3_1_port);
   U4 : NAND3_X1 port map( A1 => n2, A2 => n3, A3 => WB_EN, ZN => n1);
   U5 : INV_X1 port map( A => n4, ZN => N50);
   U6 : AOI21_X1 port map( B1 => SEL3_0_port, B2 => n5, A => S2, ZN => n4);
   U7 : INV_X1 port map( A => n6, ZN => n5);
   U8 : OAI211_X1 port map( C1 => n7, C2 => n8, A => SEL3_0_port, B => N51, ZN 
                           => N49);
   U9 : NOR2_X1 port map( A1 => n6, A2 => S2, ZN => N51);
   U10 : OAI21_X1 port map( B1 => n9, B2 => n2, A => n3, ZN => n6);
   U11 : INV_X1 port map( A => n7, ZN => n2);
   U12 : NAND3_X1 port map( A1 => n3, A2 => n10, A3 => n9, ZN => SEL3_0_port);
   U13 : AND4_X1 port map( A1 => n11, A2 => n12, A3 => n13, A4 => n14, ZN => n9
                           );
   U14 : NOR2_X1 port map( A1 => n15, A2 => n16, ZN => n14);
   U15 : XOR2_X1 port map( A => RSB(4), B => MEM_RD(4), Z => n16);
   U16 : XOR2_X1 port map( A => RSB(3), B => MEM_RD(3), Z => n15);
   U17 : XNOR2_X1 port map( A => MEM_RD(1), B => RSB(1), ZN => n13);
   U18 : XNOR2_X1 port map( A => MEM_RD(2), B => RSB(2), ZN => n12);
   U19 : XNOR2_X1 port map( A => MEM_RD(0), B => RSB(0), ZN => n11);
   U20 : INV_X1 port map( A => LD_EN, ZN => n10);
   U21 : OR4_X1 port map( A1 => RSB(3), A2 => RSB(4), A3 => RSB(2), A4 => n17, 
                           ZN => n3);
   U22 : OR2_X1 port map( A1 => RSB(1), A2 => RSB(0), ZN => n17);
   U23 : NAND4_X1 port map( A1 => n18, A2 => n19, A3 => n20, A4 => n21, ZN => 
                           n7);
   U24 : NOR2_X1 port map( A1 => n22, A2 => n23, ZN => n21);
   U25 : XOR2_X1 port map( A => WB_RD(4), B => RSB(4), Z => n23);
   U26 : XOR2_X1 port map( A => WB_RD(3), B => RSB(3), Z => n22);
   U27 : XNOR2_X1 port map( A => RSB(1), B => WB_RD(1), ZN => n20);
   U28 : XNOR2_X1 port map( A => RSB(2), B => WB_RD(2), ZN => n19);
   U29 : XNOR2_X1 port map( A => RSB(0), B => WB_RD(0), ZN => n18);
   U30 : AOI21_X1 port map( B1 => n24, B2 => n25, A => n26, ZN => N31);
   U31 : INV_X1 port map( A => n27, ZN => n25);
   U32 : NOR2_X1 port map( A1 => LD_EN, A2 => n28, ZN => n24);
   U33 : OAI221_X1 port map( B1 => LD_EN, B2 => n27, C1 => n8, C2 => n29, A => 
                           N32, ZN => N30);
   U34 : NOR2_X1 port map( A1 => n26, A2 => n28, ZN => N32);
   U35 : INV_X1 port map( A => n30_port, ZN => n28);
   U36 : AOI21_X1 port map( B1 => n27, B2 => n29, A => n31_port, ZN => n30_port
                           );
   U37 : NOR4_X1 port map( A1 => RSA(3), A2 => RSA(4), A3 => RSA(2), A4 => 
                           n32_port, ZN => n31_port);
   U38 : OR2_X1 port map( A1 => RSA(1), A2 => RSA(0), ZN => n32_port);
   U39 : INV_X1 port map( A => S1, ZN => n26);
   U40 : NAND4_X1 port map( A1 => n33, A2 => n34, A3 => n35, A4 => n36, ZN => 
                           n29);
   U41 : NOR2_X1 port map( A1 => n37, A2 => n38, ZN => n36);
   U42 : XOR2_X1 port map( A => WB_RD(4), B => RSA(4), Z => n38);
   U43 : XOR2_X1 port map( A => WB_RD(3), B => RSA(3), Z => n37);
   U44 : XNOR2_X1 port map( A => RSA(1), B => WB_RD(1), ZN => n35);
   U45 : XNOR2_X1 port map( A => RSA(2), B => WB_RD(2), ZN => n34);
   U46 : XNOR2_X1 port map( A => RSA(0), B => WB_RD(0), ZN => n33);
   U47 : INV_X1 port map( A => WB_EN, ZN => n8);
   U48 : NAND4_X1 port map( A1 => n39, A2 => n40, A3 => n41, A4 => n42, ZN => 
                           n27);
   U49 : NOR2_X1 port map( A1 => n43, A2 => n44, ZN => n42);
   U50 : XOR2_X1 port map( A => RSA(4), B => MEM_RD(4), Z => n44);
   U51 : XOR2_X1 port map( A => RSA(3), B => MEM_RD(3), Z => n43);
   U52 : XNOR2_X1 port map( A => MEM_RD(1), B => RSA(1), ZN => n41);
   U53 : XNOR2_X1 port map( A => MEM_RD(2), B => RSA(2), ZN => n40);
   U54 : XNOR2_X1 port map( A => MEM_RD(0), B => RSA(0), ZN => n39);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity register_file_NBIT32_NREG32 is

   port( RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, ADD_RD2 
         : in std_logic_vector (4 downto 0);  DATAIN : in std_logic_vector (31 
         downto 0);  OUT1, OUT2 : out std_logic_vector (31 downto 0));

end register_file_NBIT32_NREG32;

architecture SYN_Behavioral of register_file_NBIT32_NREG32 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal REGISTERS_0_31_port, REGISTERS_0_30_port, REGISTERS_0_29_port, 
      REGISTERS_0_28_port, REGISTERS_0_27_port, REGISTERS_0_26_port, 
      REGISTERS_0_25_port, REGISTERS_0_24_port, REGISTERS_0_23_port, 
      REGISTERS_0_22_port, REGISTERS_0_21_port, REGISTERS_0_20_port, 
      REGISTERS_0_19_port, REGISTERS_0_18_port, REGISTERS_0_17_port, 
      REGISTERS_0_16_port, REGISTERS_0_15_port, REGISTERS_0_14_port, 
      REGISTERS_0_13_port, REGISTERS_0_12_port, REGISTERS_0_11_port, 
      REGISTERS_0_10_port, REGISTERS_0_9_port, REGISTERS_0_8_port, 
      REGISTERS_0_7_port, REGISTERS_0_6_port, REGISTERS_0_5_port, 
      REGISTERS_0_4_port, REGISTERS_0_3_port, REGISTERS_0_2_port, 
      REGISTERS_0_1_port, REGISTERS_0_0_port, REGISTERS_1_31_port, 
      REGISTERS_1_30_port, REGISTERS_1_29_port, REGISTERS_1_28_port, 
      REGISTERS_1_27_port, REGISTERS_1_26_port, REGISTERS_1_25_port, 
      REGISTERS_1_24_port, REGISTERS_1_23_port, REGISTERS_1_22_port, 
      REGISTERS_1_21_port, REGISTERS_1_20_port, REGISTERS_1_19_port, 
      REGISTERS_1_18_port, REGISTERS_1_17_port, REGISTERS_1_16_port, 
      REGISTERS_1_15_port, REGISTERS_1_14_port, REGISTERS_1_13_port, 
      REGISTERS_1_12_port, REGISTERS_1_11_port, REGISTERS_1_10_port, 
      REGISTERS_1_9_port, REGISTERS_1_8_port, REGISTERS_1_7_port, 
      REGISTERS_1_6_port, REGISTERS_1_5_port, REGISTERS_1_4_port, 
      REGISTERS_1_3_port, REGISTERS_1_2_port, REGISTERS_1_1_port, 
      REGISTERS_1_0_port, REGISTERS_2_31_port, REGISTERS_2_30_port, 
      REGISTERS_2_29_port, REGISTERS_2_28_port, REGISTERS_2_27_port, 
      REGISTERS_2_26_port, REGISTERS_2_25_port, REGISTERS_2_24_port, 
      REGISTERS_2_23_port, REGISTERS_2_22_port, REGISTERS_2_21_port, 
      REGISTERS_2_20_port, REGISTERS_2_19_port, REGISTERS_2_18_port, 
      REGISTERS_2_17_port, REGISTERS_2_16_port, REGISTERS_2_15_port, 
      REGISTERS_2_14_port, REGISTERS_2_13_port, REGISTERS_2_12_port, 
      REGISTERS_2_11_port, REGISTERS_2_10_port, REGISTERS_2_9_port, 
      REGISTERS_2_8_port, REGISTERS_2_7_port, REGISTERS_2_6_port, 
      REGISTERS_2_5_port, REGISTERS_2_4_port, REGISTERS_2_3_port, 
      REGISTERS_2_2_port, REGISTERS_2_1_port, REGISTERS_2_0_port, 
      REGISTERS_3_31_port, REGISTERS_3_30_port, REGISTERS_3_29_port, 
      REGISTERS_3_28_port, REGISTERS_3_27_port, REGISTERS_3_26_port, 
      REGISTERS_3_25_port, REGISTERS_3_24_port, REGISTERS_3_23_port, 
      REGISTERS_3_22_port, REGISTERS_3_21_port, REGISTERS_3_20_port, 
      REGISTERS_3_19_port, REGISTERS_3_18_port, REGISTERS_3_17_port, 
      REGISTERS_3_16_port, REGISTERS_3_15_port, REGISTERS_3_14_port, 
      REGISTERS_3_13_port, REGISTERS_3_12_port, REGISTERS_3_11_port, 
      REGISTERS_3_10_port, REGISTERS_3_9_port, REGISTERS_3_8_port, 
      REGISTERS_3_7_port, REGISTERS_3_6_port, REGISTERS_3_5_port, 
      REGISTERS_3_4_port, REGISTERS_3_3_port, REGISTERS_3_2_port, 
      REGISTERS_3_1_port, REGISTERS_3_0_port, REGISTERS_4_31_port, 
      REGISTERS_4_30_port, REGISTERS_4_29_port, REGISTERS_4_28_port, 
      REGISTERS_4_27_port, REGISTERS_4_26_port, REGISTERS_4_25_port, 
      REGISTERS_4_24_port, REGISTERS_4_23_port, REGISTERS_4_22_port, 
      REGISTERS_4_21_port, REGISTERS_4_20_port, REGISTERS_4_19_port, 
      REGISTERS_4_18_port, REGISTERS_4_17_port, REGISTERS_4_16_port, 
      REGISTERS_4_15_port, REGISTERS_4_14_port, REGISTERS_4_13_port, 
      REGISTERS_4_12_port, REGISTERS_4_11_port, REGISTERS_4_10_port, 
      REGISTERS_4_9_port, REGISTERS_4_8_port, REGISTERS_4_7_port, 
      REGISTERS_4_6_port, REGISTERS_4_5_port, REGISTERS_4_4_port, 
      REGISTERS_4_3_port, REGISTERS_4_2_port, REGISTERS_4_1_port, 
      REGISTERS_4_0_port, REGISTERS_5_31_port, REGISTERS_5_30_port, 
      REGISTERS_5_29_port, REGISTERS_5_28_port, REGISTERS_5_27_port, 
      REGISTERS_5_26_port, REGISTERS_5_25_port, REGISTERS_5_24_port, 
      REGISTERS_5_23_port, REGISTERS_5_22_port, REGISTERS_5_21_port, 
      REGISTERS_5_20_port, REGISTERS_5_19_port, REGISTERS_5_18_port, 
      REGISTERS_5_17_port, REGISTERS_5_16_port, REGISTERS_5_15_port, 
      REGISTERS_5_14_port, REGISTERS_5_13_port, REGISTERS_5_12_port, 
      REGISTERS_5_11_port, REGISTERS_5_10_port, REGISTERS_5_9_port, 
      REGISTERS_5_8_port, REGISTERS_5_7_port, REGISTERS_5_6_port, 
      REGISTERS_5_5_port, REGISTERS_5_4_port, REGISTERS_5_3_port, 
      REGISTERS_5_2_port, REGISTERS_5_1_port, REGISTERS_5_0_port, 
      REGISTERS_6_31_port, REGISTERS_6_30_port, REGISTERS_6_29_port, 
      REGISTERS_6_28_port, REGISTERS_6_27_port, REGISTERS_6_26_port, 
      REGISTERS_6_25_port, REGISTERS_6_24_port, REGISTERS_6_23_port, 
      REGISTERS_6_22_port, REGISTERS_6_21_port, REGISTERS_6_20_port, 
      REGISTERS_6_19_port, REGISTERS_6_18_port, REGISTERS_6_17_port, 
      REGISTERS_6_16_port, REGISTERS_6_15_port, REGISTERS_6_14_port, 
      REGISTERS_6_13_port, REGISTERS_6_12_port, REGISTERS_6_11_port, 
      REGISTERS_6_10_port, REGISTERS_6_9_port, REGISTERS_6_8_port, 
      REGISTERS_6_7_port, REGISTERS_6_6_port, REGISTERS_6_5_port, 
      REGISTERS_6_4_port, REGISTERS_6_3_port, REGISTERS_6_2_port, 
      REGISTERS_6_1_port, REGISTERS_6_0_port, REGISTERS_7_31_port, 
      REGISTERS_7_30_port, REGISTERS_7_29_port, REGISTERS_7_28_port, 
      REGISTERS_7_27_port, REGISTERS_7_26_port, REGISTERS_7_25_port, 
      REGISTERS_7_24_port, REGISTERS_7_23_port, REGISTERS_7_22_port, 
      REGISTERS_7_21_port, REGISTERS_7_20_port, REGISTERS_7_19_port, 
      REGISTERS_7_18_port, REGISTERS_7_17_port, REGISTERS_7_16_port, 
      REGISTERS_7_15_port, REGISTERS_7_14_port, REGISTERS_7_13_port, 
      REGISTERS_7_12_port, REGISTERS_7_11_port, REGISTERS_7_10_port, 
      REGISTERS_7_9_port, REGISTERS_7_8_port, REGISTERS_7_7_port, 
      REGISTERS_7_6_port, REGISTERS_7_5_port, REGISTERS_7_4_port, 
      REGISTERS_7_3_port, REGISTERS_7_2_port, REGISTERS_7_1_port, 
      REGISTERS_7_0_port, REGISTERS_8_31_port, REGISTERS_8_30_port, 
      REGISTERS_8_29_port, REGISTERS_8_28_port, REGISTERS_8_27_port, 
      REGISTERS_8_26_port, REGISTERS_8_25_port, REGISTERS_8_24_port, 
      REGISTERS_8_23_port, REGISTERS_8_22_port, REGISTERS_8_21_port, 
      REGISTERS_8_20_port, REGISTERS_8_19_port, REGISTERS_8_18_port, 
      REGISTERS_8_17_port, REGISTERS_8_16_port, REGISTERS_8_15_port, 
      REGISTERS_8_14_port, REGISTERS_8_13_port, REGISTERS_8_12_port, 
      REGISTERS_8_11_port, REGISTERS_8_10_port, REGISTERS_8_9_port, 
      REGISTERS_8_8_port, REGISTERS_8_7_port, REGISTERS_8_6_port, 
      REGISTERS_8_5_port, REGISTERS_8_4_port, REGISTERS_8_3_port, 
      REGISTERS_8_2_port, REGISTERS_8_1_port, REGISTERS_8_0_port, 
      REGISTERS_9_31_port, REGISTERS_9_30_port, REGISTERS_9_29_port, 
      REGISTERS_9_28_port, REGISTERS_9_27_port, REGISTERS_9_26_port, 
      REGISTERS_9_25_port, REGISTERS_9_24_port, REGISTERS_9_23_port, 
      REGISTERS_9_22_port, REGISTERS_9_21_port, REGISTERS_9_20_port, 
      REGISTERS_9_19_port, REGISTERS_9_18_port, REGISTERS_9_17_port, 
      REGISTERS_9_16_port, REGISTERS_9_15_port, REGISTERS_9_14_port, 
      REGISTERS_9_13_port, REGISTERS_9_12_port, REGISTERS_9_11_port, 
      REGISTERS_9_10_port, REGISTERS_9_9_port, REGISTERS_9_8_port, 
      REGISTERS_9_7_port, REGISTERS_9_6_port, REGISTERS_9_5_port, 
      REGISTERS_9_4_port, REGISTERS_9_3_port, REGISTERS_9_2_port, 
      REGISTERS_9_1_port, REGISTERS_9_0_port, REGISTERS_10_31_port, 
      REGISTERS_10_30_port, REGISTERS_10_29_port, REGISTERS_10_28_port, 
      REGISTERS_10_27_port, REGISTERS_10_26_port, REGISTERS_10_25_port, 
      REGISTERS_10_24_port, REGISTERS_10_23_port, REGISTERS_10_22_port, 
      REGISTERS_10_21_port, REGISTERS_10_20_port, REGISTERS_10_19_port, 
      REGISTERS_10_18_port, REGISTERS_10_17_port, REGISTERS_10_16_port, 
      REGISTERS_10_15_port, REGISTERS_10_14_port, REGISTERS_10_13_port, 
      REGISTERS_10_12_port, REGISTERS_10_11_port, REGISTERS_10_10_port, 
      REGISTERS_10_9_port, REGISTERS_10_8_port, REGISTERS_10_7_port, 
      REGISTERS_10_6_port, REGISTERS_10_5_port, REGISTERS_10_4_port, 
      REGISTERS_10_3_port, REGISTERS_10_2_port, REGISTERS_10_1_port, 
      REGISTERS_10_0_port, REGISTERS_11_31_port, REGISTERS_11_30_port, 
      REGISTERS_11_29_port, REGISTERS_11_28_port, REGISTERS_11_27_port, 
      REGISTERS_11_26_port, REGISTERS_11_25_port, REGISTERS_11_24_port, 
      REGISTERS_11_23_port, REGISTERS_11_22_port, REGISTERS_11_21_port, 
      REGISTERS_11_20_port, REGISTERS_11_19_port, REGISTERS_11_18_port, 
      REGISTERS_11_17_port, REGISTERS_11_16_port, REGISTERS_11_15_port, 
      REGISTERS_11_14_port, REGISTERS_11_13_port, REGISTERS_11_12_port, 
      REGISTERS_11_11_port, REGISTERS_11_10_port, REGISTERS_11_9_port, 
      REGISTERS_11_8_port, REGISTERS_11_7_port, REGISTERS_11_6_port, 
      REGISTERS_11_5_port, REGISTERS_11_4_port, REGISTERS_11_3_port, 
      REGISTERS_11_2_port, REGISTERS_11_1_port, REGISTERS_11_0_port, 
      REGISTERS_12_31_port, REGISTERS_12_30_port, REGISTERS_12_29_port, 
      REGISTERS_12_28_port, REGISTERS_12_27_port, REGISTERS_12_26_port, 
      REGISTERS_12_25_port, REGISTERS_12_24_port, REGISTERS_12_23_port, 
      REGISTERS_12_22_port, REGISTERS_12_21_port, REGISTERS_12_20_port, 
      REGISTERS_12_19_port, REGISTERS_12_18_port, REGISTERS_12_17_port, 
      REGISTERS_12_16_port, REGISTERS_12_15_port, REGISTERS_12_14_port, 
      REGISTERS_12_13_port, REGISTERS_12_12_port, REGISTERS_12_11_port, 
      REGISTERS_12_10_port, REGISTERS_12_9_port, REGISTERS_12_8_port, 
      REGISTERS_12_7_port, REGISTERS_12_6_port, REGISTERS_12_5_port, 
      REGISTERS_12_4_port, REGISTERS_12_3_port, REGISTERS_12_2_port, 
      REGISTERS_12_1_port, REGISTERS_12_0_port, REGISTERS_13_31_port, 
      REGISTERS_13_30_port, REGISTERS_13_29_port, REGISTERS_13_28_port, 
      REGISTERS_13_27_port, REGISTERS_13_26_port, REGISTERS_13_25_port, 
      REGISTERS_13_24_port, REGISTERS_13_23_port, REGISTERS_13_22_port, 
      REGISTERS_13_21_port, REGISTERS_13_20_port, REGISTERS_13_19_port, 
      REGISTERS_13_18_port, REGISTERS_13_17_port, REGISTERS_13_16_port, 
      REGISTERS_13_15_port, REGISTERS_13_14_port, REGISTERS_13_13_port, 
      REGISTERS_13_12_port, REGISTERS_13_11_port, REGISTERS_13_10_port, 
      REGISTERS_13_9_port, REGISTERS_13_8_port, REGISTERS_13_7_port, 
      REGISTERS_13_6_port, REGISTERS_13_5_port, REGISTERS_13_4_port, 
      REGISTERS_13_3_port, REGISTERS_13_2_port, REGISTERS_13_1_port, 
      REGISTERS_13_0_port, REGISTERS_14_31_port, REGISTERS_14_30_port, 
      REGISTERS_14_29_port, REGISTERS_14_28_port, REGISTERS_14_27_port, 
      REGISTERS_14_26_port, REGISTERS_14_25_port, REGISTERS_14_24_port, 
      REGISTERS_14_23_port, REGISTERS_14_22_port, REGISTERS_14_21_port, 
      REGISTERS_14_20_port, REGISTERS_14_19_port, REGISTERS_14_18_port, 
      REGISTERS_14_17_port, REGISTERS_14_16_port, REGISTERS_14_15_port, 
      REGISTERS_14_14_port, REGISTERS_14_13_port, REGISTERS_14_12_port, 
      REGISTERS_14_11_port, REGISTERS_14_10_port, REGISTERS_14_9_port, 
      REGISTERS_14_8_port, REGISTERS_14_7_port, REGISTERS_14_6_port, 
      REGISTERS_14_5_port, REGISTERS_14_4_port, REGISTERS_14_3_port, 
      REGISTERS_14_2_port, REGISTERS_14_1_port, REGISTERS_14_0_port, 
      REGISTERS_15_31_port, REGISTERS_15_30_port, REGISTERS_15_29_port, 
      REGISTERS_15_28_port, REGISTERS_15_27_port, REGISTERS_15_26_port, 
      REGISTERS_15_25_port, REGISTERS_15_24_port, REGISTERS_15_23_port, 
      REGISTERS_15_22_port, REGISTERS_15_21_port, REGISTERS_15_20_port, 
      REGISTERS_15_19_port, REGISTERS_15_18_port, REGISTERS_15_17_port, 
      REGISTERS_15_16_port, REGISTERS_15_15_port, REGISTERS_15_14_port, 
      REGISTERS_15_13_port, REGISTERS_15_12_port, REGISTERS_15_11_port, 
      REGISTERS_15_10_port, REGISTERS_15_9_port, REGISTERS_15_8_port, 
      REGISTERS_15_7_port, REGISTERS_15_6_port, REGISTERS_15_5_port, 
      REGISTERS_15_4_port, REGISTERS_15_3_port, REGISTERS_15_2_port, 
      REGISTERS_15_1_port, REGISTERS_15_0_port, REGISTERS_16_31_port, 
      REGISTERS_16_30_port, REGISTERS_16_29_port, REGISTERS_16_28_port, 
      REGISTERS_16_27_port, REGISTERS_16_26_port, REGISTERS_16_25_port, 
      REGISTERS_16_24_port, REGISTERS_16_23_port, REGISTERS_16_22_port, 
      REGISTERS_16_21_port, REGISTERS_16_20_port, REGISTERS_16_19_port, 
      REGISTERS_16_18_port, REGISTERS_16_17_port, REGISTERS_16_16_port, 
      REGISTERS_16_15_port, REGISTERS_16_14_port, REGISTERS_16_13_port, 
      REGISTERS_16_12_port, REGISTERS_16_11_port, REGISTERS_16_10_port, 
      REGISTERS_16_9_port, REGISTERS_16_8_port, REGISTERS_16_7_port, 
      REGISTERS_16_6_port, REGISTERS_16_5_port, REGISTERS_16_4_port, 
      REGISTERS_16_3_port, REGISTERS_16_2_port, REGISTERS_16_1_port, 
      REGISTERS_16_0_port, REGISTERS_17_31_port, REGISTERS_17_30_port, 
      REGISTERS_17_29_port, REGISTERS_17_28_port, REGISTERS_17_27_port, 
      REGISTERS_17_26_port, REGISTERS_17_25_port, REGISTERS_17_24_port, 
      REGISTERS_17_23_port, REGISTERS_17_22_port, REGISTERS_17_21_port, 
      REGISTERS_17_20_port, REGISTERS_17_19_port, REGISTERS_17_18_port, 
      REGISTERS_17_17_port, REGISTERS_17_16_port, REGISTERS_17_15_port, 
      REGISTERS_17_14_port, REGISTERS_17_13_port, REGISTERS_17_12_port, 
      REGISTERS_17_11_port, REGISTERS_17_10_port, REGISTERS_17_9_port, 
      REGISTERS_17_8_port, REGISTERS_17_7_port, REGISTERS_17_6_port, 
      REGISTERS_17_5_port, REGISTERS_17_4_port, REGISTERS_17_3_port, 
      REGISTERS_17_2_port, REGISTERS_17_1_port, REGISTERS_17_0_port, 
      REGISTERS_18_31_port, REGISTERS_18_30_port, REGISTERS_18_29_port, 
      REGISTERS_18_28_port, REGISTERS_18_27_port, REGISTERS_18_26_port, 
      REGISTERS_18_25_port, REGISTERS_18_24_port, REGISTERS_18_23_port, 
      REGISTERS_18_22_port, REGISTERS_18_21_port, REGISTERS_18_20_port, 
      REGISTERS_18_19_port, REGISTERS_18_18_port, REGISTERS_18_17_port, 
      REGISTERS_18_16_port, REGISTERS_18_15_port, REGISTERS_18_14_port, 
      REGISTERS_18_13_port, REGISTERS_18_12_port, REGISTERS_18_11_port, 
      REGISTERS_18_10_port, REGISTERS_18_9_port, REGISTERS_18_8_port, 
      REGISTERS_18_7_port, REGISTERS_18_6_port, REGISTERS_18_5_port, 
      REGISTERS_18_4_port, REGISTERS_18_3_port, REGISTERS_18_2_port, 
      REGISTERS_18_1_port, REGISTERS_18_0_port, REGISTERS_19_31_port, 
      REGISTERS_19_30_port, REGISTERS_19_29_port, REGISTERS_19_28_port, 
      REGISTERS_19_27_port, REGISTERS_19_26_port, REGISTERS_19_25_port, 
      REGISTERS_19_24_port, REGISTERS_19_23_port, REGISTERS_19_22_port, 
      REGISTERS_19_21_port, REGISTERS_19_20_port, REGISTERS_19_19_port, 
      REGISTERS_19_18_port, REGISTERS_19_17_port, REGISTERS_19_16_port, 
      REGISTERS_19_15_port, REGISTERS_19_14_port, REGISTERS_19_13_port, 
      REGISTERS_19_12_port, REGISTERS_19_11_port, REGISTERS_19_10_port, 
      REGISTERS_19_9_port, REGISTERS_19_8_port, REGISTERS_19_7_port, 
      REGISTERS_19_6_port, REGISTERS_19_5_port, REGISTERS_19_4_port, 
      REGISTERS_19_3_port, REGISTERS_19_2_port, REGISTERS_19_1_port, 
      REGISTERS_19_0_port, REGISTERS_20_31_port, REGISTERS_20_30_port, 
      REGISTERS_20_29_port, REGISTERS_20_28_port, REGISTERS_20_27_port, 
      REGISTERS_20_26_port, REGISTERS_20_25_port, REGISTERS_20_24_port, 
      REGISTERS_20_23_port, REGISTERS_20_22_port, REGISTERS_20_21_port, 
      REGISTERS_20_20_port, REGISTERS_20_19_port, REGISTERS_20_18_port, 
      REGISTERS_20_17_port, REGISTERS_20_16_port, REGISTERS_20_15_port, 
      REGISTERS_20_14_port, REGISTERS_20_13_port, REGISTERS_20_12_port, 
      REGISTERS_20_11_port, REGISTERS_20_10_port, REGISTERS_20_9_port, 
      REGISTERS_20_8_port, REGISTERS_20_7_port, REGISTERS_20_6_port, 
      REGISTERS_20_5_port, REGISTERS_20_4_port, REGISTERS_20_3_port, 
      REGISTERS_20_2_port, REGISTERS_20_1_port, REGISTERS_20_0_port, 
      REGISTERS_21_31_port, REGISTERS_21_30_port, REGISTERS_21_29_port, 
      REGISTERS_21_28_port, REGISTERS_21_27_port, REGISTERS_21_26_port, 
      REGISTERS_21_25_port, REGISTERS_21_24_port, REGISTERS_21_23_port, 
      REGISTERS_21_22_port, REGISTERS_21_21_port, REGISTERS_21_20_port, 
      REGISTERS_21_19_port, REGISTERS_21_18_port, REGISTERS_21_17_port, 
      REGISTERS_21_16_port, REGISTERS_21_15_port, REGISTERS_21_14_port, 
      REGISTERS_21_13_port, REGISTERS_21_12_port, REGISTERS_21_11_port, 
      REGISTERS_21_10_port, REGISTERS_21_9_port, REGISTERS_21_8_port, 
      REGISTERS_21_7_port, REGISTERS_21_6_port, REGISTERS_21_5_port, 
      REGISTERS_21_4_port, REGISTERS_21_3_port, REGISTERS_21_2_port, 
      REGISTERS_21_1_port, REGISTERS_21_0_port, REGISTERS_22_31_port, 
      REGISTERS_22_30_port, REGISTERS_22_29_port, REGISTERS_22_28_port, 
      REGISTERS_22_27_port, REGISTERS_22_26_port, REGISTERS_22_25_port, 
      REGISTERS_22_24_port, REGISTERS_22_23_port, REGISTERS_22_22_port, 
      REGISTERS_22_21_port, REGISTERS_22_20_port, REGISTERS_22_19_port, 
      REGISTERS_22_18_port, REGISTERS_22_17_port, REGISTERS_22_16_port, 
      REGISTERS_22_15_port, REGISTERS_22_14_port, REGISTERS_22_13_port, 
      REGISTERS_22_12_port, REGISTERS_22_11_port, REGISTERS_22_10_port, 
      REGISTERS_22_9_port, REGISTERS_22_8_port, REGISTERS_22_7_port, 
      REGISTERS_22_6_port, REGISTERS_22_5_port, REGISTERS_22_4_port, 
      REGISTERS_22_3_port, REGISTERS_22_2_port, REGISTERS_22_1_port, 
      REGISTERS_22_0_port, REGISTERS_23_31_port, REGISTERS_23_30_port, 
      REGISTERS_23_29_port, REGISTERS_23_28_port, REGISTERS_23_27_port, 
      REGISTERS_23_26_port, REGISTERS_23_25_port, REGISTERS_23_24_port, 
      REGISTERS_23_23_port, REGISTERS_23_22_port, REGISTERS_23_21_port, 
      REGISTERS_23_20_port, REGISTERS_23_19_port, REGISTERS_23_18_port, 
      REGISTERS_23_17_port, REGISTERS_23_16_port, REGISTERS_23_15_port, 
      REGISTERS_23_14_port, REGISTERS_23_13_port, REGISTERS_23_12_port, 
      REGISTERS_23_11_port, REGISTERS_23_10_port, REGISTERS_23_9_port, 
      REGISTERS_23_8_port, REGISTERS_23_7_port, REGISTERS_23_6_port, 
      REGISTERS_23_5_port, REGISTERS_23_4_port, REGISTERS_23_3_port, 
      REGISTERS_23_2_port, REGISTERS_23_1_port, REGISTERS_23_0_port, 
      REGISTERS_24_31_port, REGISTERS_24_30_port, REGISTERS_24_29_port, 
      REGISTERS_24_28_port, REGISTERS_24_27_port, REGISTERS_24_26_port, 
      REGISTERS_24_25_port, REGISTERS_24_24_port, REGISTERS_24_23_port, 
      REGISTERS_24_22_port, REGISTERS_24_21_port, REGISTERS_24_20_port, 
      REGISTERS_24_19_port, REGISTERS_24_18_port, REGISTERS_24_17_port, 
      REGISTERS_24_16_port, REGISTERS_24_15_port, REGISTERS_24_14_port, 
      REGISTERS_24_13_port, REGISTERS_24_12_port, REGISTERS_24_11_port, 
      REGISTERS_24_10_port, REGISTERS_24_9_port, REGISTERS_24_8_port, 
      REGISTERS_24_7_port, REGISTERS_24_6_port, REGISTERS_24_5_port, 
      REGISTERS_24_4_port, REGISTERS_24_3_port, REGISTERS_24_2_port, 
      REGISTERS_24_1_port, REGISTERS_24_0_port, REGISTERS_25_31_port, 
      REGISTERS_25_30_port, REGISTERS_25_29_port, REGISTERS_25_28_port, 
      REGISTERS_25_27_port, REGISTERS_25_26_port, REGISTERS_25_25_port, 
      REGISTERS_25_24_port, REGISTERS_25_23_port, REGISTERS_25_22_port, 
      REGISTERS_25_21_port, REGISTERS_25_20_port, REGISTERS_25_19_port, 
      REGISTERS_25_18_port, REGISTERS_25_17_port, REGISTERS_25_16_port, 
      REGISTERS_25_15_port, REGISTERS_25_14_port, REGISTERS_25_13_port, 
      REGISTERS_25_12_port, REGISTERS_25_11_port, REGISTERS_25_10_port, 
      REGISTERS_25_9_port, REGISTERS_25_8_port, REGISTERS_25_7_port, 
      REGISTERS_25_6_port, REGISTERS_25_5_port, REGISTERS_25_4_port, 
      REGISTERS_25_3_port, REGISTERS_25_2_port, REGISTERS_25_1_port, 
      REGISTERS_25_0_port, REGISTERS_26_31_port, REGISTERS_26_30_port, 
      REGISTERS_26_29_port, REGISTERS_26_28_port, REGISTERS_26_27_port, 
      REGISTERS_26_26_port, REGISTERS_26_25_port, REGISTERS_26_24_port, 
      REGISTERS_26_23_port, REGISTERS_26_22_port, REGISTERS_26_21_port, 
      REGISTERS_26_20_port, REGISTERS_26_19_port, REGISTERS_26_18_port, 
      REGISTERS_26_17_port, REGISTERS_26_16_port, REGISTERS_26_15_port, 
      REGISTERS_26_14_port, REGISTERS_26_13_port, REGISTERS_26_12_port, 
      REGISTERS_26_11_port, REGISTERS_26_10_port, REGISTERS_26_9_port, 
      REGISTERS_26_8_port, REGISTERS_26_7_port, REGISTERS_26_6_port, 
      REGISTERS_26_5_port, REGISTERS_26_4_port, REGISTERS_26_3_port, 
      REGISTERS_26_2_port, REGISTERS_26_1_port, REGISTERS_26_0_port, 
      REGISTERS_27_31_port, REGISTERS_27_30_port, REGISTERS_27_29_port, 
      REGISTERS_27_28_port, REGISTERS_27_27_port, REGISTERS_27_26_port, 
      REGISTERS_27_25_port, REGISTERS_27_24_port, REGISTERS_27_23_port, 
      REGISTERS_27_22_port, REGISTERS_27_21_port, REGISTERS_27_20_port, 
      REGISTERS_27_19_port, REGISTERS_27_18_port, REGISTERS_27_17_port, 
      REGISTERS_27_16_port, REGISTERS_27_15_port, REGISTERS_27_14_port, 
      REGISTERS_27_13_port, REGISTERS_27_12_port, REGISTERS_27_11_port, 
      REGISTERS_27_10_port, REGISTERS_27_9_port, REGISTERS_27_8_port, 
      REGISTERS_27_7_port, REGISTERS_27_6_port, REGISTERS_27_5_port, 
      REGISTERS_27_4_port, REGISTERS_27_3_port, REGISTERS_27_2_port, 
      REGISTERS_27_1_port, REGISTERS_27_0_port, REGISTERS_28_31_port, 
      REGISTERS_28_30_port, REGISTERS_28_29_port, REGISTERS_28_28_port, 
      REGISTERS_28_27_port, REGISTERS_28_26_port, REGISTERS_28_25_port, 
      REGISTERS_28_24_port, REGISTERS_28_23_port, REGISTERS_28_22_port, 
      REGISTERS_28_21_port, REGISTERS_28_20_port, REGISTERS_28_19_port, 
      REGISTERS_28_18_port, REGISTERS_28_17_port, REGISTERS_28_16_port, 
      REGISTERS_28_15_port, REGISTERS_28_14_port, REGISTERS_28_13_port, 
      REGISTERS_28_12_port, REGISTERS_28_11_port, REGISTERS_28_10_port, 
      REGISTERS_28_9_port, REGISTERS_28_8_port, REGISTERS_28_7_port, 
      REGISTERS_28_6_port, REGISTERS_28_5_port, REGISTERS_28_4_port, 
      REGISTERS_28_3_port, REGISTERS_28_2_port, REGISTERS_28_1_port, 
      REGISTERS_28_0_port, REGISTERS_29_31_port, REGISTERS_29_30_port, 
      REGISTERS_29_29_port, REGISTERS_29_28_port, REGISTERS_29_27_port, 
      REGISTERS_29_26_port, REGISTERS_29_25_port, REGISTERS_29_24_port, 
      REGISTERS_29_23_port, REGISTERS_29_22_port, REGISTERS_29_21_port, 
      REGISTERS_29_20_port, REGISTERS_29_19_port, REGISTERS_29_18_port, 
      REGISTERS_29_17_port, REGISTERS_29_16_port, REGISTERS_29_15_port, 
      REGISTERS_29_14_port, REGISTERS_29_13_port, REGISTERS_29_12_port, 
      REGISTERS_29_11_port, REGISTERS_29_10_port, REGISTERS_29_9_port, 
      REGISTERS_29_8_port, REGISTERS_29_7_port, REGISTERS_29_6_port, 
      REGISTERS_29_5_port, REGISTERS_29_4_port, REGISTERS_29_3_port, 
      REGISTERS_29_2_port, REGISTERS_29_1_port, REGISTERS_29_0_port, 
      REGISTERS_30_31_port, REGISTERS_30_30_port, REGISTERS_30_29_port, 
      REGISTERS_30_28_port, REGISTERS_30_27_port, REGISTERS_30_26_port, 
      REGISTERS_30_25_port, REGISTERS_30_24_port, REGISTERS_30_23_port, 
      REGISTERS_30_22_port, REGISTERS_30_21_port, REGISTERS_30_20_port, 
      REGISTERS_30_19_port, REGISTERS_30_18_port, REGISTERS_30_17_port, 
      REGISTERS_30_16_port, REGISTERS_30_15_port, REGISTERS_30_14_port, 
      REGISTERS_30_13_port, REGISTERS_30_12_port, REGISTERS_30_11_port, 
      REGISTERS_30_10_port, REGISTERS_30_9_port, REGISTERS_30_8_port, 
      REGISTERS_30_7_port, REGISTERS_30_6_port, REGISTERS_30_5_port, 
      REGISTERS_30_4_port, REGISTERS_30_3_port, REGISTERS_30_2_port, 
      REGISTERS_30_1_port, REGISTERS_30_0_port, REGISTERS_31_31_port, 
      REGISTERS_31_30_port, REGISTERS_31_29_port, REGISTERS_31_28_port, 
      REGISTERS_31_27_port, REGISTERS_31_26_port, REGISTERS_31_25_port, 
      REGISTERS_31_24_port, REGISTERS_31_23_port, REGISTERS_31_22_port, 
      REGISTERS_31_21_port, REGISTERS_31_20_port, REGISTERS_31_19_port, 
      REGISTERS_31_18_port, REGISTERS_31_17_port, REGISTERS_31_16_port, 
      REGISTERS_31_15_port, REGISTERS_31_14_port, REGISTERS_31_13_port, 
      REGISTERS_31_12_port, REGISTERS_31_11_port, REGISTERS_31_10_port, 
      REGISTERS_31_9_port, REGISTERS_31_8_port, REGISTERS_31_7_port, 
      REGISTERS_31_6_port, REGISTERS_31_5_port, REGISTERS_31_4_port, 
      REGISTERS_31_3_port, REGISTERS_31_2_port, REGISTERS_31_1_port, 
      REGISTERS_31_0_port, N312, N313, N314, N315, N316, N317, N318, N319, N320
      , N321, N322, N323, N324, N325, N326, N327, N328, N329, N330, N331, N332,
      N333, N334, N335, N336, N337, N338, N339, N340, N341, N342, N343, N344, 
      N345, N346, N347, N348, N349, N350, N351, N352, N353, N354, N355, N356, 
      N357, N358, N359, N360, N361, N362, N363, N364, N365, N366, N367, N368, 
      N369, N370, N371, N372, N373, N374, N375, N376, N377, N378, N379, N380, 
      N381, N382, N383, N384, N385, N386, N387, N388, N389, N390, N391, N392, 
      N393, N394, N395, N396, N397, N398, N399, N400, N401, N402, N403, N404, 
      N405, N406, N407, N408, N409, N410, N411, N412, N413, N414, N415, N416, 
      N417, N418, N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, 
      N429, N430, N431, N432, N433, N434, N435, N436, N437, N438, N439, N440, 
      N441, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, 
      n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, 
      n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, 
      n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, 
      n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, 
      n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, 
      n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, 
      n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, 
      n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, 
      n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, 
      n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, 
      n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, 
      n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, 
      n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, 
      n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, 
      n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, 
      n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, 
      n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, 
      n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, 
      n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, 
      n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, 
      n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, 
      n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, 
      n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, 
      n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, 
      n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, 
      n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, 
      n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, 
      n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, 
      n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, 
      n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, 
      n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, 
      n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, 
      n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, 
      n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, 
      n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, 
      n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, 
      n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, 
      n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, 
      n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, 
      n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, 
      n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, 
      n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, 
      n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, 
      n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, 
      n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, 
      n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, 
      n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, 
      n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, 
      n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, 
      n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, 
      n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, 
      n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, 
      n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, 
      n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, 
      n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, 
      n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, 
      n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, 
      n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, 
      n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, 
      n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, 
      n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, 
      n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, 
      n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, 
      n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, 
      n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, 
      n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, 
      n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, 
      n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, 
      n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, 
      n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, 
      n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, 
      n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, 
      n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, 
      n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, 
      n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, 
      n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, 
      n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, 
      n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, 
      n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, 
      n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, 
      n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, 
      n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, 
      n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, 
      n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, 
      n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, 
      n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, 
      n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, 
      n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, 
      n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, 
      n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, 
      n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, 
      n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, 
      n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, 
      n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, 
      n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, 
      n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, 
      n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, 
      n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, 
      n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, 
      n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, 
      n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, 
      n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, 
      n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, 
      n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, 
      n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, 
      n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, 
      n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, 
      n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, 
      n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, 
      n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, 
      n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, 
      n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, 
      n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, 
      n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, 
      n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, 
      n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, 
      n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, 
      n1785, n1786, n1787, n1788, n1789, n1790, n1, n2, n3, n4, n5, n6, n7, n8,
      n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
      n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38
      , n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, 
      n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67
      , n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, 
      n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96
      , n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, 
      n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, 
      n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, 
      n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, 
      n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, 
      n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, 
      n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, 
      n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, 
      n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, 
      n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, 
      n312_port, n313_port, n314_port, n315_port, n316_port, n317_port, 
      n318_port, n319_port, n320_port, n321_port, n322_port, n323_port, 
      n324_port, n325_port, n326_port, n327_port, n328_port, n329_port, 
      n330_port, n331_port, n332_port, n333_port, n334_port, n335_port, 
      n336_port, n337_port, n338_port, n339_port, n340_port, n341_port, 
      n342_port, n343_port, n344_port, n345_port, n346_port, n347_port, 
      n348_port, n349_port, n350_port, n351_port, n352_port, n353_port, 
      n354_port, n355_port, n356_port, n357_port, n358_port, n359_port, 
      n360_port, n361_port, n362_port, n363_port, n364_port, n365_port, 
      n366_port, n367_port, n368_port, n369_port, n370_port, n371_port, 
      n372_port, n373_port, n374_port, n375_port, n376_port, n377_port, 
      n378_port, n379_port, n380_port, n381_port, n382_port, n383_port, 
      n384_port, n385_port, n386_port, n387_port, n388_port, n389_port, 
      n390_port, n391_port, n392_port, n393_port, n394_port, n395_port, 
      n396_port, n397_port, n398_port, n399_port, n400_port, n401_port, 
      n402_port, n403_port, n404_port, n405_port, n406_port, n407_port, 
      n408_port, n409_port, n410_port, n411_port, n412_port, n413_port, 
      n414_port, n415_port, n416_port, n417_port, n418_port, n419_port, 
      n420_port, n421_port, n422_port, n423_port, n424_port, n425_port, 
      n426_port, n427_port, n428_port, n429_port, n430_port, n431_port, 
      n432_port, n433_port, n434_port, n435_port, n436_port, n437_port, 
      n438_port, n439_port, n440_port, n441_port, n442, n443, n444, n445, n446,
      n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, 
      n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, 
      n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, 
      n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, 
      n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, 
      n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, 
      n519, n520, n521, n522, n523, n524, n525, n526, n1791, n1792, n1793, 
      n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, 
      n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, 
      n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, 
      n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, 
      n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, 
      n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, 
      n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, 
      n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, 
      n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, 
      n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, 
      n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, 
      n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, 
      n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, 
      n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, 
      n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, 
      n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, 
      n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, 
      n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, 
      n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, 
      n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, 
      n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, 
      n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, 
      n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, 
      n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, 
      n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, 
      n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, 
      n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, 
      n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, 
      n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, 
      n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, 
      n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, 
      n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, 
      n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, 
      n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, 
      n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, 
      n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, 
      n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, 
      n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, 
      n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, 
      n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, 
      n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, 
      n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, 
      n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, 
      n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, 
      n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, 
      n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, 
      n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263 : 
      std_logic;

begin
   
   REGISTERS_reg_0_31_inst : DLH_X1 port map( G => n204, D => n328_port, Q => 
                           REGISTERS_0_31_port);
   REGISTERS_reg_0_30_inst : DLH_X1 port map( G => n204, D => n332_port, Q => 
                           REGISTERS_0_30_port);
   REGISTERS_reg_0_29_inst : DLH_X1 port map( G => n204, D => n336_port, Q => 
                           REGISTERS_0_29_port);
   REGISTERS_reg_0_28_inst : DLH_X1 port map( G => n204, D => n340_port, Q => 
                           REGISTERS_0_28_port);
   REGISTERS_reg_0_27_inst : DLH_X1 port map( G => n204, D => n344_port, Q => 
                           REGISTERS_0_27_port);
   REGISTERS_reg_0_26_inst : DLH_X1 port map( G => n204, D => n348_port, Q => 
                           REGISTERS_0_26_port);
   REGISTERS_reg_0_25_inst : DLH_X1 port map( G => n204, D => n352_port, Q => 
                           REGISTERS_0_25_port);
   REGISTERS_reg_0_24_inst : DLH_X1 port map( G => n204, D => n356_port, Q => 
                           REGISTERS_0_24_port);
   REGISTERS_reg_0_23_inst : DLH_X1 port map( G => n204, D => n360_port, Q => 
                           REGISTERS_0_23_port);
   REGISTERS_reg_0_22_inst : DLH_X1 port map( G => n204, D => n364_port, Q => 
                           REGISTERS_0_22_port);
   REGISTERS_reg_0_21_inst : DLH_X1 port map( G => n205, D => n368_port, Q => 
                           REGISTERS_0_21_port);
   REGISTERS_reg_0_20_inst : DLH_X1 port map( G => n205, D => n372_port, Q => 
                           REGISTERS_0_20_port);
   REGISTERS_reg_0_19_inst : DLH_X1 port map( G => n205, D => n376_port, Q => 
                           REGISTERS_0_19_port);
   REGISTERS_reg_0_18_inst : DLH_X1 port map( G => n205, D => n380_port, Q => 
                           REGISTERS_0_18_port);
   REGISTERS_reg_0_17_inst : DLH_X1 port map( G => n205, D => n384_port, Q => 
                           REGISTERS_0_17_port);
   REGISTERS_reg_0_16_inst : DLH_X1 port map( G => n205, D => n388_port, Q => 
                           REGISTERS_0_16_port);
   REGISTERS_reg_0_15_inst : DLH_X1 port map( G => n205, D => n392_port, Q => 
                           REGISTERS_0_15_port);
   REGISTERS_reg_0_14_inst : DLH_X1 port map( G => n205, D => n396_port, Q => 
                           REGISTERS_0_14_port);
   REGISTERS_reg_0_13_inst : DLH_X1 port map( G => n205, D => n400_port, Q => 
                           REGISTERS_0_13_port);
   REGISTERS_reg_0_12_inst : DLH_X1 port map( G => n205, D => n404_port, Q => 
                           REGISTERS_0_12_port);
   REGISTERS_reg_0_11_inst : DLH_X1 port map( G => n206, D => n408_port, Q => 
                           REGISTERS_0_11_port);
   REGISTERS_reg_0_10_inst : DLH_X1 port map( G => n206, D => n412_port, Q => 
                           REGISTERS_0_10_port);
   REGISTERS_reg_0_9_inst : DLH_X1 port map( G => n206, D => n416_port, Q => 
                           REGISTERS_0_9_port);
   REGISTERS_reg_0_8_inst : DLH_X1 port map( G => n206, D => n420_port, Q => 
                           REGISTERS_0_8_port);
   REGISTERS_reg_0_7_inst : DLH_X1 port map( G => n206, D => n424_port, Q => 
                           REGISTERS_0_7_port);
   REGISTERS_reg_0_6_inst : DLH_X1 port map( G => n206, D => n428_port, Q => 
                           REGISTERS_0_6_port);
   REGISTERS_reg_0_5_inst : DLH_X1 port map( G => n206, D => n432_port, Q => 
                           REGISTERS_0_5_port);
   REGISTERS_reg_0_4_inst : DLH_X1 port map( G => n206, D => n436_port, Q => 
                           REGISTERS_0_4_port);
   REGISTERS_reg_0_3_inst : DLH_X1 port map( G => n206, D => n440_port, Q => 
                           REGISTERS_0_3_port);
   REGISTERS_reg_0_2_inst : DLH_X1 port map( G => n206, D => n444, Q => 
                           REGISTERS_0_2_port);
   REGISTERS_reg_0_1_inst : DLH_X1 port map( G => n207, D => n448, Q => 
                           REGISTERS_0_1_port);
   REGISTERS_reg_0_0_inst : DLH_X1 port map( G => n207, D => n452, Q => 
                           REGISTERS_0_0_port);
   REGISTERS_reg_1_31_inst : DLH_X1 port map( G => n211, D => n328_port, Q => 
                           REGISTERS_1_31_port);
   REGISTERS_reg_1_30_inst : DLH_X1 port map( G => n211, D => n332_port, Q => 
                           REGISTERS_1_30_port);
   REGISTERS_reg_1_29_inst : DLH_X1 port map( G => n210, D => n336_port, Q => 
                           REGISTERS_1_29_port);
   REGISTERS_reg_1_28_inst : DLH_X1 port map( G => n210, D => n340_port, Q => 
                           REGISTERS_1_28_port);
   REGISTERS_reg_1_27_inst : DLH_X1 port map( G => n210, D => n344_port, Q => 
                           REGISTERS_1_27_port);
   REGISTERS_reg_1_26_inst : DLH_X1 port map( G => n210, D => n348_port, Q => 
                           REGISTERS_1_26_port);
   REGISTERS_reg_1_25_inst : DLH_X1 port map( G => n210, D => n352_port, Q => 
                           REGISTERS_1_25_port);
   REGISTERS_reg_1_24_inst : DLH_X1 port map( G => n210, D => n356_port, Q => 
                           REGISTERS_1_24_port);
   REGISTERS_reg_1_23_inst : DLH_X1 port map( G => n210, D => n360_port, Q => 
                           REGISTERS_1_23_port);
   REGISTERS_reg_1_22_inst : DLH_X1 port map( G => n210, D => n364_port, Q => 
                           REGISTERS_1_22_port);
   REGISTERS_reg_1_21_inst : DLH_X1 port map( G => n210, D => n368_port, Q => 
                           REGISTERS_1_21_port);
   REGISTERS_reg_1_20_inst : DLH_X1 port map( G => n210, D => n372_port, Q => 
                           REGISTERS_1_20_port);
   REGISTERS_reg_1_19_inst : DLH_X1 port map( G => n209, D => n376_port, Q => 
                           REGISTERS_1_19_port);
   REGISTERS_reg_1_18_inst : DLH_X1 port map( G => n209, D => n380_port, Q => 
                           REGISTERS_1_18_port);
   REGISTERS_reg_1_17_inst : DLH_X1 port map( G => n209, D => n384_port, Q => 
                           REGISTERS_1_17_port);
   REGISTERS_reg_1_16_inst : DLH_X1 port map( G => n209, D => n388_port, Q => 
                           REGISTERS_1_16_port);
   REGISTERS_reg_1_15_inst : DLH_X1 port map( G => n209, D => n392_port, Q => 
                           REGISTERS_1_15_port);
   REGISTERS_reg_1_14_inst : DLH_X1 port map( G => n209, D => n396_port, Q => 
                           REGISTERS_1_14_port);
   REGISTERS_reg_1_13_inst : DLH_X1 port map( G => n209, D => n400_port, Q => 
                           REGISTERS_1_13_port);
   REGISTERS_reg_1_12_inst : DLH_X1 port map( G => n209, D => n404_port, Q => 
                           REGISTERS_1_12_port);
   REGISTERS_reg_1_11_inst : DLH_X1 port map( G => n209, D => n408_port, Q => 
                           REGISTERS_1_11_port);
   REGISTERS_reg_1_10_inst : DLH_X1 port map( G => n209, D => n412_port, Q => 
                           REGISTERS_1_10_port);
   REGISTERS_reg_1_9_inst : DLH_X1 port map( G => n208, D => n416_port, Q => 
                           REGISTERS_1_9_port);
   REGISTERS_reg_1_8_inst : DLH_X1 port map( G => n208, D => n420_port, Q => 
                           REGISTERS_1_8_port);
   REGISTERS_reg_1_7_inst : DLH_X1 port map( G => n208, D => n424_port, Q => 
                           REGISTERS_1_7_port);
   REGISTERS_reg_1_6_inst : DLH_X1 port map( G => n208, D => n428_port, Q => 
                           REGISTERS_1_6_port);
   REGISTERS_reg_1_5_inst : DLH_X1 port map( G => n208, D => n432_port, Q => 
                           REGISTERS_1_5_port);
   REGISTERS_reg_1_4_inst : DLH_X1 port map( G => n208, D => n436_port, Q => 
                           REGISTERS_1_4_port);
   REGISTERS_reg_1_3_inst : DLH_X1 port map( G => n208, D => n440_port, Q => 
                           REGISTERS_1_3_port);
   REGISTERS_reg_1_2_inst : DLH_X1 port map( G => n208, D => n444, Q => 
                           REGISTERS_1_2_port);
   REGISTERS_reg_1_1_inst : DLH_X1 port map( G => n208, D => n448, Q => 
                           REGISTERS_1_1_port);
   REGISTERS_reg_1_0_inst : DLH_X1 port map( G => n208, D => n452, Q => 
                           REGISTERS_1_0_port);
   REGISTERS_reg_2_31_inst : DLH_X1 port map( G => n215, D => n328_port, Q => 
                           REGISTERS_2_31_port);
   REGISTERS_reg_2_30_inst : DLH_X1 port map( G => n215, D => n332_port, Q => 
                           REGISTERS_2_30_port);
   REGISTERS_reg_2_29_inst : DLH_X1 port map( G => n214, D => n336_port, Q => 
                           REGISTERS_2_29_port);
   REGISTERS_reg_2_28_inst : DLH_X1 port map( G => n214, D => n340_port, Q => 
                           REGISTERS_2_28_port);
   REGISTERS_reg_2_27_inst : DLH_X1 port map( G => n214, D => n344_port, Q => 
                           REGISTERS_2_27_port);
   REGISTERS_reg_2_26_inst : DLH_X1 port map( G => n214, D => n348_port, Q => 
                           REGISTERS_2_26_port);
   REGISTERS_reg_2_25_inst : DLH_X1 port map( G => n214, D => n352_port, Q => 
                           REGISTERS_2_25_port);
   REGISTERS_reg_2_24_inst : DLH_X1 port map( G => n214, D => n356_port, Q => 
                           REGISTERS_2_24_port);
   REGISTERS_reg_2_23_inst : DLH_X1 port map( G => n214, D => n360_port, Q => 
                           REGISTERS_2_23_port);
   REGISTERS_reg_2_22_inst : DLH_X1 port map( G => n214, D => n364_port, Q => 
                           REGISTERS_2_22_port);
   REGISTERS_reg_2_21_inst : DLH_X1 port map( G => n214, D => n368_port, Q => 
                           REGISTERS_2_21_port);
   REGISTERS_reg_2_20_inst : DLH_X1 port map( G => n214, D => n372_port, Q => 
                           REGISTERS_2_20_port);
   REGISTERS_reg_2_19_inst : DLH_X1 port map( G => n213, D => n376_port, Q => 
                           REGISTERS_2_19_port);
   REGISTERS_reg_2_18_inst : DLH_X1 port map( G => n213, D => n380_port, Q => 
                           REGISTERS_2_18_port);
   REGISTERS_reg_2_17_inst : DLH_X1 port map( G => n213, D => n384_port, Q => 
                           REGISTERS_2_17_port);
   REGISTERS_reg_2_16_inst : DLH_X1 port map( G => n213, D => n388_port, Q => 
                           REGISTERS_2_16_port);
   REGISTERS_reg_2_15_inst : DLH_X1 port map( G => n213, D => n392_port, Q => 
                           REGISTERS_2_15_port);
   REGISTERS_reg_2_14_inst : DLH_X1 port map( G => n213, D => n396_port, Q => 
                           REGISTERS_2_14_port);
   REGISTERS_reg_2_13_inst : DLH_X1 port map( G => n213, D => n400_port, Q => 
                           REGISTERS_2_13_port);
   REGISTERS_reg_2_12_inst : DLH_X1 port map( G => n213, D => n404_port, Q => 
                           REGISTERS_2_12_port);
   REGISTERS_reg_2_11_inst : DLH_X1 port map( G => n213, D => n408_port, Q => 
                           REGISTERS_2_11_port);
   REGISTERS_reg_2_10_inst : DLH_X1 port map( G => n213, D => n412_port, Q => 
                           REGISTERS_2_10_port);
   REGISTERS_reg_2_9_inst : DLH_X1 port map( G => n212, D => n416_port, Q => 
                           REGISTERS_2_9_port);
   REGISTERS_reg_2_8_inst : DLH_X1 port map( G => n212, D => n420_port, Q => 
                           REGISTERS_2_8_port);
   REGISTERS_reg_2_7_inst : DLH_X1 port map( G => n212, D => n424_port, Q => 
                           REGISTERS_2_7_port);
   REGISTERS_reg_2_6_inst : DLH_X1 port map( G => n212, D => n428_port, Q => 
                           REGISTERS_2_6_port);
   REGISTERS_reg_2_5_inst : DLH_X1 port map( G => n212, D => n432_port, Q => 
                           REGISTERS_2_5_port);
   REGISTERS_reg_2_4_inst : DLH_X1 port map( G => n212, D => n436_port, Q => 
                           REGISTERS_2_4_port);
   REGISTERS_reg_2_3_inst : DLH_X1 port map( G => n212, D => n440_port, Q => 
                           REGISTERS_2_3_port);
   REGISTERS_reg_2_2_inst : DLH_X1 port map( G => n212, D => n444, Q => 
                           REGISTERS_2_2_port);
   REGISTERS_reg_2_1_inst : DLH_X1 port map( G => n212, D => n448, Q => 
                           REGISTERS_2_1_port);
   REGISTERS_reg_2_0_inst : DLH_X1 port map( G => n212, D => n452, Q => 
                           REGISTERS_2_0_port);
   REGISTERS_reg_3_31_inst : DLH_X1 port map( G => n219, D => n328_port, Q => 
                           REGISTERS_3_31_port);
   REGISTERS_reg_3_30_inst : DLH_X1 port map( G => n219, D => n332_port, Q => 
                           REGISTERS_3_30_port);
   REGISTERS_reg_3_29_inst : DLH_X1 port map( G => n218, D => n336_port, Q => 
                           REGISTERS_3_29_port);
   REGISTERS_reg_3_28_inst : DLH_X1 port map( G => n218, D => n340_port, Q => 
                           REGISTERS_3_28_port);
   REGISTERS_reg_3_27_inst : DLH_X1 port map( G => n218, D => n344_port, Q => 
                           REGISTERS_3_27_port);
   REGISTERS_reg_3_26_inst : DLH_X1 port map( G => n218, D => n348_port, Q => 
                           REGISTERS_3_26_port);
   REGISTERS_reg_3_25_inst : DLH_X1 port map( G => n218, D => n352_port, Q => 
                           REGISTERS_3_25_port);
   REGISTERS_reg_3_24_inst : DLH_X1 port map( G => n218, D => n356_port, Q => 
                           REGISTERS_3_24_port);
   REGISTERS_reg_3_23_inst : DLH_X1 port map( G => n218, D => n360_port, Q => 
                           REGISTERS_3_23_port);
   REGISTERS_reg_3_22_inst : DLH_X1 port map( G => n218, D => n364_port, Q => 
                           REGISTERS_3_22_port);
   REGISTERS_reg_3_21_inst : DLH_X1 port map( G => n218, D => n368_port, Q => 
                           REGISTERS_3_21_port);
   REGISTERS_reg_3_20_inst : DLH_X1 port map( G => n218, D => n372_port, Q => 
                           REGISTERS_3_20_port);
   REGISTERS_reg_3_19_inst : DLH_X1 port map( G => n217, D => n376_port, Q => 
                           REGISTERS_3_19_port);
   REGISTERS_reg_3_18_inst : DLH_X1 port map( G => n217, D => n380_port, Q => 
                           REGISTERS_3_18_port);
   REGISTERS_reg_3_17_inst : DLH_X1 port map( G => n217, D => n384_port, Q => 
                           REGISTERS_3_17_port);
   REGISTERS_reg_3_16_inst : DLH_X1 port map( G => n217, D => n388_port, Q => 
                           REGISTERS_3_16_port);
   REGISTERS_reg_3_15_inst : DLH_X1 port map( G => n217, D => n392_port, Q => 
                           REGISTERS_3_15_port);
   REGISTERS_reg_3_14_inst : DLH_X1 port map( G => n217, D => n396_port, Q => 
                           REGISTERS_3_14_port);
   REGISTERS_reg_3_13_inst : DLH_X1 port map( G => n217, D => n400_port, Q => 
                           REGISTERS_3_13_port);
   REGISTERS_reg_3_12_inst : DLH_X1 port map( G => n217, D => n404_port, Q => 
                           REGISTERS_3_12_port);
   REGISTERS_reg_3_11_inst : DLH_X1 port map( G => n217, D => n408_port, Q => 
                           REGISTERS_3_11_port);
   REGISTERS_reg_3_10_inst : DLH_X1 port map( G => n217, D => n412_port, Q => 
                           REGISTERS_3_10_port);
   REGISTERS_reg_3_9_inst : DLH_X1 port map( G => n216, D => n416_port, Q => 
                           REGISTERS_3_9_port);
   REGISTERS_reg_3_8_inst : DLH_X1 port map( G => n216, D => n420_port, Q => 
                           REGISTERS_3_8_port);
   REGISTERS_reg_3_7_inst : DLH_X1 port map( G => n216, D => n424_port, Q => 
                           REGISTERS_3_7_port);
   REGISTERS_reg_3_6_inst : DLH_X1 port map( G => n216, D => n428_port, Q => 
                           REGISTERS_3_6_port);
   REGISTERS_reg_3_5_inst : DLH_X1 port map( G => n216, D => n432_port, Q => 
                           REGISTERS_3_5_port);
   REGISTERS_reg_3_4_inst : DLH_X1 port map( G => n216, D => n436_port, Q => 
                           REGISTERS_3_4_port);
   REGISTERS_reg_3_3_inst : DLH_X1 port map( G => n216, D => n440_port, Q => 
                           REGISTERS_3_3_port);
   REGISTERS_reg_3_2_inst : DLH_X1 port map( G => n216, D => n444, Q => 
                           REGISTERS_3_2_port);
   REGISTERS_reg_3_1_inst : DLH_X1 port map( G => n216, D => n448, Q => 
                           REGISTERS_3_1_port);
   REGISTERS_reg_3_0_inst : DLH_X1 port map( G => n216, D => n452, Q => 
                           REGISTERS_3_0_port);
   REGISTERS_reg_4_31_inst : DLH_X1 port map( G => n223, D => n328_port, Q => 
                           REGISTERS_4_31_port);
   REGISTERS_reg_4_30_inst : DLH_X1 port map( G => n223, D => n332_port, Q => 
                           REGISTERS_4_30_port);
   REGISTERS_reg_4_29_inst : DLH_X1 port map( G => n222, D => n336_port, Q => 
                           REGISTERS_4_29_port);
   REGISTERS_reg_4_28_inst : DLH_X1 port map( G => n222, D => n340_port, Q => 
                           REGISTERS_4_28_port);
   REGISTERS_reg_4_27_inst : DLH_X1 port map( G => n222, D => n344_port, Q => 
                           REGISTERS_4_27_port);
   REGISTERS_reg_4_26_inst : DLH_X1 port map( G => n222, D => n348_port, Q => 
                           REGISTERS_4_26_port);
   REGISTERS_reg_4_25_inst : DLH_X1 port map( G => n222, D => n352_port, Q => 
                           REGISTERS_4_25_port);
   REGISTERS_reg_4_24_inst : DLH_X1 port map( G => n222, D => n356_port, Q => 
                           REGISTERS_4_24_port);
   REGISTERS_reg_4_23_inst : DLH_X1 port map( G => n222, D => n360_port, Q => 
                           REGISTERS_4_23_port);
   REGISTERS_reg_4_22_inst : DLH_X1 port map( G => n222, D => n364_port, Q => 
                           REGISTERS_4_22_port);
   REGISTERS_reg_4_21_inst : DLH_X1 port map( G => n222, D => n368_port, Q => 
                           REGISTERS_4_21_port);
   REGISTERS_reg_4_20_inst : DLH_X1 port map( G => n222, D => n372_port, Q => 
                           REGISTERS_4_20_port);
   REGISTERS_reg_4_19_inst : DLH_X1 port map( G => n221, D => n376_port, Q => 
                           REGISTERS_4_19_port);
   REGISTERS_reg_4_18_inst : DLH_X1 port map( G => n221, D => n380_port, Q => 
                           REGISTERS_4_18_port);
   REGISTERS_reg_4_17_inst : DLH_X1 port map( G => n221, D => n384_port, Q => 
                           REGISTERS_4_17_port);
   REGISTERS_reg_4_16_inst : DLH_X1 port map( G => n221, D => n388_port, Q => 
                           REGISTERS_4_16_port);
   REGISTERS_reg_4_15_inst : DLH_X1 port map( G => n221, D => n392_port, Q => 
                           REGISTERS_4_15_port);
   REGISTERS_reg_4_14_inst : DLH_X1 port map( G => n221, D => n396_port, Q => 
                           REGISTERS_4_14_port);
   REGISTERS_reg_4_13_inst : DLH_X1 port map( G => n221, D => n400_port, Q => 
                           REGISTERS_4_13_port);
   REGISTERS_reg_4_12_inst : DLH_X1 port map( G => n221, D => n404_port, Q => 
                           REGISTERS_4_12_port);
   REGISTERS_reg_4_11_inst : DLH_X1 port map( G => n221, D => n408_port, Q => 
                           REGISTERS_4_11_port);
   REGISTERS_reg_4_10_inst : DLH_X1 port map( G => n221, D => n412_port, Q => 
                           REGISTERS_4_10_port);
   REGISTERS_reg_4_9_inst : DLH_X1 port map( G => n220, D => n416_port, Q => 
                           REGISTERS_4_9_port);
   REGISTERS_reg_4_8_inst : DLH_X1 port map( G => n220, D => n420_port, Q => 
                           REGISTERS_4_8_port);
   REGISTERS_reg_4_7_inst : DLH_X1 port map( G => n220, D => n424_port, Q => 
                           REGISTERS_4_7_port);
   REGISTERS_reg_4_6_inst : DLH_X1 port map( G => n220, D => n428_port, Q => 
                           REGISTERS_4_6_port);
   REGISTERS_reg_4_5_inst : DLH_X1 port map( G => n220, D => n432_port, Q => 
                           REGISTERS_4_5_port);
   REGISTERS_reg_4_4_inst : DLH_X1 port map( G => n220, D => n436_port, Q => 
                           REGISTERS_4_4_port);
   REGISTERS_reg_4_3_inst : DLH_X1 port map( G => n220, D => n440_port, Q => 
                           REGISTERS_4_3_port);
   REGISTERS_reg_4_2_inst : DLH_X1 port map( G => n220, D => n444, Q => 
                           REGISTERS_4_2_port);
   REGISTERS_reg_4_1_inst : DLH_X1 port map( G => n220, D => n448, Q => 
                           REGISTERS_4_1_port);
   REGISTERS_reg_4_0_inst : DLH_X1 port map( G => n220, D => n452, Q => 
                           REGISTERS_4_0_port);
   REGISTERS_reg_5_31_inst : DLH_X1 port map( G => n227, D => n328_port, Q => 
                           REGISTERS_5_31_port);
   REGISTERS_reg_5_30_inst : DLH_X1 port map( G => n227, D => n332_port, Q => 
                           REGISTERS_5_30_port);
   REGISTERS_reg_5_29_inst : DLH_X1 port map( G => n226, D => n336_port, Q => 
                           REGISTERS_5_29_port);
   REGISTERS_reg_5_28_inst : DLH_X1 port map( G => n226, D => n340_port, Q => 
                           REGISTERS_5_28_port);
   REGISTERS_reg_5_27_inst : DLH_X1 port map( G => n226, D => n344_port, Q => 
                           REGISTERS_5_27_port);
   REGISTERS_reg_5_26_inst : DLH_X1 port map( G => n226, D => n348_port, Q => 
                           REGISTERS_5_26_port);
   REGISTERS_reg_5_25_inst : DLH_X1 port map( G => n226, D => n352_port, Q => 
                           REGISTERS_5_25_port);
   REGISTERS_reg_5_24_inst : DLH_X1 port map( G => n226, D => n356_port, Q => 
                           REGISTERS_5_24_port);
   REGISTERS_reg_5_23_inst : DLH_X1 port map( G => n226, D => n360_port, Q => 
                           REGISTERS_5_23_port);
   REGISTERS_reg_5_22_inst : DLH_X1 port map( G => n226, D => n364_port, Q => 
                           REGISTERS_5_22_port);
   REGISTERS_reg_5_21_inst : DLH_X1 port map( G => n226, D => n368_port, Q => 
                           REGISTERS_5_21_port);
   REGISTERS_reg_5_20_inst : DLH_X1 port map( G => n226, D => n372_port, Q => 
                           REGISTERS_5_20_port);
   REGISTERS_reg_5_19_inst : DLH_X1 port map( G => n225, D => n376_port, Q => 
                           REGISTERS_5_19_port);
   REGISTERS_reg_5_18_inst : DLH_X1 port map( G => n225, D => n380_port, Q => 
                           REGISTERS_5_18_port);
   REGISTERS_reg_5_17_inst : DLH_X1 port map( G => n225, D => n384_port, Q => 
                           REGISTERS_5_17_port);
   REGISTERS_reg_5_16_inst : DLH_X1 port map( G => n225, D => n388_port, Q => 
                           REGISTERS_5_16_port);
   REGISTERS_reg_5_15_inst : DLH_X1 port map( G => n225, D => n392_port, Q => 
                           REGISTERS_5_15_port);
   REGISTERS_reg_5_14_inst : DLH_X1 port map( G => n225, D => n396_port, Q => 
                           REGISTERS_5_14_port);
   REGISTERS_reg_5_13_inst : DLH_X1 port map( G => n225, D => n400_port, Q => 
                           REGISTERS_5_13_port);
   REGISTERS_reg_5_12_inst : DLH_X1 port map( G => n225, D => n404_port, Q => 
                           REGISTERS_5_12_port);
   REGISTERS_reg_5_11_inst : DLH_X1 port map( G => n225, D => n408_port, Q => 
                           REGISTERS_5_11_port);
   REGISTERS_reg_5_10_inst : DLH_X1 port map( G => n225, D => n412_port, Q => 
                           REGISTERS_5_10_port);
   REGISTERS_reg_5_9_inst : DLH_X1 port map( G => n224, D => n416_port, Q => 
                           REGISTERS_5_9_port);
   REGISTERS_reg_5_8_inst : DLH_X1 port map( G => n224, D => n420_port, Q => 
                           REGISTERS_5_8_port);
   REGISTERS_reg_5_7_inst : DLH_X1 port map( G => n224, D => n424_port, Q => 
                           REGISTERS_5_7_port);
   REGISTERS_reg_5_6_inst : DLH_X1 port map( G => n224, D => n428_port, Q => 
                           REGISTERS_5_6_port);
   REGISTERS_reg_5_5_inst : DLH_X1 port map( G => n224, D => n432_port, Q => 
                           REGISTERS_5_5_port);
   REGISTERS_reg_5_4_inst : DLH_X1 port map( G => n224, D => n436_port, Q => 
                           REGISTERS_5_4_port);
   REGISTERS_reg_5_3_inst : DLH_X1 port map( G => n224, D => n440_port, Q => 
                           REGISTERS_5_3_port);
   REGISTERS_reg_5_2_inst : DLH_X1 port map( G => n224, D => n444, Q => 
                           REGISTERS_5_2_port);
   REGISTERS_reg_5_1_inst : DLH_X1 port map( G => n224, D => n448, Q => 
                           REGISTERS_5_1_port);
   REGISTERS_reg_5_0_inst : DLH_X1 port map( G => n224, D => n452, Q => 
                           REGISTERS_5_0_port);
   REGISTERS_reg_6_31_inst : DLH_X1 port map( G => n231, D => n328_port, Q => 
                           REGISTERS_6_31_port);
   REGISTERS_reg_6_30_inst : DLH_X1 port map( G => n231, D => n332_port, Q => 
                           REGISTERS_6_30_port);
   REGISTERS_reg_6_29_inst : DLH_X1 port map( G => n230, D => n336_port, Q => 
                           REGISTERS_6_29_port);
   REGISTERS_reg_6_28_inst : DLH_X1 port map( G => n230, D => n340_port, Q => 
                           REGISTERS_6_28_port);
   REGISTERS_reg_6_27_inst : DLH_X1 port map( G => n230, D => n344_port, Q => 
                           REGISTERS_6_27_port);
   REGISTERS_reg_6_26_inst : DLH_X1 port map( G => n230, D => n348_port, Q => 
                           REGISTERS_6_26_port);
   REGISTERS_reg_6_25_inst : DLH_X1 port map( G => n230, D => n352_port, Q => 
                           REGISTERS_6_25_port);
   REGISTERS_reg_6_24_inst : DLH_X1 port map( G => n230, D => n356_port, Q => 
                           REGISTERS_6_24_port);
   REGISTERS_reg_6_23_inst : DLH_X1 port map( G => n230, D => n360_port, Q => 
                           REGISTERS_6_23_port);
   REGISTERS_reg_6_22_inst : DLH_X1 port map( G => n230, D => n364_port, Q => 
                           REGISTERS_6_22_port);
   REGISTERS_reg_6_21_inst : DLH_X1 port map( G => n230, D => n368_port, Q => 
                           REGISTERS_6_21_port);
   REGISTERS_reg_6_20_inst : DLH_X1 port map( G => n230, D => n372_port, Q => 
                           REGISTERS_6_20_port);
   REGISTERS_reg_6_19_inst : DLH_X1 port map( G => n229, D => n376_port, Q => 
                           REGISTERS_6_19_port);
   REGISTERS_reg_6_18_inst : DLH_X1 port map( G => n229, D => n380_port, Q => 
                           REGISTERS_6_18_port);
   REGISTERS_reg_6_17_inst : DLH_X1 port map( G => n229, D => n384_port, Q => 
                           REGISTERS_6_17_port);
   REGISTERS_reg_6_16_inst : DLH_X1 port map( G => n229, D => n388_port, Q => 
                           REGISTERS_6_16_port);
   REGISTERS_reg_6_15_inst : DLH_X1 port map( G => n229, D => n392_port, Q => 
                           REGISTERS_6_15_port);
   REGISTERS_reg_6_14_inst : DLH_X1 port map( G => n229, D => n396_port, Q => 
                           REGISTERS_6_14_port);
   REGISTERS_reg_6_13_inst : DLH_X1 port map( G => n229, D => n400_port, Q => 
                           REGISTERS_6_13_port);
   REGISTERS_reg_6_12_inst : DLH_X1 port map( G => n229, D => n404_port, Q => 
                           REGISTERS_6_12_port);
   REGISTERS_reg_6_11_inst : DLH_X1 port map( G => n229, D => n408_port, Q => 
                           REGISTERS_6_11_port);
   REGISTERS_reg_6_10_inst : DLH_X1 port map( G => n229, D => n412_port, Q => 
                           REGISTERS_6_10_port);
   REGISTERS_reg_6_9_inst : DLH_X1 port map( G => n228, D => n416_port, Q => 
                           REGISTERS_6_9_port);
   REGISTERS_reg_6_8_inst : DLH_X1 port map( G => n228, D => n420_port, Q => 
                           REGISTERS_6_8_port);
   REGISTERS_reg_6_7_inst : DLH_X1 port map( G => n228, D => n424_port, Q => 
                           REGISTERS_6_7_port);
   REGISTERS_reg_6_6_inst : DLH_X1 port map( G => n228, D => n428_port, Q => 
                           REGISTERS_6_6_port);
   REGISTERS_reg_6_5_inst : DLH_X1 port map( G => n228, D => n432_port, Q => 
                           REGISTERS_6_5_port);
   REGISTERS_reg_6_4_inst : DLH_X1 port map( G => n228, D => n436_port, Q => 
                           REGISTERS_6_4_port);
   REGISTERS_reg_6_3_inst : DLH_X1 port map( G => n228, D => n440_port, Q => 
                           REGISTERS_6_3_port);
   REGISTERS_reg_6_2_inst : DLH_X1 port map( G => n228, D => n444, Q => 
                           REGISTERS_6_2_port);
   REGISTERS_reg_6_1_inst : DLH_X1 port map( G => n228, D => n448, Q => 
                           REGISTERS_6_1_port);
   REGISTERS_reg_6_0_inst : DLH_X1 port map( G => n228, D => n452, Q => 
                           REGISTERS_6_0_port);
   REGISTERS_reg_7_31_inst : DLH_X1 port map( G => n235, D => n328_port, Q => 
                           REGISTERS_7_31_port);
   REGISTERS_reg_7_30_inst : DLH_X1 port map( G => n235, D => n332_port, Q => 
                           REGISTERS_7_30_port);
   REGISTERS_reg_7_29_inst : DLH_X1 port map( G => n234, D => n336_port, Q => 
                           REGISTERS_7_29_port);
   REGISTERS_reg_7_28_inst : DLH_X1 port map( G => n234, D => n340_port, Q => 
                           REGISTERS_7_28_port);
   REGISTERS_reg_7_27_inst : DLH_X1 port map( G => n234, D => n344_port, Q => 
                           REGISTERS_7_27_port);
   REGISTERS_reg_7_26_inst : DLH_X1 port map( G => n234, D => n348_port, Q => 
                           REGISTERS_7_26_port);
   REGISTERS_reg_7_25_inst : DLH_X1 port map( G => n234, D => n352_port, Q => 
                           REGISTERS_7_25_port);
   REGISTERS_reg_7_24_inst : DLH_X1 port map( G => n234, D => n356_port, Q => 
                           REGISTERS_7_24_port);
   REGISTERS_reg_7_23_inst : DLH_X1 port map( G => n234, D => n360_port, Q => 
                           REGISTERS_7_23_port);
   REGISTERS_reg_7_22_inst : DLH_X1 port map( G => n234, D => n364_port, Q => 
                           REGISTERS_7_22_port);
   REGISTERS_reg_7_21_inst : DLH_X1 port map( G => n234, D => n368_port, Q => 
                           REGISTERS_7_21_port);
   REGISTERS_reg_7_20_inst : DLH_X1 port map( G => n234, D => n372_port, Q => 
                           REGISTERS_7_20_port);
   REGISTERS_reg_7_19_inst : DLH_X1 port map( G => n233, D => n376_port, Q => 
                           REGISTERS_7_19_port);
   REGISTERS_reg_7_18_inst : DLH_X1 port map( G => n233, D => n380_port, Q => 
                           REGISTERS_7_18_port);
   REGISTERS_reg_7_17_inst : DLH_X1 port map( G => n233, D => n384_port, Q => 
                           REGISTERS_7_17_port);
   REGISTERS_reg_7_16_inst : DLH_X1 port map( G => n233, D => n388_port, Q => 
                           REGISTERS_7_16_port);
   REGISTERS_reg_7_15_inst : DLH_X1 port map( G => n233, D => n392_port, Q => 
                           REGISTERS_7_15_port);
   REGISTERS_reg_7_14_inst : DLH_X1 port map( G => n233, D => n396_port, Q => 
                           REGISTERS_7_14_port);
   REGISTERS_reg_7_13_inst : DLH_X1 port map( G => n233, D => n400_port, Q => 
                           REGISTERS_7_13_port);
   REGISTERS_reg_7_12_inst : DLH_X1 port map( G => n233, D => n404_port, Q => 
                           REGISTERS_7_12_port);
   REGISTERS_reg_7_11_inst : DLH_X1 port map( G => n233, D => n408_port, Q => 
                           REGISTERS_7_11_port);
   REGISTERS_reg_7_10_inst : DLH_X1 port map( G => n233, D => n412_port, Q => 
                           REGISTERS_7_10_port);
   REGISTERS_reg_7_9_inst : DLH_X1 port map( G => n232, D => n416_port, Q => 
                           REGISTERS_7_9_port);
   REGISTERS_reg_7_8_inst : DLH_X1 port map( G => n232, D => n420_port, Q => 
                           REGISTERS_7_8_port);
   REGISTERS_reg_7_7_inst : DLH_X1 port map( G => n232, D => n424_port, Q => 
                           REGISTERS_7_7_port);
   REGISTERS_reg_7_6_inst : DLH_X1 port map( G => n232, D => n428_port, Q => 
                           REGISTERS_7_6_port);
   REGISTERS_reg_7_5_inst : DLH_X1 port map( G => n232, D => n432_port, Q => 
                           REGISTERS_7_5_port);
   REGISTERS_reg_7_4_inst : DLH_X1 port map( G => n232, D => n436_port, Q => 
                           REGISTERS_7_4_port);
   REGISTERS_reg_7_3_inst : DLH_X1 port map( G => n232, D => n440_port, Q => 
                           REGISTERS_7_3_port);
   REGISTERS_reg_7_2_inst : DLH_X1 port map( G => n232, D => n444, Q => 
                           REGISTERS_7_2_port);
   REGISTERS_reg_7_1_inst : DLH_X1 port map( G => n232, D => n448, Q => 
                           REGISTERS_7_1_port);
   REGISTERS_reg_7_0_inst : DLH_X1 port map( G => n232, D => n452, Q => 
                           REGISTERS_7_0_port);
   REGISTERS_reg_8_31_inst : DLH_X1 port map( G => n239, D => n328_port, Q => 
                           REGISTERS_8_31_port);
   REGISTERS_reg_8_30_inst : DLH_X1 port map( G => n239, D => n332_port, Q => 
                           REGISTERS_8_30_port);
   REGISTERS_reg_8_29_inst : DLH_X1 port map( G => n238, D => n336_port, Q => 
                           REGISTERS_8_29_port);
   REGISTERS_reg_8_28_inst : DLH_X1 port map( G => n238, D => n340_port, Q => 
                           REGISTERS_8_28_port);
   REGISTERS_reg_8_27_inst : DLH_X1 port map( G => n238, D => n344_port, Q => 
                           REGISTERS_8_27_port);
   REGISTERS_reg_8_26_inst : DLH_X1 port map( G => n238, D => n348_port, Q => 
                           REGISTERS_8_26_port);
   REGISTERS_reg_8_25_inst : DLH_X1 port map( G => n238, D => n352_port, Q => 
                           REGISTERS_8_25_port);
   REGISTERS_reg_8_24_inst : DLH_X1 port map( G => n238, D => n356_port, Q => 
                           REGISTERS_8_24_port);
   REGISTERS_reg_8_23_inst : DLH_X1 port map( G => n238, D => n360_port, Q => 
                           REGISTERS_8_23_port);
   REGISTERS_reg_8_22_inst : DLH_X1 port map( G => n238, D => n364_port, Q => 
                           REGISTERS_8_22_port);
   REGISTERS_reg_8_21_inst : DLH_X1 port map( G => n238, D => n368_port, Q => 
                           REGISTERS_8_21_port);
   REGISTERS_reg_8_20_inst : DLH_X1 port map( G => n238, D => n372_port, Q => 
                           REGISTERS_8_20_port);
   REGISTERS_reg_8_19_inst : DLH_X1 port map( G => n237, D => n376_port, Q => 
                           REGISTERS_8_19_port);
   REGISTERS_reg_8_18_inst : DLH_X1 port map( G => n237, D => n380_port, Q => 
                           REGISTERS_8_18_port);
   REGISTERS_reg_8_17_inst : DLH_X1 port map( G => n237, D => n384_port, Q => 
                           REGISTERS_8_17_port);
   REGISTERS_reg_8_16_inst : DLH_X1 port map( G => n237, D => n388_port, Q => 
                           REGISTERS_8_16_port);
   REGISTERS_reg_8_15_inst : DLH_X1 port map( G => n237, D => n392_port, Q => 
                           REGISTERS_8_15_port);
   REGISTERS_reg_8_14_inst : DLH_X1 port map( G => n237, D => n396_port, Q => 
                           REGISTERS_8_14_port);
   REGISTERS_reg_8_13_inst : DLH_X1 port map( G => n237, D => n400_port, Q => 
                           REGISTERS_8_13_port);
   REGISTERS_reg_8_12_inst : DLH_X1 port map( G => n237, D => n404_port, Q => 
                           REGISTERS_8_12_port);
   REGISTERS_reg_8_11_inst : DLH_X1 port map( G => n237, D => n408_port, Q => 
                           REGISTERS_8_11_port);
   REGISTERS_reg_8_10_inst : DLH_X1 port map( G => n237, D => n412_port, Q => 
                           REGISTERS_8_10_port);
   REGISTERS_reg_8_9_inst : DLH_X1 port map( G => n236, D => n416_port, Q => 
                           REGISTERS_8_9_port);
   REGISTERS_reg_8_8_inst : DLH_X1 port map( G => n236, D => n420_port, Q => 
                           REGISTERS_8_8_port);
   REGISTERS_reg_8_7_inst : DLH_X1 port map( G => n236, D => n424_port, Q => 
                           REGISTERS_8_7_port);
   REGISTERS_reg_8_6_inst : DLH_X1 port map( G => n236, D => n428_port, Q => 
                           REGISTERS_8_6_port);
   REGISTERS_reg_8_5_inst : DLH_X1 port map( G => n236, D => n432_port, Q => 
                           REGISTERS_8_5_port);
   REGISTERS_reg_8_4_inst : DLH_X1 port map( G => n236, D => n436_port, Q => 
                           REGISTERS_8_4_port);
   REGISTERS_reg_8_3_inst : DLH_X1 port map( G => n236, D => n440_port, Q => 
                           REGISTERS_8_3_port);
   REGISTERS_reg_8_2_inst : DLH_X1 port map( G => n236, D => n444, Q => 
                           REGISTERS_8_2_port);
   REGISTERS_reg_8_1_inst : DLH_X1 port map( G => n236, D => n448, Q => 
                           REGISTERS_8_1_port);
   REGISTERS_reg_8_0_inst : DLH_X1 port map( G => n236, D => n452, Q => 
                           REGISTERS_8_0_port);
   REGISTERS_reg_9_31_inst : DLH_X1 port map( G => n243, D => n328_port, Q => 
                           REGISTERS_9_31_port);
   REGISTERS_reg_9_30_inst : DLH_X1 port map( G => n243, D => n332_port, Q => 
                           REGISTERS_9_30_port);
   REGISTERS_reg_9_29_inst : DLH_X1 port map( G => n242, D => n336_port, Q => 
                           REGISTERS_9_29_port);
   REGISTERS_reg_9_28_inst : DLH_X1 port map( G => n242, D => n340_port, Q => 
                           REGISTERS_9_28_port);
   REGISTERS_reg_9_27_inst : DLH_X1 port map( G => n242, D => n344_port, Q => 
                           REGISTERS_9_27_port);
   REGISTERS_reg_9_26_inst : DLH_X1 port map( G => n242, D => n348_port, Q => 
                           REGISTERS_9_26_port);
   REGISTERS_reg_9_25_inst : DLH_X1 port map( G => n242, D => n352_port, Q => 
                           REGISTERS_9_25_port);
   REGISTERS_reg_9_24_inst : DLH_X1 port map( G => n242, D => n356_port, Q => 
                           REGISTERS_9_24_port);
   REGISTERS_reg_9_23_inst : DLH_X1 port map( G => n242, D => n360_port, Q => 
                           REGISTERS_9_23_port);
   REGISTERS_reg_9_22_inst : DLH_X1 port map( G => n242, D => n364_port, Q => 
                           REGISTERS_9_22_port);
   REGISTERS_reg_9_21_inst : DLH_X1 port map( G => n242, D => n368_port, Q => 
                           REGISTERS_9_21_port);
   REGISTERS_reg_9_20_inst : DLH_X1 port map( G => n242, D => n372_port, Q => 
                           REGISTERS_9_20_port);
   REGISTERS_reg_9_19_inst : DLH_X1 port map( G => n241, D => n376_port, Q => 
                           REGISTERS_9_19_port);
   REGISTERS_reg_9_18_inst : DLH_X1 port map( G => n241, D => n380_port, Q => 
                           REGISTERS_9_18_port);
   REGISTERS_reg_9_17_inst : DLH_X1 port map( G => n241, D => n384_port, Q => 
                           REGISTERS_9_17_port);
   REGISTERS_reg_9_16_inst : DLH_X1 port map( G => n241, D => n388_port, Q => 
                           REGISTERS_9_16_port);
   REGISTERS_reg_9_15_inst : DLH_X1 port map( G => n241, D => n392_port, Q => 
                           REGISTERS_9_15_port);
   REGISTERS_reg_9_14_inst : DLH_X1 port map( G => n241, D => n396_port, Q => 
                           REGISTERS_9_14_port);
   REGISTERS_reg_9_13_inst : DLH_X1 port map( G => n241, D => n400_port, Q => 
                           REGISTERS_9_13_port);
   REGISTERS_reg_9_12_inst : DLH_X1 port map( G => n241, D => n404_port, Q => 
                           REGISTERS_9_12_port);
   REGISTERS_reg_9_11_inst : DLH_X1 port map( G => n241, D => n408_port, Q => 
                           REGISTERS_9_11_port);
   REGISTERS_reg_9_10_inst : DLH_X1 port map( G => n241, D => n412_port, Q => 
                           REGISTERS_9_10_port);
   REGISTERS_reg_9_9_inst : DLH_X1 port map( G => n240, D => n416_port, Q => 
                           REGISTERS_9_9_port);
   REGISTERS_reg_9_8_inst : DLH_X1 port map( G => n240, D => n420_port, Q => 
                           REGISTERS_9_8_port);
   REGISTERS_reg_9_7_inst : DLH_X1 port map( G => n240, D => n424_port, Q => 
                           REGISTERS_9_7_port);
   REGISTERS_reg_9_6_inst : DLH_X1 port map( G => n240, D => n428_port, Q => 
                           REGISTERS_9_6_port);
   REGISTERS_reg_9_5_inst : DLH_X1 port map( G => n240, D => n432_port, Q => 
                           REGISTERS_9_5_port);
   REGISTERS_reg_9_4_inst : DLH_X1 port map( G => n240, D => n436_port, Q => 
                           REGISTERS_9_4_port);
   REGISTERS_reg_9_3_inst : DLH_X1 port map( G => n240, D => n440_port, Q => 
                           REGISTERS_9_3_port);
   REGISTERS_reg_9_2_inst : DLH_X1 port map( G => n240, D => n444, Q => 
                           REGISTERS_9_2_port);
   REGISTERS_reg_9_1_inst : DLH_X1 port map( G => n240, D => n448, Q => 
                           REGISTERS_9_1_port);
   REGISTERS_reg_9_0_inst : DLH_X1 port map( G => n240, D => n452, Q => 
                           REGISTERS_9_0_port);
   REGISTERS_reg_10_31_inst : DLH_X1 port map( G => n247, D => n329_port, Q => 
                           REGISTERS_10_31_port);
   REGISTERS_reg_10_30_inst : DLH_X1 port map( G => n247, D => n333_port, Q => 
                           REGISTERS_10_30_port);
   REGISTERS_reg_10_29_inst : DLH_X1 port map( G => n246, D => n337_port, Q => 
                           REGISTERS_10_29_port);
   REGISTERS_reg_10_28_inst : DLH_X1 port map( G => n246, D => n341_port, Q => 
                           REGISTERS_10_28_port);
   REGISTERS_reg_10_27_inst : DLH_X1 port map( G => n246, D => n345_port, Q => 
                           REGISTERS_10_27_port);
   REGISTERS_reg_10_26_inst : DLH_X1 port map( G => n246, D => n349_port, Q => 
                           REGISTERS_10_26_port);
   REGISTERS_reg_10_25_inst : DLH_X1 port map( G => n246, D => n353_port, Q => 
                           REGISTERS_10_25_port);
   REGISTERS_reg_10_24_inst : DLH_X1 port map( G => n246, D => n357_port, Q => 
                           REGISTERS_10_24_port);
   REGISTERS_reg_10_23_inst : DLH_X1 port map( G => n246, D => n361_port, Q => 
                           REGISTERS_10_23_port);
   REGISTERS_reg_10_22_inst : DLH_X1 port map( G => n246, D => n365_port, Q => 
                           REGISTERS_10_22_port);
   REGISTERS_reg_10_21_inst : DLH_X1 port map( G => n246, D => n369_port, Q => 
                           REGISTERS_10_21_port);
   REGISTERS_reg_10_20_inst : DLH_X1 port map( G => n246, D => n373_port, Q => 
                           REGISTERS_10_20_port);
   REGISTERS_reg_10_19_inst : DLH_X1 port map( G => n245, D => n377_port, Q => 
                           REGISTERS_10_19_port);
   REGISTERS_reg_10_18_inst : DLH_X1 port map( G => n245, D => n381_port, Q => 
                           REGISTERS_10_18_port);
   REGISTERS_reg_10_17_inst : DLH_X1 port map( G => n245, D => n385_port, Q => 
                           REGISTERS_10_17_port);
   REGISTERS_reg_10_16_inst : DLH_X1 port map( G => n245, D => n389_port, Q => 
                           REGISTERS_10_16_port);
   REGISTERS_reg_10_15_inst : DLH_X1 port map( G => n245, D => n393_port, Q => 
                           REGISTERS_10_15_port);
   REGISTERS_reg_10_14_inst : DLH_X1 port map( G => n245, D => n397_port, Q => 
                           REGISTERS_10_14_port);
   REGISTERS_reg_10_13_inst : DLH_X1 port map( G => n245, D => n401_port, Q => 
                           REGISTERS_10_13_port);
   REGISTERS_reg_10_12_inst : DLH_X1 port map( G => n245, D => n405_port, Q => 
                           REGISTERS_10_12_port);
   REGISTERS_reg_10_11_inst : DLH_X1 port map( G => n245, D => n409_port, Q => 
                           REGISTERS_10_11_port);
   REGISTERS_reg_10_10_inst : DLH_X1 port map( G => n245, D => n413_port, Q => 
                           REGISTERS_10_10_port);
   REGISTERS_reg_10_9_inst : DLH_X1 port map( G => n244, D => n417_port, Q => 
                           REGISTERS_10_9_port);
   REGISTERS_reg_10_8_inst : DLH_X1 port map( G => n244, D => n421_port, Q => 
                           REGISTERS_10_8_port);
   REGISTERS_reg_10_7_inst : DLH_X1 port map( G => n244, D => n425_port, Q => 
                           REGISTERS_10_7_port);
   REGISTERS_reg_10_6_inst : DLH_X1 port map( G => n244, D => n429_port, Q => 
                           REGISTERS_10_6_port);
   REGISTERS_reg_10_5_inst : DLH_X1 port map( G => n244, D => n433_port, Q => 
                           REGISTERS_10_5_port);
   REGISTERS_reg_10_4_inst : DLH_X1 port map( G => n244, D => n437_port, Q => 
                           REGISTERS_10_4_port);
   REGISTERS_reg_10_3_inst : DLH_X1 port map( G => n244, D => n441_port, Q => 
                           REGISTERS_10_3_port);
   REGISTERS_reg_10_2_inst : DLH_X1 port map( G => n244, D => n445, Q => 
                           REGISTERS_10_2_port);
   REGISTERS_reg_10_1_inst : DLH_X1 port map( G => n244, D => n449, Q => 
                           REGISTERS_10_1_port);
   REGISTERS_reg_10_0_inst : DLH_X1 port map( G => n244, D => n453, Q => 
                           REGISTERS_10_0_port);
   REGISTERS_reg_11_31_inst : DLH_X1 port map( G => n251, D => n329_port, Q => 
                           REGISTERS_11_31_port);
   REGISTERS_reg_11_30_inst : DLH_X1 port map( G => n251, D => n333_port, Q => 
                           REGISTERS_11_30_port);
   REGISTERS_reg_11_29_inst : DLH_X1 port map( G => n250, D => n337_port, Q => 
                           REGISTERS_11_29_port);
   REGISTERS_reg_11_28_inst : DLH_X1 port map( G => n250, D => n341_port, Q => 
                           REGISTERS_11_28_port);
   REGISTERS_reg_11_27_inst : DLH_X1 port map( G => n250, D => n345_port, Q => 
                           REGISTERS_11_27_port);
   REGISTERS_reg_11_26_inst : DLH_X1 port map( G => n250, D => n349_port, Q => 
                           REGISTERS_11_26_port);
   REGISTERS_reg_11_25_inst : DLH_X1 port map( G => n250, D => n353_port, Q => 
                           REGISTERS_11_25_port);
   REGISTERS_reg_11_24_inst : DLH_X1 port map( G => n250, D => n357_port, Q => 
                           REGISTERS_11_24_port);
   REGISTERS_reg_11_23_inst : DLH_X1 port map( G => n250, D => n361_port, Q => 
                           REGISTERS_11_23_port);
   REGISTERS_reg_11_22_inst : DLH_X1 port map( G => n250, D => n365_port, Q => 
                           REGISTERS_11_22_port);
   REGISTERS_reg_11_21_inst : DLH_X1 port map( G => n250, D => n369_port, Q => 
                           REGISTERS_11_21_port);
   REGISTERS_reg_11_20_inst : DLH_X1 port map( G => n250, D => n373_port, Q => 
                           REGISTERS_11_20_port);
   REGISTERS_reg_11_19_inst : DLH_X1 port map( G => n249, D => n377_port, Q => 
                           REGISTERS_11_19_port);
   REGISTERS_reg_11_18_inst : DLH_X1 port map( G => n249, D => n381_port, Q => 
                           REGISTERS_11_18_port);
   REGISTERS_reg_11_17_inst : DLH_X1 port map( G => n249, D => n385_port, Q => 
                           REGISTERS_11_17_port);
   REGISTERS_reg_11_16_inst : DLH_X1 port map( G => n249, D => n389_port, Q => 
                           REGISTERS_11_16_port);
   REGISTERS_reg_11_15_inst : DLH_X1 port map( G => n249, D => n393_port, Q => 
                           REGISTERS_11_15_port);
   REGISTERS_reg_11_14_inst : DLH_X1 port map( G => n249, D => n397_port, Q => 
                           REGISTERS_11_14_port);
   REGISTERS_reg_11_13_inst : DLH_X1 port map( G => n249, D => n401_port, Q => 
                           REGISTERS_11_13_port);
   REGISTERS_reg_11_12_inst : DLH_X1 port map( G => n249, D => n405_port, Q => 
                           REGISTERS_11_12_port);
   REGISTERS_reg_11_11_inst : DLH_X1 port map( G => n249, D => n409_port, Q => 
                           REGISTERS_11_11_port);
   REGISTERS_reg_11_10_inst : DLH_X1 port map( G => n249, D => n413_port, Q => 
                           REGISTERS_11_10_port);
   REGISTERS_reg_11_9_inst : DLH_X1 port map( G => n248, D => n417_port, Q => 
                           REGISTERS_11_9_port);
   REGISTERS_reg_11_8_inst : DLH_X1 port map( G => n248, D => n421_port, Q => 
                           REGISTERS_11_8_port);
   REGISTERS_reg_11_7_inst : DLH_X1 port map( G => n248, D => n425_port, Q => 
                           REGISTERS_11_7_port);
   REGISTERS_reg_11_6_inst : DLH_X1 port map( G => n248, D => n429_port, Q => 
                           REGISTERS_11_6_port);
   REGISTERS_reg_11_5_inst : DLH_X1 port map( G => n248, D => n433_port, Q => 
                           REGISTERS_11_5_port);
   REGISTERS_reg_11_4_inst : DLH_X1 port map( G => n248, D => n437_port, Q => 
                           REGISTERS_11_4_port);
   REGISTERS_reg_11_3_inst : DLH_X1 port map( G => n248, D => n441_port, Q => 
                           REGISTERS_11_3_port);
   REGISTERS_reg_11_2_inst : DLH_X1 port map( G => n248, D => n445, Q => 
                           REGISTERS_11_2_port);
   REGISTERS_reg_11_1_inst : DLH_X1 port map( G => n248, D => n449, Q => 
                           REGISTERS_11_1_port);
   REGISTERS_reg_11_0_inst : DLH_X1 port map( G => n248, D => n453, Q => 
                           REGISTERS_11_0_port);
   REGISTERS_reg_12_31_inst : DLH_X1 port map( G => n255, D => n329_port, Q => 
                           REGISTERS_12_31_port);
   REGISTERS_reg_12_30_inst : DLH_X1 port map( G => n255, D => n333_port, Q => 
                           REGISTERS_12_30_port);
   REGISTERS_reg_12_29_inst : DLH_X1 port map( G => n254, D => n337_port, Q => 
                           REGISTERS_12_29_port);
   REGISTERS_reg_12_28_inst : DLH_X1 port map( G => n254, D => n341_port, Q => 
                           REGISTERS_12_28_port);
   REGISTERS_reg_12_27_inst : DLH_X1 port map( G => n254, D => n345_port, Q => 
                           REGISTERS_12_27_port);
   REGISTERS_reg_12_26_inst : DLH_X1 port map( G => n254, D => n349_port, Q => 
                           REGISTERS_12_26_port);
   REGISTERS_reg_12_25_inst : DLH_X1 port map( G => n254, D => n353_port, Q => 
                           REGISTERS_12_25_port);
   REGISTERS_reg_12_24_inst : DLH_X1 port map( G => n254, D => n357_port, Q => 
                           REGISTERS_12_24_port);
   REGISTERS_reg_12_23_inst : DLH_X1 port map( G => n254, D => n361_port, Q => 
                           REGISTERS_12_23_port);
   REGISTERS_reg_12_22_inst : DLH_X1 port map( G => n254, D => n365_port, Q => 
                           REGISTERS_12_22_port);
   REGISTERS_reg_12_21_inst : DLH_X1 port map( G => n254, D => n369_port, Q => 
                           REGISTERS_12_21_port);
   REGISTERS_reg_12_20_inst : DLH_X1 port map( G => n254, D => n373_port, Q => 
                           REGISTERS_12_20_port);
   REGISTERS_reg_12_19_inst : DLH_X1 port map( G => n253, D => n377_port, Q => 
                           REGISTERS_12_19_port);
   REGISTERS_reg_12_18_inst : DLH_X1 port map( G => n253, D => n381_port, Q => 
                           REGISTERS_12_18_port);
   REGISTERS_reg_12_17_inst : DLH_X1 port map( G => n253, D => n385_port, Q => 
                           REGISTERS_12_17_port);
   REGISTERS_reg_12_16_inst : DLH_X1 port map( G => n253, D => n389_port, Q => 
                           REGISTERS_12_16_port);
   REGISTERS_reg_12_15_inst : DLH_X1 port map( G => n253, D => n393_port, Q => 
                           REGISTERS_12_15_port);
   REGISTERS_reg_12_14_inst : DLH_X1 port map( G => n253, D => n397_port, Q => 
                           REGISTERS_12_14_port);
   REGISTERS_reg_12_13_inst : DLH_X1 port map( G => n253, D => n401_port, Q => 
                           REGISTERS_12_13_port);
   REGISTERS_reg_12_12_inst : DLH_X1 port map( G => n253, D => n405_port, Q => 
                           REGISTERS_12_12_port);
   REGISTERS_reg_12_11_inst : DLH_X1 port map( G => n253, D => n409_port, Q => 
                           REGISTERS_12_11_port);
   REGISTERS_reg_12_10_inst : DLH_X1 port map( G => n253, D => n413_port, Q => 
                           REGISTERS_12_10_port);
   REGISTERS_reg_12_9_inst : DLH_X1 port map( G => n252, D => n417_port, Q => 
                           REGISTERS_12_9_port);
   REGISTERS_reg_12_8_inst : DLH_X1 port map( G => n252, D => n421_port, Q => 
                           REGISTERS_12_8_port);
   REGISTERS_reg_12_7_inst : DLH_X1 port map( G => n252, D => n425_port, Q => 
                           REGISTERS_12_7_port);
   REGISTERS_reg_12_6_inst : DLH_X1 port map( G => n252, D => n429_port, Q => 
                           REGISTERS_12_6_port);
   REGISTERS_reg_12_5_inst : DLH_X1 port map( G => n252, D => n433_port, Q => 
                           REGISTERS_12_5_port);
   REGISTERS_reg_12_4_inst : DLH_X1 port map( G => n252, D => n437_port, Q => 
                           REGISTERS_12_4_port);
   REGISTERS_reg_12_3_inst : DLH_X1 port map( G => n252, D => n441_port, Q => 
                           REGISTERS_12_3_port);
   REGISTERS_reg_12_2_inst : DLH_X1 port map( G => n252, D => n445, Q => 
                           REGISTERS_12_2_port);
   REGISTERS_reg_12_1_inst : DLH_X1 port map( G => n252, D => n449, Q => 
                           REGISTERS_12_1_port);
   REGISTERS_reg_12_0_inst : DLH_X1 port map( G => n252, D => n453, Q => 
                           REGISTERS_12_0_port);
   REGISTERS_reg_13_31_inst : DLH_X1 port map( G => n259, D => n329_port, Q => 
                           REGISTERS_13_31_port);
   REGISTERS_reg_13_30_inst : DLH_X1 port map( G => n259, D => n333_port, Q => 
                           REGISTERS_13_30_port);
   REGISTERS_reg_13_29_inst : DLH_X1 port map( G => n258, D => n337_port, Q => 
                           REGISTERS_13_29_port);
   REGISTERS_reg_13_28_inst : DLH_X1 port map( G => n258, D => n341_port, Q => 
                           REGISTERS_13_28_port);
   REGISTERS_reg_13_27_inst : DLH_X1 port map( G => n258, D => n345_port, Q => 
                           REGISTERS_13_27_port);
   REGISTERS_reg_13_26_inst : DLH_X1 port map( G => n258, D => n349_port, Q => 
                           REGISTERS_13_26_port);
   REGISTERS_reg_13_25_inst : DLH_X1 port map( G => n258, D => n353_port, Q => 
                           REGISTERS_13_25_port);
   REGISTERS_reg_13_24_inst : DLH_X1 port map( G => n258, D => n357_port, Q => 
                           REGISTERS_13_24_port);
   REGISTERS_reg_13_23_inst : DLH_X1 port map( G => n258, D => n361_port, Q => 
                           REGISTERS_13_23_port);
   REGISTERS_reg_13_22_inst : DLH_X1 port map( G => n258, D => n365_port, Q => 
                           REGISTERS_13_22_port);
   REGISTERS_reg_13_21_inst : DLH_X1 port map( G => n258, D => n369_port, Q => 
                           REGISTERS_13_21_port);
   REGISTERS_reg_13_20_inst : DLH_X1 port map( G => n258, D => n373_port, Q => 
                           REGISTERS_13_20_port);
   REGISTERS_reg_13_19_inst : DLH_X1 port map( G => n257, D => n377_port, Q => 
                           REGISTERS_13_19_port);
   REGISTERS_reg_13_18_inst : DLH_X1 port map( G => n257, D => n381_port, Q => 
                           REGISTERS_13_18_port);
   REGISTERS_reg_13_17_inst : DLH_X1 port map( G => n257, D => n385_port, Q => 
                           REGISTERS_13_17_port);
   REGISTERS_reg_13_16_inst : DLH_X1 port map( G => n257, D => n389_port, Q => 
                           REGISTERS_13_16_port);
   REGISTERS_reg_13_15_inst : DLH_X1 port map( G => n257, D => n393_port, Q => 
                           REGISTERS_13_15_port);
   REGISTERS_reg_13_14_inst : DLH_X1 port map( G => n257, D => n397_port, Q => 
                           REGISTERS_13_14_port);
   REGISTERS_reg_13_13_inst : DLH_X1 port map( G => n257, D => n401_port, Q => 
                           REGISTERS_13_13_port);
   REGISTERS_reg_13_12_inst : DLH_X1 port map( G => n257, D => n405_port, Q => 
                           REGISTERS_13_12_port);
   REGISTERS_reg_13_11_inst : DLH_X1 port map( G => n257, D => n409_port, Q => 
                           REGISTERS_13_11_port);
   REGISTERS_reg_13_10_inst : DLH_X1 port map( G => n257, D => n413_port, Q => 
                           REGISTERS_13_10_port);
   REGISTERS_reg_13_9_inst : DLH_X1 port map( G => n256, D => n417_port, Q => 
                           REGISTERS_13_9_port);
   REGISTERS_reg_13_8_inst : DLH_X1 port map( G => n256, D => n421_port, Q => 
                           REGISTERS_13_8_port);
   REGISTERS_reg_13_7_inst : DLH_X1 port map( G => n256, D => n425_port, Q => 
                           REGISTERS_13_7_port);
   REGISTERS_reg_13_6_inst : DLH_X1 port map( G => n256, D => n429_port, Q => 
                           REGISTERS_13_6_port);
   REGISTERS_reg_13_5_inst : DLH_X1 port map( G => n256, D => n433_port, Q => 
                           REGISTERS_13_5_port);
   REGISTERS_reg_13_4_inst : DLH_X1 port map( G => n256, D => n437_port, Q => 
                           REGISTERS_13_4_port);
   REGISTERS_reg_13_3_inst : DLH_X1 port map( G => n256, D => n441_port, Q => 
                           REGISTERS_13_3_port);
   REGISTERS_reg_13_2_inst : DLH_X1 port map( G => n256, D => n445, Q => 
                           REGISTERS_13_2_port);
   REGISTERS_reg_13_1_inst : DLH_X1 port map( G => n256, D => n449, Q => 
                           REGISTERS_13_1_port);
   REGISTERS_reg_13_0_inst : DLH_X1 port map( G => n256, D => n453, Q => 
                           REGISTERS_13_0_port);
   REGISTERS_reg_14_31_inst : DLH_X1 port map( G => n263, D => n329_port, Q => 
                           REGISTERS_14_31_port);
   REGISTERS_reg_14_30_inst : DLH_X1 port map( G => n263, D => n333_port, Q => 
                           REGISTERS_14_30_port);
   REGISTERS_reg_14_29_inst : DLH_X1 port map( G => n262, D => n337_port, Q => 
                           REGISTERS_14_29_port);
   REGISTERS_reg_14_28_inst : DLH_X1 port map( G => n262, D => n341_port, Q => 
                           REGISTERS_14_28_port);
   REGISTERS_reg_14_27_inst : DLH_X1 port map( G => n262, D => n345_port, Q => 
                           REGISTERS_14_27_port);
   REGISTERS_reg_14_26_inst : DLH_X1 port map( G => n262, D => n349_port, Q => 
                           REGISTERS_14_26_port);
   REGISTERS_reg_14_25_inst : DLH_X1 port map( G => n262, D => n353_port, Q => 
                           REGISTERS_14_25_port);
   REGISTERS_reg_14_24_inst : DLH_X1 port map( G => n262, D => n357_port, Q => 
                           REGISTERS_14_24_port);
   REGISTERS_reg_14_23_inst : DLH_X1 port map( G => n262, D => n361_port, Q => 
                           REGISTERS_14_23_port);
   REGISTERS_reg_14_22_inst : DLH_X1 port map( G => n262, D => n365_port, Q => 
                           REGISTERS_14_22_port);
   REGISTERS_reg_14_21_inst : DLH_X1 port map( G => n262, D => n369_port, Q => 
                           REGISTERS_14_21_port);
   REGISTERS_reg_14_20_inst : DLH_X1 port map( G => n262, D => n373_port, Q => 
                           REGISTERS_14_20_port);
   REGISTERS_reg_14_19_inst : DLH_X1 port map( G => n261, D => n377_port, Q => 
                           REGISTERS_14_19_port);
   REGISTERS_reg_14_18_inst : DLH_X1 port map( G => n261, D => n381_port, Q => 
                           REGISTERS_14_18_port);
   REGISTERS_reg_14_17_inst : DLH_X1 port map( G => n261, D => n385_port, Q => 
                           REGISTERS_14_17_port);
   REGISTERS_reg_14_16_inst : DLH_X1 port map( G => n261, D => n389_port, Q => 
                           REGISTERS_14_16_port);
   REGISTERS_reg_14_15_inst : DLH_X1 port map( G => n261, D => n393_port, Q => 
                           REGISTERS_14_15_port);
   REGISTERS_reg_14_14_inst : DLH_X1 port map( G => n261, D => n397_port, Q => 
                           REGISTERS_14_14_port);
   REGISTERS_reg_14_13_inst : DLH_X1 port map( G => n261, D => n401_port, Q => 
                           REGISTERS_14_13_port);
   REGISTERS_reg_14_12_inst : DLH_X1 port map( G => n261, D => n405_port, Q => 
                           REGISTERS_14_12_port);
   REGISTERS_reg_14_11_inst : DLH_X1 port map( G => n261, D => n409_port, Q => 
                           REGISTERS_14_11_port);
   REGISTERS_reg_14_10_inst : DLH_X1 port map( G => n261, D => n413_port, Q => 
                           REGISTERS_14_10_port);
   REGISTERS_reg_14_9_inst : DLH_X1 port map( G => n260, D => n417_port, Q => 
                           REGISTERS_14_9_port);
   REGISTERS_reg_14_8_inst : DLH_X1 port map( G => n260, D => n421_port, Q => 
                           REGISTERS_14_8_port);
   REGISTERS_reg_14_7_inst : DLH_X1 port map( G => n260, D => n425_port, Q => 
                           REGISTERS_14_7_port);
   REGISTERS_reg_14_6_inst : DLH_X1 port map( G => n260, D => n429_port, Q => 
                           REGISTERS_14_6_port);
   REGISTERS_reg_14_5_inst : DLH_X1 port map( G => n260, D => n433_port, Q => 
                           REGISTERS_14_5_port);
   REGISTERS_reg_14_4_inst : DLH_X1 port map( G => n260, D => n437_port, Q => 
                           REGISTERS_14_4_port);
   REGISTERS_reg_14_3_inst : DLH_X1 port map( G => n260, D => n441_port, Q => 
                           REGISTERS_14_3_port);
   REGISTERS_reg_14_2_inst : DLH_X1 port map( G => n260, D => n445, Q => 
                           REGISTERS_14_2_port);
   REGISTERS_reg_14_1_inst : DLH_X1 port map( G => n260, D => n449, Q => 
                           REGISTERS_14_1_port);
   REGISTERS_reg_14_0_inst : DLH_X1 port map( G => n260, D => n453, Q => 
                           REGISTERS_14_0_port);
   REGISTERS_reg_15_31_inst : DLH_X1 port map( G => n267, D => n329_port, Q => 
                           REGISTERS_15_31_port);
   REGISTERS_reg_15_30_inst : DLH_X1 port map( G => n267, D => n333_port, Q => 
                           REGISTERS_15_30_port);
   REGISTERS_reg_15_29_inst : DLH_X1 port map( G => n266, D => n337_port, Q => 
                           REGISTERS_15_29_port);
   REGISTERS_reg_15_28_inst : DLH_X1 port map( G => n266, D => n341_port, Q => 
                           REGISTERS_15_28_port);
   REGISTERS_reg_15_27_inst : DLH_X1 port map( G => n266, D => n345_port, Q => 
                           REGISTERS_15_27_port);
   REGISTERS_reg_15_26_inst : DLH_X1 port map( G => n266, D => n349_port, Q => 
                           REGISTERS_15_26_port);
   REGISTERS_reg_15_25_inst : DLH_X1 port map( G => n266, D => n353_port, Q => 
                           REGISTERS_15_25_port);
   REGISTERS_reg_15_24_inst : DLH_X1 port map( G => n266, D => n357_port, Q => 
                           REGISTERS_15_24_port);
   REGISTERS_reg_15_23_inst : DLH_X1 port map( G => n266, D => n361_port, Q => 
                           REGISTERS_15_23_port);
   REGISTERS_reg_15_22_inst : DLH_X1 port map( G => n266, D => n365_port, Q => 
                           REGISTERS_15_22_port);
   REGISTERS_reg_15_21_inst : DLH_X1 port map( G => n266, D => n369_port, Q => 
                           REGISTERS_15_21_port);
   REGISTERS_reg_15_20_inst : DLH_X1 port map( G => n266, D => n373_port, Q => 
                           REGISTERS_15_20_port);
   REGISTERS_reg_15_19_inst : DLH_X1 port map( G => n265, D => n377_port, Q => 
                           REGISTERS_15_19_port);
   REGISTERS_reg_15_18_inst : DLH_X1 port map( G => n265, D => n381_port, Q => 
                           REGISTERS_15_18_port);
   REGISTERS_reg_15_17_inst : DLH_X1 port map( G => n265, D => n385_port, Q => 
                           REGISTERS_15_17_port);
   REGISTERS_reg_15_16_inst : DLH_X1 port map( G => n265, D => n389_port, Q => 
                           REGISTERS_15_16_port);
   REGISTERS_reg_15_15_inst : DLH_X1 port map( G => n265, D => n393_port, Q => 
                           REGISTERS_15_15_port);
   REGISTERS_reg_15_14_inst : DLH_X1 port map( G => n265, D => n397_port, Q => 
                           REGISTERS_15_14_port);
   REGISTERS_reg_15_13_inst : DLH_X1 port map( G => n265, D => n401_port, Q => 
                           REGISTERS_15_13_port);
   REGISTERS_reg_15_12_inst : DLH_X1 port map( G => n265, D => n405_port, Q => 
                           REGISTERS_15_12_port);
   REGISTERS_reg_15_11_inst : DLH_X1 port map( G => n265, D => n409_port, Q => 
                           REGISTERS_15_11_port);
   REGISTERS_reg_15_10_inst : DLH_X1 port map( G => n265, D => n413_port, Q => 
                           REGISTERS_15_10_port);
   REGISTERS_reg_15_9_inst : DLH_X1 port map( G => n264, D => n417_port, Q => 
                           REGISTERS_15_9_port);
   REGISTERS_reg_15_8_inst : DLH_X1 port map( G => n264, D => n421_port, Q => 
                           REGISTERS_15_8_port);
   REGISTERS_reg_15_7_inst : DLH_X1 port map( G => n264, D => n425_port, Q => 
                           REGISTERS_15_7_port);
   REGISTERS_reg_15_6_inst : DLH_X1 port map( G => n264, D => n429_port, Q => 
                           REGISTERS_15_6_port);
   REGISTERS_reg_15_5_inst : DLH_X1 port map( G => n264, D => n433_port, Q => 
                           REGISTERS_15_5_port);
   REGISTERS_reg_15_4_inst : DLH_X1 port map( G => n264, D => n437_port, Q => 
                           REGISTERS_15_4_port);
   REGISTERS_reg_15_3_inst : DLH_X1 port map( G => n264, D => n441_port, Q => 
                           REGISTERS_15_3_port);
   REGISTERS_reg_15_2_inst : DLH_X1 port map( G => n264, D => n445, Q => 
                           REGISTERS_15_2_port);
   REGISTERS_reg_15_1_inst : DLH_X1 port map( G => n264, D => n449, Q => 
                           REGISTERS_15_1_port);
   REGISTERS_reg_15_0_inst : DLH_X1 port map( G => n264, D => n453, Q => 
                           REGISTERS_15_0_port);
   REGISTERS_reg_16_31_inst : DLH_X1 port map( G => n271, D => n329_port, Q => 
                           REGISTERS_16_31_port);
   REGISTERS_reg_16_30_inst : DLH_X1 port map( G => n271, D => n333_port, Q => 
                           REGISTERS_16_30_port);
   REGISTERS_reg_16_29_inst : DLH_X1 port map( G => n270, D => n337_port, Q => 
                           REGISTERS_16_29_port);
   REGISTERS_reg_16_28_inst : DLH_X1 port map( G => n270, D => n341_port, Q => 
                           REGISTERS_16_28_port);
   REGISTERS_reg_16_27_inst : DLH_X1 port map( G => n270, D => n345_port, Q => 
                           REGISTERS_16_27_port);
   REGISTERS_reg_16_26_inst : DLH_X1 port map( G => n270, D => n349_port, Q => 
                           REGISTERS_16_26_port);
   REGISTERS_reg_16_25_inst : DLH_X1 port map( G => n270, D => n353_port, Q => 
                           REGISTERS_16_25_port);
   REGISTERS_reg_16_24_inst : DLH_X1 port map( G => n270, D => n357_port, Q => 
                           REGISTERS_16_24_port);
   REGISTERS_reg_16_23_inst : DLH_X1 port map( G => n270, D => n361_port, Q => 
                           REGISTERS_16_23_port);
   REGISTERS_reg_16_22_inst : DLH_X1 port map( G => n270, D => n365_port, Q => 
                           REGISTERS_16_22_port);
   REGISTERS_reg_16_21_inst : DLH_X1 port map( G => n270, D => n369_port, Q => 
                           REGISTERS_16_21_port);
   REGISTERS_reg_16_20_inst : DLH_X1 port map( G => n270, D => n373_port, Q => 
                           REGISTERS_16_20_port);
   REGISTERS_reg_16_19_inst : DLH_X1 port map( G => n269, D => n377_port, Q => 
                           REGISTERS_16_19_port);
   REGISTERS_reg_16_18_inst : DLH_X1 port map( G => n269, D => n381_port, Q => 
                           REGISTERS_16_18_port);
   REGISTERS_reg_16_17_inst : DLH_X1 port map( G => n269, D => n385_port, Q => 
                           REGISTERS_16_17_port);
   REGISTERS_reg_16_16_inst : DLH_X1 port map( G => n269, D => n389_port, Q => 
                           REGISTERS_16_16_port);
   REGISTERS_reg_16_15_inst : DLH_X1 port map( G => n269, D => n393_port, Q => 
                           REGISTERS_16_15_port);
   REGISTERS_reg_16_14_inst : DLH_X1 port map( G => n269, D => n397_port, Q => 
                           REGISTERS_16_14_port);
   REGISTERS_reg_16_13_inst : DLH_X1 port map( G => n269, D => n401_port, Q => 
                           REGISTERS_16_13_port);
   REGISTERS_reg_16_12_inst : DLH_X1 port map( G => n269, D => n405_port, Q => 
                           REGISTERS_16_12_port);
   REGISTERS_reg_16_11_inst : DLH_X1 port map( G => n269, D => n409_port, Q => 
                           REGISTERS_16_11_port);
   REGISTERS_reg_16_10_inst : DLH_X1 port map( G => n269, D => n413_port, Q => 
                           REGISTERS_16_10_port);
   REGISTERS_reg_16_9_inst : DLH_X1 port map( G => n268, D => n417_port, Q => 
                           REGISTERS_16_9_port);
   REGISTERS_reg_16_8_inst : DLH_X1 port map( G => n268, D => n421_port, Q => 
                           REGISTERS_16_8_port);
   REGISTERS_reg_16_7_inst : DLH_X1 port map( G => n268, D => n425_port, Q => 
                           REGISTERS_16_7_port);
   REGISTERS_reg_16_6_inst : DLH_X1 port map( G => n268, D => n429_port, Q => 
                           REGISTERS_16_6_port);
   REGISTERS_reg_16_5_inst : DLH_X1 port map( G => n268, D => n433_port, Q => 
                           REGISTERS_16_5_port);
   REGISTERS_reg_16_4_inst : DLH_X1 port map( G => n268, D => n437_port, Q => 
                           REGISTERS_16_4_port);
   REGISTERS_reg_16_3_inst : DLH_X1 port map( G => n268, D => n441_port, Q => 
                           REGISTERS_16_3_port);
   REGISTERS_reg_16_2_inst : DLH_X1 port map( G => n268, D => n445, Q => 
                           REGISTERS_16_2_port);
   REGISTERS_reg_16_1_inst : DLH_X1 port map( G => n268, D => n449, Q => 
                           REGISTERS_16_1_port);
   REGISTERS_reg_16_0_inst : DLH_X1 port map( G => n268, D => n453, Q => 
                           REGISTERS_16_0_port);
   REGISTERS_reg_17_31_inst : DLH_X1 port map( G => n275, D => n329_port, Q => 
                           REGISTERS_17_31_port);
   REGISTERS_reg_17_30_inst : DLH_X1 port map( G => n275, D => n333_port, Q => 
                           REGISTERS_17_30_port);
   REGISTERS_reg_17_29_inst : DLH_X1 port map( G => n274, D => n337_port, Q => 
                           REGISTERS_17_29_port);
   REGISTERS_reg_17_28_inst : DLH_X1 port map( G => n274, D => n341_port, Q => 
                           REGISTERS_17_28_port);
   REGISTERS_reg_17_27_inst : DLH_X1 port map( G => n274, D => n345_port, Q => 
                           REGISTERS_17_27_port);
   REGISTERS_reg_17_26_inst : DLH_X1 port map( G => n274, D => n349_port, Q => 
                           REGISTERS_17_26_port);
   REGISTERS_reg_17_25_inst : DLH_X1 port map( G => n274, D => n353_port, Q => 
                           REGISTERS_17_25_port);
   REGISTERS_reg_17_24_inst : DLH_X1 port map( G => n274, D => n357_port, Q => 
                           REGISTERS_17_24_port);
   REGISTERS_reg_17_23_inst : DLH_X1 port map( G => n274, D => n361_port, Q => 
                           REGISTERS_17_23_port);
   REGISTERS_reg_17_22_inst : DLH_X1 port map( G => n274, D => n365_port, Q => 
                           REGISTERS_17_22_port);
   REGISTERS_reg_17_21_inst : DLH_X1 port map( G => n274, D => n369_port, Q => 
                           REGISTERS_17_21_port);
   REGISTERS_reg_17_20_inst : DLH_X1 port map( G => n274, D => n373_port, Q => 
                           REGISTERS_17_20_port);
   REGISTERS_reg_17_19_inst : DLH_X1 port map( G => n273, D => n377_port, Q => 
                           REGISTERS_17_19_port);
   REGISTERS_reg_17_18_inst : DLH_X1 port map( G => n273, D => n381_port, Q => 
                           REGISTERS_17_18_port);
   REGISTERS_reg_17_17_inst : DLH_X1 port map( G => n273, D => n385_port, Q => 
                           REGISTERS_17_17_port);
   REGISTERS_reg_17_16_inst : DLH_X1 port map( G => n273, D => n389_port, Q => 
                           REGISTERS_17_16_port);
   REGISTERS_reg_17_15_inst : DLH_X1 port map( G => n273, D => n393_port, Q => 
                           REGISTERS_17_15_port);
   REGISTERS_reg_17_14_inst : DLH_X1 port map( G => n273, D => n397_port, Q => 
                           REGISTERS_17_14_port);
   REGISTERS_reg_17_13_inst : DLH_X1 port map( G => n273, D => n401_port, Q => 
                           REGISTERS_17_13_port);
   REGISTERS_reg_17_12_inst : DLH_X1 port map( G => n273, D => n405_port, Q => 
                           REGISTERS_17_12_port);
   REGISTERS_reg_17_11_inst : DLH_X1 port map( G => n273, D => n409_port, Q => 
                           REGISTERS_17_11_port);
   REGISTERS_reg_17_10_inst : DLH_X1 port map( G => n273, D => n413_port, Q => 
                           REGISTERS_17_10_port);
   REGISTERS_reg_17_9_inst : DLH_X1 port map( G => n272, D => n417_port, Q => 
                           REGISTERS_17_9_port);
   REGISTERS_reg_17_8_inst : DLH_X1 port map( G => n272, D => n421_port, Q => 
                           REGISTERS_17_8_port);
   REGISTERS_reg_17_7_inst : DLH_X1 port map( G => n272, D => n425_port, Q => 
                           REGISTERS_17_7_port);
   REGISTERS_reg_17_6_inst : DLH_X1 port map( G => n272, D => n429_port, Q => 
                           REGISTERS_17_6_port);
   REGISTERS_reg_17_5_inst : DLH_X1 port map( G => n272, D => n433_port, Q => 
                           REGISTERS_17_5_port);
   REGISTERS_reg_17_4_inst : DLH_X1 port map( G => n272, D => n437_port, Q => 
                           REGISTERS_17_4_port);
   REGISTERS_reg_17_3_inst : DLH_X1 port map( G => n272, D => n441_port, Q => 
                           REGISTERS_17_3_port);
   REGISTERS_reg_17_2_inst : DLH_X1 port map( G => n272, D => n445, Q => 
                           REGISTERS_17_2_port);
   REGISTERS_reg_17_1_inst : DLH_X1 port map( G => n272, D => n449, Q => 
                           REGISTERS_17_1_port);
   REGISTERS_reg_17_0_inst : DLH_X1 port map( G => n272, D => n453, Q => 
                           REGISTERS_17_0_port);
   REGISTERS_reg_18_31_inst : DLH_X1 port map( G => n279, D => n329_port, Q => 
                           REGISTERS_18_31_port);
   REGISTERS_reg_18_30_inst : DLH_X1 port map( G => n279, D => n333_port, Q => 
                           REGISTERS_18_30_port);
   REGISTERS_reg_18_29_inst : DLH_X1 port map( G => n278, D => n337_port, Q => 
                           REGISTERS_18_29_port);
   REGISTERS_reg_18_28_inst : DLH_X1 port map( G => n278, D => n341_port, Q => 
                           REGISTERS_18_28_port);
   REGISTERS_reg_18_27_inst : DLH_X1 port map( G => n278, D => n345_port, Q => 
                           REGISTERS_18_27_port);
   REGISTERS_reg_18_26_inst : DLH_X1 port map( G => n278, D => n349_port, Q => 
                           REGISTERS_18_26_port);
   REGISTERS_reg_18_25_inst : DLH_X1 port map( G => n278, D => n353_port, Q => 
                           REGISTERS_18_25_port);
   REGISTERS_reg_18_24_inst : DLH_X1 port map( G => n278, D => n357_port, Q => 
                           REGISTERS_18_24_port);
   REGISTERS_reg_18_23_inst : DLH_X1 port map( G => n278, D => n361_port, Q => 
                           REGISTERS_18_23_port);
   REGISTERS_reg_18_22_inst : DLH_X1 port map( G => n278, D => n365_port, Q => 
                           REGISTERS_18_22_port);
   REGISTERS_reg_18_21_inst : DLH_X1 port map( G => n278, D => n369_port, Q => 
                           REGISTERS_18_21_port);
   REGISTERS_reg_18_20_inst : DLH_X1 port map( G => n278, D => n373_port, Q => 
                           REGISTERS_18_20_port);
   REGISTERS_reg_18_19_inst : DLH_X1 port map( G => n277, D => n377_port, Q => 
                           REGISTERS_18_19_port);
   REGISTERS_reg_18_18_inst : DLH_X1 port map( G => n277, D => n381_port, Q => 
                           REGISTERS_18_18_port);
   REGISTERS_reg_18_17_inst : DLH_X1 port map( G => n277, D => n385_port, Q => 
                           REGISTERS_18_17_port);
   REGISTERS_reg_18_16_inst : DLH_X1 port map( G => n277, D => n389_port, Q => 
                           REGISTERS_18_16_port);
   REGISTERS_reg_18_15_inst : DLH_X1 port map( G => n277, D => n393_port, Q => 
                           REGISTERS_18_15_port);
   REGISTERS_reg_18_14_inst : DLH_X1 port map( G => n277, D => n397_port, Q => 
                           REGISTERS_18_14_port);
   REGISTERS_reg_18_13_inst : DLH_X1 port map( G => n277, D => n401_port, Q => 
                           REGISTERS_18_13_port);
   REGISTERS_reg_18_12_inst : DLH_X1 port map( G => n277, D => n405_port, Q => 
                           REGISTERS_18_12_port);
   REGISTERS_reg_18_11_inst : DLH_X1 port map( G => n277, D => n409_port, Q => 
                           REGISTERS_18_11_port);
   REGISTERS_reg_18_10_inst : DLH_X1 port map( G => n277, D => n413_port, Q => 
                           REGISTERS_18_10_port);
   REGISTERS_reg_18_9_inst : DLH_X1 port map( G => n276, D => n417_port, Q => 
                           REGISTERS_18_9_port);
   REGISTERS_reg_18_8_inst : DLH_X1 port map( G => n276, D => n421_port, Q => 
                           REGISTERS_18_8_port);
   REGISTERS_reg_18_7_inst : DLH_X1 port map( G => n276, D => n425_port, Q => 
                           REGISTERS_18_7_port);
   REGISTERS_reg_18_6_inst : DLH_X1 port map( G => n276, D => n429_port, Q => 
                           REGISTERS_18_6_port);
   REGISTERS_reg_18_5_inst : DLH_X1 port map( G => n276, D => n433_port, Q => 
                           REGISTERS_18_5_port);
   REGISTERS_reg_18_4_inst : DLH_X1 port map( G => n276, D => n437_port, Q => 
                           REGISTERS_18_4_port);
   REGISTERS_reg_18_3_inst : DLH_X1 port map( G => n276, D => n441_port, Q => 
                           REGISTERS_18_3_port);
   REGISTERS_reg_18_2_inst : DLH_X1 port map( G => n276, D => n445, Q => 
                           REGISTERS_18_2_port);
   REGISTERS_reg_18_1_inst : DLH_X1 port map( G => n276, D => n449, Q => 
                           REGISTERS_18_1_port);
   REGISTERS_reg_18_0_inst : DLH_X1 port map( G => n276, D => n453, Q => 
                           REGISTERS_18_0_port);
   REGISTERS_reg_19_31_inst : DLH_X1 port map( G => n283, D => n329_port, Q => 
                           REGISTERS_19_31_port);
   REGISTERS_reg_19_30_inst : DLH_X1 port map( G => n283, D => n333_port, Q => 
                           REGISTERS_19_30_port);
   REGISTERS_reg_19_29_inst : DLH_X1 port map( G => n282, D => n337_port, Q => 
                           REGISTERS_19_29_port);
   REGISTERS_reg_19_28_inst : DLH_X1 port map( G => n282, D => n341_port, Q => 
                           REGISTERS_19_28_port);
   REGISTERS_reg_19_27_inst : DLH_X1 port map( G => n282, D => n345_port, Q => 
                           REGISTERS_19_27_port);
   REGISTERS_reg_19_26_inst : DLH_X1 port map( G => n282, D => n349_port, Q => 
                           REGISTERS_19_26_port);
   REGISTERS_reg_19_25_inst : DLH_X1 port map( G => n282, D => n353_port, Q => 
                           REGISTERS_19_25_port);
   REGISTERS_reg_19_24_inst : DLH_X1 port map( G => n282, D => n357_port, Q => 
                           REGISTERS_19_24_port);
   REGISTERS_reg_19_23_inst : DLH_X1 port map( G => n282, D => n361_port, Q => 
                           REGISTERS_19_23_port);
   REGISTERS_reg_19_22_inst : DLH_X1 port map( G => n282, D => n365_port, Q => 
                           REGISTERS_19_22_port);
   REGISTERS_reg_19_21_inst : DLH_X1 port map( G => n282, D => n369_port, Q => 
                           REGISTERS_19_21_port);
   REGISTERS_reg_19_20_inst : DLH_X1 port map( G => n282, D => n373_port, Q => 
                           REGISTERS_19_20_port);
   REGISTERS_reg_19_19_inst : DLH_X1 port map( G => n281, D => n377_port, Q => 
                           REGISTERS_19_19_port);
   REGISTERS_reg_19_18_inst : DLH_X1 port map( G => n281, D => n381_port, Q => 
                           REGISTERS_19_18_port);
   REGISTERS_reg_19_17_inst : DLH_X1 port map( G => n281, D => n385_port, Q => 
                           REGISTERS_19_17_port);
   REGISTERS_reg_19_16_inst : DLH_X1 port map( G => n281, D => n389_port, Q => 
                           REGISTERS_19_16_port);
   REGISTERS_reg_19_15_inst : DLH_X1 port map( G => n281, D => n393_port, Q => 
                           REGISTERS_19_15_port);
   REGISTERS_reg_19_14_inst : DLH_X1 port map( G => n281, D => n397_port, Q => 
                           REGISTERS_19_14_port);
   REGISTERS_reg_19_13_inst : DLH_X1 port map( G => n281, D => n401_port, Q => 
                           REGISTERS_19_13_port);
   REGISTERS_reg_19_12_inst : DLH_X1 port map( G => n281, D => n405_port, Q => 
                           REGISTERS_19_12_port);
   REGISTERS_reg_19_11_inst : DLH_X1 port map( G => n281, D => n409_port, Q => 
                           REGISTERS_19_11_port);
   REGISTERS_reg_19_10_inst : DLH_X1 port map( G => n281, D => n413_port, Q => 
                           REGISTERS_19_10_port);
   REGISTERS_reg_19_9_inst : DLH_X1 port map( G => n280, D => n417_port, Q => 
                           REGISTERS_19_9_port);
   REGISTERS_reg_19_8_inst : DLH_X1 port map( G => n280, D => n421_port, Q => 
                           REGISTERS_19_8_port);
   REGISTERS_reg_19_7_inst : DLH_X1 port map( G => n280, D => n425_port, Q => 
                           REGISTERS_19_7_port);
   REGISTERS_reg_19_6_inst : DLH_X1 port map( G => n280, D => n429_port, Q => 
                           REGISTERS_19_6_port);
   REGISTERS_reg_19_5_inst : DLH_X1 port map( G => n280, D => n433_port, Q => 
                           REGISTERS_19_5_port);
   REGISTERS_reg_19_4_inst : DLH_X1 port map( G => n280, D => n437_port, Q => 
                           REGISTERS_19_4_port);
   REGISTERS_reg_19_3_inst : DLH_X1 port map( G => n280, D => n441_port, Q => 
                           REGISTERS_19_3_port);
   REGISTERS_reg_19_2_inst : DLH_X1 port map( G => n280, D => n445, Q => 
                           REGISTERS_19_2_port);
   REGISTERS_reg_19_1_inst : DLH_X1 port map( G => n280, D => n449, Q => 
                           REGISTERS_19_1_port);
   REGISTERS_reg_19_0_inst : DLH_X1 port map( G => n280, D => n453, Q => 
                           REGISTERS_19_0_port);
   REGISTERS_reg_20_31_inst : DLH_X1 port map( G => n287, D => n330_port, Q => 
                           REGISTERS_20_31_port);
   REGISTERS_reg_20_30_inst : DLH_X1 port map( G => n287, D => n334_port, Q => 
                           REGISTERS_20_30_port);
   REGISTERS_reg_20_29_inst : DLH_X1 port map( G => n286, D => n338_port, Q => 
                           REGISTERS_20_29_port);
   REGISTERS_reg_20_28_inst : DLH_X1 port map( G => n286, D => n342_port, Q => 
                           REGISTERS_20_28_port);
   REGISTERS_reg_20_27_inst : DLH_X1 port map( G => n286, D => n346_port, Q => 
                           REGISTERS_20_27_port);
   REGISTERS_reg_20_26_inst : DLH_X1 port map( G => n286, D => n350_port, Q => 
                           REGISTERS_20_26_port);
   REGISTERS_reg_20_25_inst : DLH_X1 port map( G => n286, D => n354_port, Q => 
                           REGISTERS_20_25_port);
   REGISTERS_reg_20_24_inst : DLH_X1 port map( G => n286, D => n358_port, Q => 
                           REGISTERS_20_24_port);
   REGISTERS_reg_20_23_inst : DLH_X1 port map( G => n286, D => n362_port, Q => 
                           REGISTERS_20_23_port);
   REGISTERS_reg_20_22_inst : DLH_X1 port map( G => n286, D => n366_port, Q => 
                           REGISTERS_20_22_port);
   REGISTERS_reg_20_21_inst : DLH_X1 port map( G => n286, D => n370_port, Q => 
                           REGISTERS_20_21_port);
   REGISTERS_reg_20_20_inst : DLH_X1 port map( G => n286, D => n374_port, Q => 
                           REGISTERS_20_20_port);
   REGISTERS_reg_20_19_inst : DLH_X1 port map( G => n285, D => n378_port, Q => 
                           REGISTERS_20_19_port);
   REGISTERS_reg_20_18_inst : DLH_X1 port map( G => n285, D => n382_port, Q => 
                           REGISTERS_20_18_port);
   REGISTERS_reg_20_17_inst : DLH_X1 port map( G => n285, D => n386_port, Q => 
                           REGISTERS_20_17_port);
   REGISTERS_reg_20_16_inst : DLH_X1 port map( G => n285, D => n390_port, Q => 
                           REGISTERS_20_16_port);
   REGISTERS_reg_20_15_inst : DLH_X1 port map( G => n285, D => n394_port, Q => 
                           REGISTERS_20_15_port);
   REGISTERS_reg_20_14_inst : DLH_X1 port map( G => n285, D => n398_port, Q => 
                           REGISTERS_20_14_port);
   REGISTERS_reg_20_13_inst : DLH_X1 port map( G => n285, D => n402_port, Q => 
                           REGISTERS_20_13_port);
   REGISTERS_reg_20_12_inst : DLH_X1 port map( G => n285, D => n406_port, Q => 
                           REGISTERS_20_12_port);
   REGISTERS_reg_20_11_inst : DLH_X1 port map( G => n285, D => n410_port, Q => 
                           REGISTERS_20_11_port);
   REGISTERS_reg_20_10_inst : DLH_X1 port map( G => n285, D => n414_port, Q => 
                           REGISTERS_20_10_port);
   REGISTERS_reg_20_9_inst : DLH_X1 port map( G => n284, D => n418_port, Q => 
                           REGISTERS_20_9_port);
   REGISTERS_reg_20_8_inst : DLH_X1 port map( G => n284, D => n422_port, Q => 
                           REGISTERS_20_8_port);
   REGISTERS_reg_20_7_inst : DLH_X1 port map( G => n284, D => n426_port, Q => 
                           REGISTERS_20_7_port);
   REGISTERS_reg_20_6_inst : DLH_X1 port map( G => n284, D => n430_port, Q => 
                           REGISTERS_20_6_port);
   REGISTERS_reg_20_5_inst : DLH_X1 port map( G => n284, D => n434_port, Q => 
                           REGISTERS_20_5_port);
   REGISTERS_reg_20_4_inst : DLH_X1 port map( G => n284, D => n438_port, Q => 
                           REGISTERS_20_4_port);
   REGISTERS_reg_20_3_inst : DLH_X1 port map( G => n284, D => n442, Q => 
                           REGISTERS_20_3_port);
   REGISTERS_reg_20_2_inst : DLH_X1 port map( G => n284, D => n446, Q => 
                           REGISTERS_20_2_port);
   REGISTERS_reg_20_1_inst : DLH_X1 port map( G => n284, D => n450, Q => 
                           REGISTERS_20_1_port);
   REGISTERS_reg_20_0_inst : DLH_X1 port map( G => n284, D => n454, Q => 
                           REGISTERS_20_0_port);
   REGISTERS_reg_21_31_inst : DLH_X1 port map( G => n291, D => n330_port, Q => 
                           REGISTERS_21_31_port);
   REGISTERS_reg_21_30_inst : DLH_X1 port map( G => n291, D => n334_port, Q => 
                           REGISTERS_21_30_port);
   REGISTERS_reg_21_29_inst : DLH_X1 port map( G => n290, D => n338_port, Q => 
                           REGISTERS_21_29_port);
   REGISTERS_reg_21_28_inst : DLH_X1 port map( G => n290, D => n342_port, Q => 
                           REGISTERS_21_28_port);
   REGISTERS_reg_21_27_inst : DLH_X1 port map( G => n290, D => n346_port, Q => 
                           REGISTERS_21_27_port);
   REGISTERS_reg_21_26_inst : DLH_X1 port map( G => n290, D => n350_port, Q => 
                           REGISTERS_21_26_port);
   REGISTERS_reg_21_25_inst : DLH_X1 port map( G => n290, D => n354_port, Q => 
                           REGISTERS_21_25_port);
   REGISTERS_reg_21_24_inst : DLH_X1 port map( G => n290, D => n358_port, Q => 
                           REGISTERS_21_24_port);
   REGISTERS_reg_21_23_inst : DLH_X1 port map( G => n290, D => n362_port, Q => 
                           REGISTERS_21_23_port);
   REGISTERS_reg_21_22_inst : DLH_X1 port map( G => n290, D => n366_port, Q => 
                           REGISTERS_21_22_port);
   REGISTERS_reg_21_21_inst : DLH_X1 port map( G => n290, D => n370_port, Q => 
                           REGISTERS_21_21_port);
   REGISTERS_reg_21_20_inst : DLH_X1 port map( G => n290, D => n374_port, Q => 
                           REGISTERS_21_20_port);
   REGISTERS_reg_21_19_inst : DLH_X1 port map( G => n289, D => n378_port, Q => 
                           REGISTERS_21_19_port);
   REGISTERS_reg_21_18_inst : DLH_X1 port map( G => n289, D => n382_port, Q => 
                           REGISTERS_21_18_port);
   REGISTERS_reg_21_17_inst : DLH_X1 port map( G => n289, D => n386_port, Q => 
                           REGISTERS_21_17_port);
   REGISTERS_reg_21_16_inst : DLH_X1 port map( G => n289, D => n390_port, Q => 
                           REGISTERS_21_16_port);
   REGISTERS_reg_21_15_inst : DLH_X1 port map( G => n289, D => n394_port, Q => 
                           REGISTERS_21_15_port);
   REGISTERS_reg_21_14_inst : DLH_X1 port map( G => n289, D => n398_port, Q => 
                           REGISTERS_21_14_port);
   REGISTERS_reg_21_13_inst : DLH_X1 port map( G => n289, D => n402_port, Q => 
                           REGISTERS_21_13_port);
   REGISTERS_reg_21_12_inst : DLH_X1 port map( G => n289, D => n406_port, Q => 
                           REGISTERS_21_12_port);
   REGISTERS_reg_21_11_inst : DLH_X1 port map( G => n289, D => n410_port, Q => 
                           REGISTERS_21_11_port);
   REGISTERS_reg_21_10_inst : DLH_X1 port map( G => n289, D => n414_port, Q => 
                           REGISTERS_21_10_port);
   REGISTERS_reg_21_9_inst : DLH_X1 port map( G => n288, D => n418_port, Q => 
                           REGISTERS_21_9_port);
   REGISTERS_reg_21_8_inst : DLH_X1 port map( G => n288, D => n422_port, Q => 
                           REGISTERS_21_8_port);
   REGISTERS_reg_21_7_inst : DLH_X1 port map( G => n288, D => n426_port, Q => 
                           REGISTERS_21_7_port);
   REGISTERS_reg_21_6_inst : DLH_X1 port map( G => n288, D => n430_port, Q => 
                           REGISTERS_21_6_port);
   REGISTERS_reg_21_5_inst : DLH_X1 port map( G => n288, D => n434_port, Q => 
                           REGISTERS_21_5_port);
   REGISTERS_reg_21_4_inst : DLH_X1 port map( G => n288, D => n438_port, Q => 
                           REGISTERS_21_4_port);
   REGISTERS_reg_21_3_inst : DLH_X1 port map( G => n288, D => n442, Q => 
                           REGISTERS_21_3_port);
   REGISTERS_reg_21_2_inst : DLH_X1 port map( G => n288, D => n446, Q => 
                           REGISTERS_21_2_port);
   REGISTERS_reg_21_1_inst : DLH_X1 port map( G => n288, D => n450, Q => 
                           REGISTERS_21_1_port);
   REGISTERS_reg_21_0_inst : DLH_X1 port map( G => n288, D => n454, Q => 
                           REGISTERS_21_0_port);
   REGISTERS_reg_22_31_inst : DLH_X1 port map( G => n295, D => n330_port, Q => 
                           REGISTERS_22_31_port);
   REGISTERS_reg_22_30_inst : DLH_X1 port map( G => n295, D => n334_port, Q => 
                           REGISTERS_22_30_port);
   REGISTERS_reg_22_29_inst : DLH_X1 port map( G => n294, D => n338_port, Q => 
                           REGISTERS_22_29_port);
   REGISTERS_reg_22_28_inst : DLH_X1 port map( G => n294, D => n342_port, Q => 
                           REGISTERS_22_28_port);
   REGISTERS_reg_22_27_inst : DLH_X1 port map( G => n294, D => n346_port, Q => 
                           REGISTERS_22_27_port);
   REGISTERS_reg_22_26_inst : DLH_X1 port map( G => n294, D => n350_port, Q => 
                           REGISTERS_22_26_port);
   REGISTERS_reg_22_25_inst : DLH_X1 port map( G => n294, D => n354_port, Q => 
                           REGISTERS_22_25_port);
   REGISTERS_reg_22_24_inst : DLH_X1 port map( G => n294, D => n358_port, Q => 
                           REGISTERS_22_24_port);
   REGISTERS_reg_22_23_inst : DLH_X1 port map( G => n294, D => n362_port, Q => 
                           REGISTERS_22_23_port);
   REGISTERS_reg_22_22_inst : DLH_X1 port map( G => n294, D => n366_port, Q => 
                           REGISTERS_22_22_port);
   REGISTERS_reg_22_21_inst : DLH_X1 port map( G => n294, D => n370_port, Q => 
                           REGISTERS_22_21_port);
   REGISTERS_reg_22_20_inst : DLH_X1 port map( G => n294, D => n374_port, Q => 
                           REGISTERS_22_20_port);
   REGISTERS_reg_22_19_inst : DLH_X1 port map( G => n293, D => n378_port, Q => 
                           REGISTERS_22_19_port);
   REGISTERS_reg_22_18_inst : DLH_X1 port map( G => n293, D => n382_port, Q => 
                           REGISTERS_22_18_port);
   REGISTERS_reg_22_17_inst : DLH_X1 port map( G => n293, D => n386_port, Q => 
                           REGISTERS_22_17_port);
   REGISTERS_reg_22_16_inst : DLH_X1 port map( G => n293, D => n390_port, Q => 
                           REGISTERS_22_16_port);
   REGISTERS_reg_22_15_inst : DLH_X1 port map( G => n293, D => n394_port, Q => 
                           REGISTERS_22_15_port);
   REGISTERS_reg_22_14_inst : DLH_X1 port map( G => n293, D => n398_port, Q => 
                           REGISTERS_22_14_port);
   REGISTERS_reg_22_13_inst : DLH_X1 port map( G => n293, D => n402_port, Q => 
                           REGISTERS_22_13_port);
   REGISTERS_reg_22_12_inst : DLH_X1 port map( G => n293, D => n406_port, Q => 
                           REGISTERS_22_12_port);
   REGISTERS_reg_22_11_inst : DLH_X1 port map( G => n293, D => n410_port, Q => 
                           REGISTERS_22_11_port);
   REGISTERS_reg_22_10_inst : DLH_X1 port map( G => n293, D => n414_port, Q => 
                           REGISTERS_22_10_port);
   REGISTERS_reg_22_9_inst : DLH_X1 port map( G => n292, D => n418_port, Q => 
                           REGISTERS_22_9_port);
   REGISTERS_reg_22_8_inst : DLH_X1 port map( G => n292, D => n422_port, Q => 
                           REGISTERS_22_8_port);
   REGISTERS_reg_22_7_inst : DLH_X1 port map( G => n292, D => n426_port, Q => 
                           REGISTERS_22_7_port);
   REGISTERS_reg_22_6_inst : DLH_X1 port map( G => n292, D => n430_port, Q => 
                           REGISTERS_22_6_port);
   REGISTERS_reg_22_5_inst : DLH_X1 port map( G => n292, D => n434_port, Q => 
                           REGISTERS_22_5_port);
   REGISTERS_reg_22_4_inst : DLH_X1 port map( G => n292, D => n438_port, Q => 
                           REGISTERS_22_4_port);
   REGISTERS_reg_22_3_inst : DLH_X1 port map( G => n292, D => n442, Q => 
                           REGISTERS_22_3_port);
   REGISTERS_reg_22_2_inst : DLH_X1 port map( G => n292, D => n446, Q => 
                           REGISTERS_22_2_port);
   REGISTERS_reg_22_1_inst : DLH_X1 port map( G => n292, D => n450, Q => 
                           REGISTERS_22_1_port);
   REGISTERS_reg_22_0_inst : DLH_X1 port map( G => n292, D => n454, Q => 
                           REGISTERS_22_0_port);
   REGISTERS_reg_23_31_inst : DLH_X1 port map( G => n299, D => n330_port, Q => 
                           REGISTERS_23_31_port);
   REGISTERS_reg_23_30_inst : DLH_X1 port map( G => n299, D => n334_port, Q => 
                           REGISTERS_23_30_port);
   REGISTERS_reg_23_29_inst : DLH_X1 port map( G => n298, D => n338_port, Q => 
                           REGISTERS_23_29_port);
   REGISTERS_reg_23_28_inst : DLH_X1 port map( G => n298, D => n342_port, Q => 
                           REGISTERS_23_28_port);
   REGISTERS_reg_23_27_inst : DLH_X1 port map( G => n298, D => n346_port, Q => 
                           REGISTERS_23_27_port);
   REGISTERS_reg_23_26_inst : DLH_X1 port map( G => n298, D => n350_port, Q => 
                           REGISTERS_23_26_port);
   REGISTERS_reg_23_25_inst : DLH_X1 port map( G => n298, D => n354_port, Q => 
                           REGISTERS_23_25_port);
   REGISTERS_reg_23_24_inst : DLH_X1 port map( G => n298, D => n358_port, Q => 
                           REGISTERS_23_24_port);
   REGISTERS_reg_23_23_inst : DLH_X1 port map( G => n298, D => n362_port, Q => 
                           REGISTERS_23_23_port);
   REGISTERS_reg_23_22_inst : DLH_X1 port map( G => n298, D => n366_port, Q => 
                           REGISTERS_23_22_port);
   REGISTERS_reg_23_21_inst : DLH_X1 port map( G => n298, D => n370_port, Q => 
                           REGISTERS_23_21_port);
   REGISTERS_reg_23_20_inst : DLH_X1 port map( G => n298, D => n374_port, Q => 
                           REGISTERS_23_20_port);
   REGISTERS_reg_23_19_inst : DLH_X1 port map( G => n297, D => n378_port, Q => 
                           REGISTERS_23_19_port);
   REGISTERS_reg_23_18_inst : DLH_X1 port map( G => n297, D => n382_port, Q => 
                           REGISTERS_23_18_port);
   REGISTERS_reg_23_17_inst : DLH_X1 port map( G => n297, D => n386_port, Q => 
                           REGISTERS_23_17_port);
   REGISTERS_reg_23_16_inst : DLH_X1 port map( G => n297, D => n390_port, Q => 
                           REGISTERS_23_16_port);
   REGISTERS_reg_23_15_inst : DLH_X1 port map( G => n297, D => n394_port, Q => 
                           REGISTERS_23_15_port);
   REGISTERS_reg_23_14_inst : DLH_X1 port map( G => n297, D => n398_port, Q => 
                           REGISTERS_23_14_port);
   REGISTERS_reg_23_13_inst : DLH_X1 port map( G => n297, D => n402_port, Q => 
                           REGISTERS_23_13_port);
   REGISTERS_reg_23_12_inst : DLH_X1 port map( G => n297, D => n406_port, Q => 
                           REGISTERS_23_12_port);
   REGISTERS_reg_23_11_inst : DLH_X1 port map( G => n297, D => n410_port, Q => 
                           REGISTERS_23_11_port);
   REGISTERS_reg_23_10_inst : DLH_X1 port map( G => n297, D => n414_port, Q => 
                           REGISTERS_23_10_port);
   REGISTERS_reg_23_9_inst : DLH_X1 port map( G => n296, D => n418_port, Q => 
                           REGISTERS_23_9_port);
   REGISTERS_reg_23_8_inst : DLH_X1 port map( G => n296, D => n422_port, Q => 
                           REGISTERS_23_8_port);
   REGISTERS_reg_23_7_inst : DLH_X1 port map( G => n296, D => n426_port, Q => 
                           REGISTERS_23_7_port);
   REGISTERS_reg_23_6_inst : DLH_X1 port map( G => n296, D => n430_port, Q => 
                           REGISTERS_23_6_port);
   REGISTERS_reg_23_5_inst : DLH_X1 port map( G => n296, D => n434_port, Q => 
                           REGISTERS_23_5_port);
   REGISTERS_reg_23_4_inst : DLH_X1 port map( G => n296, D => n438_port, Q => 
                           REGISTERS_23_4_port);
   REGISTERS_reg_23_3_inst : DLH_X1 port map( G => n296, D => n442, Q => 
                           REGISTERS_23_3_port);
   REGISTERS_reg_23_2_inst : DLH_X1 port map( G => n296, D => n446, Q => 
                           REGISTERS_23_2_port);
   REGISTERS_reg_23_1_inst : DLH_X1 port map( G => n296, D => n450, Q => 
                           REGISTERS_23_1_port);
   REGISTERS_reg_23_0_inst : DLH_X1 port map( G => n296, D => n454, Q => 
                           REGISTERS_23_0_port);
   REGISTERS_reg_24_31_inst : DLH_X1 port map( G => n303, D => n330_port, Q => 
                           REGISTERS_24_31_port);
   REGISTERS_reg_24_30_inst : DLH_X1 port map( G => n303, D => n334_port, Q => 
                           REGISTERS_24_30_port);
   REGISTERS_reg_24_29_inst : DLH_X1 port map( G => n302, D => n338_port, Q => 
                           REGISTERS_24_29_port);
   REGISTERS_reg_24_28_inst : DLH_X1 port map( G => n302, D => n342_port, Q => 
                           REGISTERS_24_28_port);
   REGISTERS_reg_24_27_inst : DLH_X1 port map( G => n302, D => n346_port, Q => 
                           REGISTERS_24_27_port);
   REGISTERS_reg_24_26_inst : DLH_X1 port map( G => n302, D => n350_port, Q => 
                           REGISTERS_24_26_port);
   REGISTERS_reg_24_25_inst : DLH_X1 port map( G => n302, D => n354_port, Q => 
                           REGISTERS_24_25_port);
   REGISTERS_reg_24_24_inst : DLH_X1 port map( G => n302, D => n358_port, Q => 
                           REGISTERS_24_24_port);
   REGISTERS_reg_24_23_inst : DLH_X1 port map( G => n302, D => n362_port, Q => 
                           REGISTERS_24_23_port);
   REGISTERS_reg_24_22_inst : DLH_X1 port map( G => n302, D => n366_port, Q => 
                           REGISTERS_24_22_port);
   REGISTERS_reg_24_21_inst : DLH_X1 port map( G => n302, D => n370_port, Q => 
                           REGISTERS_24_21_port);
   REGISTERS_reg_24_20_inst : DLH_X1 port map( G => n302, D => n374_port, Q => 
                           REGISTERS_24_20_port);
   REGISTERS_reg_24_19_inst : DLH_X1 port map( G => n301, D => n378_port, Q => 
                           REGISTERS_24_19_port);
   REGISTERS_reg_24_18_inst : DLH_X1 port map( G => n301, D => n382_port, Q => 
                           REGISTERS_24_18_port);
   REGISTERS_reg_24_17_inst : DLH_X1 port map( G => n301, D => n386_port, Q => 
                           REGISTERS_24_17_port);
   REGISTERS_reg_24_16_inst : DLH_X1 port map( G => n301, D => n390_port, Q => 
                           REGISTERS_24_16_port);
   REGISTERS_reg_24_15_inst : DLH_X1 port map( G => n301, D => n394_port, Q => 
                           REGISTERS_24_15_port);
   REGISTERS_reg_24_14_inst : DLH_X1 port map( G => n301, D => n398_port, Q => 
                           REGISTERS_24_14_port);
   REGISTERS_reg_24_13_inst : DLH_X1 port map( G => n301, D => n402_port, Q => 
                           REGISTERS_24_13_port);
   REGISTERS_reg_24_12_inst : DLH_X1 port map( G => n301, D => n406_port, Q => 
                           REGISTERS_24_12_port);
   REGISTERS_reg_24_11_inst : DLH_X1 port map( G => n301, D => n410_port, Q => 
                           REGISTERS_24_11_port);
   REGISTERS_reg_24_10_inst : DLH_X1 port map( G => n301, D => n414_port, Q => 
                           REGISTERS_24_10_port);
   REGISTERS_reg_24_9_inst : DLH_X1 port map( G => n300, D => n418_port, Q => 
                           REGISTERS_24_9_port);
   REGISTERS_reg_24_8_inst : DLH_X1 port map( G => n300, D => n422_port, Q => 
                           REGISTERS_24_8_port);
   REGISTERS_reg_24_7_inst : DLH_X1 port map( G => n300, D => n426_port, Q => 
                           REGISTERS_24_7_port);
   REGISTERS_reg_24_6_inst : DLH_X1 port map( G => n300, D => n430_port, Q => 
                           REGISTERS_24_6_port);
   REGISTERS_reg_24_5_inst : DLH_X1 port map( G => n300, D => n434_port, Q => 
                           REGISTERS_24_5_port);
   REGISTERS_reg_24_4_inst : DLH_X1 port map( G => n300, D => n438_port, Q => 
                           REGISTERS_24_4_port);
   REGISTERS_reg_24_3_inst : DLH_X1 port map( G => n300, D => n442, Q => 
                           REGISTERS_24_3_port);
   REGISTERS_reg_24_2_inst : DLH_X1 port map( G => n300, D => n446, Q => 
                           REGISTERS_24_2_port);
   REGISTERS_reg_24_1_inst : DLH_X1 port map( G => n300, D => n450, Q => 
                           REGISTERS_24_1_port);
   REGISTERS_reg_24_0_inst : DLH_X1 port map( G => n300, D => n454, Q => 
                           REGISTERS_24_0_port);
   REGISTERS_reg_25_31_inst : DLH_X1 port map( G => n307, D => n330_port, Q => 
                           REGISTERS_25_31_port);
   REGISTERS_reg_25_30_inst : DLH_X1 port map( G => n307, D => n334_port, Q => 
                           REGISTERS_25_30_port);
   REGISTERS_reg_25_29_inst : DLH_X1 port map( G => n306, D => n338_port, Q => 
                           REGISTERS_25_29_port);
   REGISTERS_reg_25_28_inst : DLH_X1 port map( G => n306, D => n342_port, Q => 
                           REGISTERS_25_28_port);
   REGISTERS_reg_25_27_inst : DLH_X1 port map( G => n306, D => n346_port, Q => 
                           REGISTERS_25_27_port);
   REGISTERS_reg_25_26_inst : DLH_X1 port map( G => n306, D => n350_port, Q => 
                           REGISTERS_25_26_port);
   REGISTERS_reg_25_25_inst : DLH_X1 port map( G => n306, D => n354_port, Q => 
                           REGISTERS_25_25_port);
   REGISTERS_reg_25_24_inst : DLH_X1 port map( G => n306, D => n358_port, Q => 
                           REGISTERS_25_24_port);
   REGISTERS_reg_25_23_inst : DLH_X1 port map( G => n306, D => n362_port, Q => 
                           REGISTERS_25_23_port);
   REGISTERS_reg_25_22_inst : DLH_X1 port map( G => n306, D => n366_port, Q => 
                           REGISTERS_25_22_port);
   REGISTERS_reg_25_21_inst : DLH_X1 port map( G => n306, D => n370_port, Q => 
                           REGISTERS_25_21_port);
   REGISTERS_reg_25_20_inst : DLH_X1 port map( G => n306, D => n374_port, Q => 
                           REGISTERS_25_20_port);
   REGISTERS_reg_25_19_inst : DLH_X1 port map( G => n305, D => n378_port, Q => 
                           REGISTERS_25_19_port);
   REGISTERS_reg_25_18_inst : DLH_X1 port map( G => n305, D => n382_port, Q => 
                           REGISTERS_25_18_port);
   REGISTERS_reg_25_17_inst : DLH_X1 port map( G => n305, D => n386_port, Q => 
                           REGISTERS_25_17_port);
   REGISTERS_reg_25_16_inst : DLH_X1 port map( G => n305, D => n390_port, Q => 
                           REGISTERS_25_16_port);
   REGISTERS_reg_25_15_inst : DLH_X1 port map( G => n305, D => n394_port, Q => 
                           REGISTERS_25_15_port);
   REGISTERS_reg_25_14_inst : DLH_X1 port map( G => n305, D => n398_port, Q => 
                           REGISTERS_25_14_port);
   REGISTERS_reg_25_13_inst : DLH_X1 port map( G => n305, D => n402_port, Q => 
                           REGISTERS_25_13_port);
   REGISTERS_reg_25_12_inst : DLH_X1 port map( G => n305, D => n406_port, Q => 
                           REGISTERS_25_12_port);
   REGISTERS_reg_25_11_inst : DLH_X1 port map( G => n305, D => n410_port, Q => 
                           REGISTERS_25_11_port);
   REGISTERS_reg_25_10_inst : DLH_X1 port map( G => n305, D => n414_port, Q => 
                           REGISTERS_25_10_port);
   REGISTERS_reg_25_9_inst : DLH_X1 port map( G => n304, D => n418_port, Q => 
                           REGISTERS_25_9_port);
   REGISTERS_reg_25_8_inst : DLH_X1 port map( G => n304, D => n422_port, Q => 
                           REGISTERS_25_8_port);
   REGISTERS_reg_25_7_inst : DLH_X1 port map( G => n304, D => n426_port, Q => 
                           REGISTERS_25_7_port);
   REGISTERS_reg_25_6_inst : DLH_X1 port map( G => n304, D => n430_port, Q => 
                           REGISTERS_25_6_port);
   REGISTERS_reg_25_5_inst : DLH_X1 port map( G => n304, D => n434_port, Q => 
                           REGISTERS_25_5_port);
   REGISTERS_reg_25_4_inst : DLH_X1 port map( G => n304, D => n438_port, Q => 
                           REGISTERS_25_4_port);
   REGISTERS_reg_25_3_inst : DLH_X1 port map( G => n304, D => n442, Q => 
                           REGISTERS_25_3_port);
   REGISTERS_reg_25_2_inst : DLH_X1 port map( G => n304, D => n446, Q => 
                           REGISTERS_25_2_port);
   REGISTERS_reg_25_1_inst : DLH_X1 port map( G => n304, D => n450, Q => 
                           REGISTERS_25_1_port);
   REGISTERS_reg_25_0_inst : DLH_X1 port map( G => n304, D => n454, Q => 
                           REGISTERS_25_0_port);
   REGISTERS_reg_26_31_inst : DLH_X1 port map( G => n311, D => n330_port, Q => 
                           REGISTERS_26_31_port);
   REGISTERS_reg_26_30_inst : DLH_X1 port map( G => n311, D => n334_port, Q => 
                           REGISTERS_26_30_port);
   REGISTERS_reg_26_29_inst : DLH_X1 port map( G => n310, D => n338_port, Q => 
                           REGISTERS_26_29_port);
   REGISTERS_reg_26_28_inst : DLH_X1 port map( G => n310, D => n342_port, Q => 
                           REGISTERS_26_28_port);
   REGISTERS_reg_26_27_inst : DLH_X1 port map( G => n310, D => n346_port, Q => 
                           REGISTERS_26_27_port);
   REGISTERS_reg_26_26_inst : DLH_X1 port map( G => n310, D => n350_port, Q => 
                           REGISTERS_26_26_port);
   REGISTERS_reg_26_25_inst : DLH_X1 port map( G => n310, D => n354_port, Q => 
                           REGISTERS_26_25_port);
   REGISTERS_reg_26_24_inst : DLH_X1 port map( G => n310, D => n358_port, Q => 
                           REGISTERS_26_24_port);
   REGISTERS_reg_26_23_inst : DLH_X1 port map( G => n310, D => n362_port, Q => 
                           REGISTERS_26_23_port);
   REGISTERS_reg_26_22_inst : DLH_X1 port map( G => n310, D => n366_port, Q => 
                           REGISTERS_26_22_port);
   REGISTERS_reg_26_21_inst : DLH_X1 port map( G => n310, D => n370_port, Q => 
                           REGISTERS_26_21_port);
   REGISTERS_reg_26_20_inst : DLH_X1 port map( G => n310, D => n374_port, Q => 
                           REGISTERS_26_20_port);
   REGISTERS_reg_26_19_inst : DLH_X1 port map( G => n309, D => n378_port, Q => 
                           REGISTERS_26_19_port);
   REGISTERS_reg_26_18_inst : DLH_X1 port map( G => n309, D => n382_port, Q => 
                           REGISTERS_26_18_port);
   REGISTERS_reg_26_17_inst : DLH_X1 port map( G => n309, D => n386_port, Q => 
                           REGISTERS_26_17_port);
   REGISTERS_reg_26_16_inst : DLH_X1 port map( G => n309, D => n390_port, Q => 
                           REGISTERS_26_16_port);
   REGISTERS_reg_26_15_inst : DLH_X1 port map( G => n309, D => n394_port, Q => 
                           REGISTERS_26_15_port);
   REGISTERS_reg_26_14_inst : DLH_X1 port map( G => n309, D => n398_port, Q => 
                           REGISTERS_26_14_port);
   REGISTERS_reg_26_13_inst : DLH_X1 port map( G => n309, D => n402_port, Q => 
                           REGISTERS_26_13_port);
   REGISTERS_reg_26_12_inst : DLH_X1 port map( G => n309, D => n406_port, Q => 
                           REGISTERS_26_12_port);
   REGISTERS_reg_26_11_inst : DLH_X1 port map( G => n309, D => n410_port, Q => 
                           REGISTERS_26_11_port);
   REGISTERS_reg_26_10_inst : DLH_X1 port map( G => n309, D => n414_port, Q => 
                           REGISTERS_26_10_port);
   REGISTERS_reg_26_9_inst : DLH_X1 port map( G => n308, D => n418_port, Q => 
                           REGISTERS_26_9_port);
   REGISTERS_reg_26_8_inst : DLH_X1 port map( G => n308, D => n422_port, Q => 
                           REGISTERS_26_8_port);
   REGISTERS_reg_26_7_inst : DLH_X1 port map( G => n308, D => n426_port, Q => 
                           REGISTERS_26_7_port);
   REGISTERS_reg_26_6_inst : DLH_X1 port map( G => n308, D => n430_port, Q => 
                           REGISTERS_26_6_port);
   REGISTERS_reg_26_5_inst : DLH_X1 port map( G => n308, D => n434_port, Q => 
                           REGISTERS_26_5_port);
   REGISTERS_reg_26_4_inst : DLH_X1 port map( G => n308, D => n438_port, Q => 
                           REGISTERS_26_4_port);
   REGISTERS_reg_26_3_inst : DLH_X1 port map( G => n308, D => n442, Q => 
                           REGISTERS_26_3_port);
   REGISTERS_reg_26_2_inst : DLH_X1 port map( G => n308, D => n446, Q => 
                           REGISTERS_26_2_port);
   REGISTERS_reg_26_1_inst : DLH_X1 port map( G => n308, D => n450, Q => 
                           REGISTERS_26_1_port);
   REGISTERS_reg_26_0_inst : DLH_X1 port map( G => n308, D => n454, Q => 
                           REGISTERS_26_0_port);
   REGISTERS_reg_27_31_inst : DLH_X1 port map( G => n315_port, D => n330_port, 
                           Q => REGISTERS_27_31_port);
   REGISTERS_reg_27_30_inst : DLH_X1 port map( G => n315_port, D => n334_port, 
                           Q => REGISTERS_27_30_port);
   REGISTERS_reg_27_29_inst : DLH_X1 port map( G => n314_port, D => n338_port, 
                           Q => REGISTERS_27_29_port);
   REGISTERS_reg_27_28_inst : DLH_X1 port map( G => n314_port, D => n342_port, 
                           Q => REGISTERS_27_28_port);
   REGISTERS_reg_27_27_inst : DLH_X1 port map( G => n314_port, D => n346_port, 
                           Q => REGISTERS_27_27_port);
   REGISTERS_reg_27_26_inst : DLH_X1 port map( G => n314_port, D => n350_port, 
                           Q => REGISTERS_27_26_port);
   REGISTERS_reg_27_25_inst : DLH_X1 port map( G => n314_port, D => n354_port, 
                           Q => REGISTERS_27_25_port);
   REGISTERS_reg_27_24_inst : DLH_X1 port map( G => n314_port, D => n358_port, 
                           Q => REGISTERS_27_24_port);
   REGISTERS_reg_27_23_inst : DLH_X1 port map( G => n314_port, D => n362_port, 
                           Q => REGISTERS_27_23_port);
   REGISTERS_reg_27_22_inst : DLH_X1 port map( G => n314_port, D => n366_port, 
                           Q => REGISTERS_27_22_port);
   REGISTERS_reg_27_21_inst : DLH_X1 port map( G => n314_port, D => n370_port, 
                           Q => REGISTERS_27_21_port);
   REGISTERS_reg_27_20_inst : DLH_X1 port map( G => n314_port, D => n374_port, 
                           Q => REGISTERS_27_20_port);
   REGISTERS_reg_27_19_inst : DLH_X1 port map( G => n313_port, D => n378_port, 
                           Q => REGISTERS_27_19_port);
   REGISTERS_reg_27_18_inst : DLH_X1 port map( G => n313_port, D => n382_port, 
                           Q => REGISTERS_27_18_port);
   REGISTERS_reg_27_17_inst : DLH_X1 port map( G => n313_port, D => n386_port, 
                           Q => REGISTERS_27_17_port);
   REGISTERS_reg_27_16_inst : DLH_X1 port map( G => n313_port, D => n390_port, 
                           Q => REGISTERS_27_16_port);
   REGISTERS_reg_27_15_inst : DLH_X1 port map( G => n313_port, D => n394_port, 
                           Q => REGISTERS_27_15_port);
   REGISTERS_reg_27_14_inst : DLH_X1 port map( G => n313_port, D => n398_port, 
                           Q => REGISTERS_27_14_port);
   REGISTERS_reg_27_13_inst : DLH_X1 port map( G => n313_port, D => n402_port, 
                           Q => REGISTERS_27_13_port);
   REGISTERS_reg_27_12_inst : DLH_X1 port map( G => n313_port, D => n406_port, 
                           Q => REGISTERS_27_12_port);
   REGISTERS_reg_27_11_inst : DLH_X1 port map( G => n313_port, D => n410_port, 
                           Q => REGISTERS_27_11_port);
   REGISTERS_reg_27_10_inst : DLH_X1 port map( G => n313_port, D => n414_port, 
                           Q => REGISTERS_27_10_port);
   REGISTERS_reg_27_9_inst : DLH_X1 port map( G => n312_port, D => n418_port, Q
                           => REGISTERS_27_9_port);
   REGISTERS_reg_27_8_inst : DLH_X1 port map( G => n312_port, D => n422_port, Q
                           => REGISTERS_27_8_port);
   REGISTERS_reg_27_7_inst : DLH_X1 port map( G => n312_port, D => n426_port, Q
                           => REGISTERS_27_7_port);
   REGISTERS_reg_27_6_inst : DLH_X1 port map( G => n312_port, D => n430_port, Q
                           => REGISTERS_27_6_port);
   REGISTERS_reg_27_5_inst : DLH_X1 port map( G => n312_port, D => n434_port, Q
                           => REGISTERS_27_5_port);
   REGISTERS_reg_27_4_inst : DLH_X1 port map( G => n312_port, D => n438_port, Q
                           => REGISTERS_27_4_port);
   REGISTERS_reg_27_3_inst : DLH_X1 port map( G => n312_port, D => n442, Q => 
                           REGISTERS_27_3_port);
   REGISTERS_reg_27_2_inst : DLH_X1 port map( G => n312_port, D => n446, Q => 
                           REGISTERS_27_2_port);
   REGISTERS_reg_27_1_inst : DLH_X1 port map( G => n312_port, D => n450, Q => 
                           REGISTERS_27_1_port);
   REGISTERS_reg_27_0_inst : DLH_X1 port map( G => n312_port, D => n454, Q => 
                           REGISTERS_27_0_port);
   REGISTERS_reg_28_31_inst : DLH_X1 port map( G => n319_port, D => n330_port, 
                           Q => REGISTERS_28_31_port);
   REGISTERS_reg_28_30_inst : DLH_X1 port map( G => n319_port, D => n334_port, 
                           Q => REGISTERS_28_30_port);
   REGISTERS_reg_28_29_inst : DLH_X1 port map( G => n318_port, D => n338_port, 
                           Q => REGISTERS_28_29_port);
   REGISTERS_reg_28_28_inst : DLH_X1 port map( G => n318_port, D => n342_port, 
                           Q => REGISTERS_28_28_port);
   REGISTERS_reg_28_27_inst : DLH_X1 port map( G => n318_port, D => n346_port, 
                           Q => REGISTERS_28_27_port);
   REGISTERS_reg_28_26_inst : DLH_X1 port map( G => n318_port, D => n350_port, 
                           Q => REGISTERS_28_26_port);
   REGISTERS_reg_28_25_inst : DLH_X1 port map( G => n318_port, D => n354_port, 
                           Q => REGISTERS_28_25_port);
   REGISTERS_reg_28_24_inst : DLH_X1 port map( G => n318_port, D => n358_port, 
                           Q => REGISTERS_28_24_port);
   REGISTERS_reg_28_23_inst : DLH_X1 port map( G => n318_port, D => n362_port, 
                           Q => REGISTERS_28_23_port);
   REGISTERS_reg_28_22_inst : DLH_X1 port map( G => n318_port, D => n366_port, 
                           Q => REGISTERS_28_22_port);
   REGISTERS_reg_28_21_inst : DLH_X1 port map( G => n318_port, D => n370_port, 
                           Q => REGISTERS_28_21_port);
   REGISTERS_reg_28_20_inst : DLH_X1 port map( G => n318_port, D => n374_port, 
                           Q => REGISTERS_28_20_port);
   REGISTERS_reg_28_19_inst : DLH_X1 port map( G => n317_port, D => n378_port, 
                           Q => REGISTERS_28_19_port);
   REGISTERS_reg_28_18_inst : DLH_X1 port map( G => n317_port, D => n382_port, 
                           Q => REGISTERS_28_18_port);
   REGISTERS_reg_28_17_inst : DLH_X1 port map( G => n317_port, D => n386_port, 
                           Q => REGISTERS_28_17_port);
   REGISTERS_reg_28_16_inst : DLH_X1 port map( G => n317_port, D => n390_port, 
                           Q => REGISTERS_28_16_port);
   REGISTERS_reg_28_15_inst : DLH_X1 port map( G => n317_port, D => n394_port, 
                           Q => REGISTERS_28_15_port);
   REGISTERS_reg_28_14_inst : DLH_X1 port map( G => n317_port, D => n398_port, 
                           Q => REGISTERS_28_14_port);
   REGISTERS_reg_28_13_inst : DLH_X1 port map( G => n317_port, D => n402_port, 
                           Q => REGISTERS_28_13_port);
   REGISTERS_reg_28_12_inst : DLH_X1 port map( G => n317_port, D => n406_port, 
                           Q => REGISTERS_28_12_port);
   REGISTERS_reg_28_11_inst : DLH_X1 port map( G => n317_port, D => n410_port, 
                           Q => REGISTERS_28_11_port);
   REGISTERS_reg_28_10_inst : DLH_X1 port map( G => n317_port, D => n414_port, 
                           Q => REGISTERS_28_10_port);
   REGISTERS_reg_28_9_inst : DLH_X1 port map( G => n316_port, D => n418_port, Q
                           => REGISTERS_28_9_port);
   REGISTERS_reg_28_8_inst : DLH_X1 port map( G => n316_port, D => n422_port, Q
                           => REGISTERS_28_8_port);
   REGISTERS_reg_28_7_inst : DLH_X1 port map( G => n316_port, D => n426_port, Q
                           => REGISTERS_28_7_port);
   REGISTERS_reg_28_6_inst : DLH_X1 port map( G => n316_port, D => n430_port, Q
                           => REGISTERS_28_6_port);
   REGISTERS_reg_28_5_inst : DLH_X1 port map( G => n316_port, D => n434_port, Q
                           => REGISTERS_28_5_port);
   REGISTERS_reg_28_4_inst : DLH_X1 port map( G => n316_port, D => n438_port, Q
                           => REGISTERS_28_4_port);
   REGISTERS_reg_28_3_inst : DLH_X1 port map( G => n316_port, D => n442, Q => 
                           REGISTERS_28_3_port);
   REGISTERS_reg_28_2_inst : DLH_X1 port map( G => n316_port, D => n446, Q => 
                           REGISTERS_28_2_port);
   REGISTERS_reg_28_1_inst : DLH_X1 port map( G => n316_port, D => n450, Q => 
                           REGISTERS_28_1_port);
   REGISTERS_reg_28_0_inst : DLH_X1 port map( G => n316_port, D => n454, Q => 
                           REGISTERS_28_0_port);
   REGISTERS_reg_29_31_inst : DLH_X1 port map( G => n323_port, D => n330_port, 
                           Q => REGISTERS_29_31_port);
   REGISTERS_reg_29_30_inst : DLH_X1 port map( G => n323_port, D => n334_port, 
                           Q => REGISTERS_29_30_port);
   REGISTERS_reg_29_29_inst : DLH_X1 port map( G => n322_port, D => n338_port, 
                           Q => REGISTERS_29_29_port);
   REGISTERS_reg_29_28_inst : DLH_X1 port map( G => n322_port, D => n342_port, 
                           Q => REGISTERS_29_28_port);
   REGISTERS_reg_29_27_inst : DLH_X1 port map( G => n322_port, D => n346_port, 
                           Q => REGISTERS_29_27_port);
   REGISTERS_reg_29_26_inst : DLH_X1 port map( G => n322_port, D => n350_port, 
                           Q => REGISTERS_29_26_port);
   REGISTERS_reg_29_25_inst : DLH_X1 port map( G => n322_port, D => n354_port, 
                           Q => REGISTERS_29_25_port);
   REGISTERS_reg_29_24_inst : DLH_X1 port map( G => n322_port, D => n358_port, 
                           Q => REGISTERS_29_24_port);
   REGISTERS_reg_29_23_inst : DLH_X1 port map( G => n322_port, D => n362_port, 
                           Q => REGISTERS_29_23_port);
   REGISTERS_reg_29_22_inst : DLH_X1 port map( G => n322_port, D => n366_port, 
                           Q => REGISTERS_29_22_port);
   REGISTERS_reg_29_21_inst : DLH_X1 port map( G => n322_port, D => n370_port, 
                           Q => REGISTERS_29_21_port);
   REGISTERS_reg_29_20_inst : DLH_X1 port map( G => n322_port, D => n374_port, 
                           Q => REGISTERS_29_20_port);
   REGISTERS_reg_29_19_inst : DLH_X1 port map( G => n321_port, D => n378_port, 
                           Q => REGISTERS_29_19_port);
   REGISTERS_reg_29_18_inst : DLH_X1 port map( G => n321_port, D => n382_port, 
                           Q => REGISTERS_29_18_port);
   REGISTERS_reg_29_17_inst : DLH_X1 port map( G => n321_port, D => n386_port, 
                           Q => REGISTERS_29_17_port);
   REGISTERS_reg_29_16_inst : DLH_X1 port map( G => n321_port, D => n390_port, 
                           Q => REGISTERS_29_16_port);
   REGISTERS_reg_29_15_inst : DLH_X1 port map( G => n321_port, D => n394_port, 
                           Q => REGISTERS_29_15_port);
   REGISTERS_reg_29_14_inst : DLH_X1 port map( G => n321_port, D => n398_port, 
                           Q => REGISTERS_29_14_port);
   REGISTERS_reg_29_13_inst : DLH_X1 port map( G => n321_port, D => n402_port, 
                           Q => REGISTERS_29_13_port);
   REGISTERS_reg_29_12_inst : DLH_X1 port map( G => n321_port, D => n406_port, 
                           Q => REGISTERS_29_12_port);
   REGISTERS_reg_29_11_inst : DLH_X1 port map( G => n321_port, D => n410_port, 
                           Q => REGISTERS_29_11_port);
   REGISTERS_reg_29_10_inst : DLH_X1 port map( G => n321_port, D => n414_port, 
                           Q => REGISTERS_29_10_port);
   REGISTERS_reg_29_9_inst : DLH_X1 port map( G => n320_port, D => n418_port, Q
                           => REGISTERS_29_9_port);
   REGISTERS_reg_29_8_inst : DLH_X1 port map( G => n320_port, D => n422_port, Q
                           => REGISTERS_29_8_port);
   REGISTERS_reg_29_7_inst : DLH_X1 port map( G => n320_port, D => n426_port, Q
                           => REGISTERS_29_7_port);
   REGISTERS_reg_29_6_inst : DLH_X1 port map( G => n320_port, D => n430_port, Q
                           => REGISTERS_29_6_port);
   REGISTERS_reg_29_5_inst : DLH_X1 port map( G => n320_port, D => n434_port, Q
                           => REGISTERS_29_5_port);
   REGISTERS_reg_29_4_inst : DLH_X1 port map( G => n320_port, D => n438_port, Q
                           => REGISTERS_29_4_port);
   REGISTERS_reg_29_3_inst : DLH_X1 port map( G => n320_port, D => n442, Q => 
                           REGISTERS_29_3_port);
   REGISTERS_reg_29_2_inst : DLH_X1 port map( G => n320_port, D => n446, Q => 
                           REGISTERS_29_2_port);
   REGISTERS_reg_29_1_inst : DLH_X1 port map( G => n320_port, D => n450, Q => 
                           REGISTERS_29_1_port);
   REGISTERS_reg_29_0_inst : DLH_X1 port map( G => n320_port, D => n454, Q => 
                           REGISTERS_29_0_port);
   REGISTERS_reg_30_31_inst : DLH_X1 port map( G => n327_port, D => n331_port, 
                           Q => REGISTERS_30_31_port);
   REGISTERS_reg_30_30_inst : DLH_X1 port map( G => n327_port, D => n335_port, 
                           Q => REGISTERS_30_30_port);
   REGISTERS_reg_30_29_inst : DLH_X1 port map( G => n326_port, D => n339_port, 
                           Q => REGISTERS_30_29_port);
   REGISTERS_reg_30_28_inst : DLH_X1 port map( G => n326_port, D => n343_port, 
                           Q => REGISTERS_30_28_port);
   REGISTERS_reg_30_27_inst : DLH_X1 port map( G => n326_port, D => n347_port, 
                           Q => REGISTERS_30_27_port);
   REGISTERS_reg_30_26_inst : DLH_X1 port map( G => n326_port, D => n351_port, 
                           Q => REGISTERS_30_26_port);
   REGISTERS_reg_30_25_inst : DLH_X1 port map( G => n326_port, D => n355_port, 
                           Q => REGISTERS_30_25_port);
   REGISTERS_reg_30_24_inst : DLH_X1 port map( G => n326_port, D => n359_port, 
                           Q => REGISTERS_30_24_port);
   REGISTERS_reg_30_23_inst : DLH_X1 port map( G => n326_port, D => n363_port, 
                           Q => REGISTERS_30_23_port);
   REGISTERS_reg_30_22_inst : DLH_X1 port map( G => n326_port, D => n367_port, 
                           Q => REGISTERS_30_22_port);
   REGISTERS_reg_30_21_inst : DLH_X1 port map( G => n326_port, D => n371_port, 
                           Q => REGISTERS_30_21_port);
   REGISTERS_reg_30_20_inst : DLH_X1 port map( G => n326_port, D => n375_port, 
                           Q => REGISTERS_30_20_port);
   REGISTERS_reg_30_19_inst : DLH_X1 port map( G => n325_port, D => n379_port, 
                           Q => REGISTERS_30_19_port);
   REGISTERS_reg_30_18_inst : DLH_X1 port map( G => n325_port, D => n383_port, 
                           Q => REGISTERS_30_18_port);
   REGISTERS_reg_30_17_inst : DLH_X1 port map( G => n325_port, D => n387_port, 
                           Q => REGISTERS_30_17_port);
   REGISTERS_reg_30_16_inst : DLH_X1 port map( G => n325_port, D => n391_port, 
                           Q => REGISTERS_30_16_port);
   REGISTERS_reg_30_15_inst : DLH_X1 port map( G => n325_port, D => n395_port, 
                           Q => REGISTERS_30_15_port);
   REGISTERS_reg_30_14_inst : DLH_X1 port map( G => n325_port, D => n399_port, 
                           Q => REGISTERS_30_14_port);
   REGISTERS_reg_30_13_inst : DLH_X1 port map( G => n325_port, D => n403_port, 
                           Q => REGISTERS_30_13_port);
   REGISTERS_reg_30_12_inst : DLH_X1 port map( G => n325_port, D => n407_port, 
                           Q => REGISTERS_30_12_port);
   REGISTERS_reg_30_11_inst : DLH_X1 port map( G => n325_port, D => n411_port, 
                           Q => REGISTERS_30_11_port);
   REGISTERS_reg_30_10_inst : DLH_X1 port map( G => n325_port, D => n415_port, 
                           Q => REGISTERS_30_10_port);
   REGISTERS_reg_30_9_inst : DLH_X1 port map( G => n324_port, D => n419_port, Q
                           => REGISTERS_30_9_port);
   REGISTERS_reg_30_8_inst : DLH_X1 port map( G => n324_port, D => n423_port, Q
                           => REGISTERS_30_8_port);
   REGISTERS_reg_30_7_inst : DLH_X1 port map( G => n324_port, D => n427_port, Q
                           => REGISTERS_30_7_port);
   REGISTERS_reg_30_6_inst : DLH_X1 port map( G => n324_port, D => n431_port, Q
                           => REGISTERS_30_6_port);
   REGISTERS_reg_30_5_inst : DLH_X1 port map( G => n324_port, D => n435_port, Q
                           => REGISTERS_30_5_port);
   REGISTERS_reg_30_4_inst : DLH_X1 port map( G => n324_port, D => n439_port, Q
                           => REGISTERS_30_4_port);
   REGISTERS_reg_30_3_inst : DLH_X1 port map( G => n324_port, D => n443, Q => 
                           REGISTERS_30_3_port);
   REGISTERS_reg_30_2_inst : DLH_X1 port map( G => n324_port, D => n447, Q => 
                           REGISTERS_30_2_port);
   REGISTERS_reg_30_1_inst : DLH_X1 port map( G => n324_port, D => n451, Q => 
                           REGISTERS_30_1_port);
   REGISTERS_reg_30_0_inst : DLH_X1 port map( G => n324_port, D => n455, Q => 
                           REGISTERS_30_0_port);
   REGISTERS_reg_31_31_inst : DLH_X1 port map( G => n459, D => n331_port, Q => 
                           REGISTERS_31_31_port);
   REGISTERS_reg_31_30_inst : DLH_X1 port map( G => n459, D => n335_port, Q => 
                           REGISTERS_31_30_port);
   REGISTERS_reg_31_29_inst : DLH_X1 port map( G => n458, D => n339_port, Q => 
                           REGISTERS_31_29_port);
   REGISTERS_reg_31_28_inst : DLH_X1 port map( G => n458, D => n343_port, Q => 
                           REGISTERS_31_28_port);
   REGISTERS_reg_31_27_inst : DLH_X1 port map( G => n458, D => n347_port, Q => 
                           REGISTERS_31_27_port);
   REGISTERS_reg_31_26_inst : DLH_X1 port map( G => n458, D => n351_port, Q => 
                           REGISTERS_31_26_port);
   REGISTERS_reg_31_25_inst : DLH_X1 port map( G => n458, D => n355_port, Q => 
                           REGISTERS_31_25_port);
   REGISTERS_reg_31_24_inst : DLH_X1 port map( G => n458, D => n359_port, Q => 
                           REGISTERS_31_24_port);
   REGISTERS_reg_31_23_inst : DLH_X1 port map( G => n458, D => n363_port, Q => 
                           REGISTERS_31_23_port);
   REGISTERS_reg_31_22_inst : DLH_X1 port map( G => n458, D => n367_port, Q => 
                           REGISTERS_31_22_port);
   REGISTERS_reg_31_21_inst : DLH_X1 port map( G => n458, D => n371_port, Q => 
                           REGISTERS_31_21_port);
   REGISTERS_reg_31_20_inst : DLH_X1 port map( G => n458, D => n375_port, Q => 
                           REGISTERS_31_20_port);
   REGISTERS_reg_31_19_inst : DLH_X1 port map( G => n457, D => n379_port, Q => 
                           REGISTERS_31_19_port);
   REGISTERS_reg_31_18_inst : DLH_X1 port map( G => n457, D => n383_port, Q => 
                           REGISTERS_31_18_port);
   REGISTERS_reg_31_17_inst : DLH_X1 port map( G => n457, D => n387_port, Q => 
                           REGISTERS_31_17_port);
   REGISTERS_reg_31_16_inst : DLH_X1 port map( G => n457, D => n391_port, Q => 
                           REGISTERS_31_16_port);
   REGISTERS_reg_31_15_inst : DLH_X1 port map( G => n457, D => n395_port, Q => 
                           REGISTERS_31_15_port);
   REGISTERS_reg_31_14_inst : DLH_X1 port map( G => n457, D => n399_port, Q => 
                           REGISTERS_31_14_port);
   REGISTERS_reg_31_13_inst : DLH_X1 port map( G => n457, D => n403_port, Q => 
                           REGISTERS_31_13_port);
   REGISTERS_reg_31_12_inst : DLH_X1 port map( G => n457, D => n407_port, Q => 
                           REGISTERS_31_12_port);
   REGISTERS_reg_31_11_inst : DLH_X1 port map( G => n457, D => n411_port, Q => 
                           REGISTERS_31_11_port);
   REGISTERS_reg_31_10_inst : DLH_X1 port map( G => n457, D => n415_port, Q => 
                           REGISTERS_31_10_port);
   REGISTERS_reg_31_9_inst : DLH_X1 port map( G => n456, D => n419_port, Q => 
                           REGISTERS_31_9_port);
   REGISTERS_reg_31_8_inst : DLH_X1 port map( G => n456, D => n423_port, Q => 
                           REGISTERS_31_8_port);
   REGISTERS_reg_31_7_inst : DLH_X1 port map( G => n456, D => n427_port, Q => 
                           REGISTERS_31_7_port);
   REGISTERS_reg_31_6_inst : DLH_X1 port map( G => n456, D => n431_port, Q => 
                           REGISTERS_31_6_port);
   REGISTERS_reg_31_5_inst : DLH_X1 port map( G => n456, D => n435_port, Q => 
                           REGISTERS_31_5_port);
   REGISTERS_reg_31_4_inst : DLH_X1 port map( G => n456, D => n439_port, Q => 
                           REGISTERS_31_4_port);
   REGISTERS_reg_31_3_inst : DLH_X1 port map( G => n456, D => n443, Q => 
                           REGISTERS_31_3_port);
   REGISTERS_reg_31_2_inst : DLH_X1 port map( G => n456, D => n447, Q => 
                           REGISTERS_31_2_port);
   REGISTERS_reg_31_1_inst : DLH_X1 port map( G => n456, D => n451, Q => 
                           REGISTERS_31_1_port);
   REGISTERS_reg_31_0_inst : DLH_X1 port map( G => n456, D => n455, Q => 
                           REGISTERS_31_0_port);
   OUT1_reg_31_inst : DLH_X1 port map( G => n200, D => N408, Q => OUT1(31));
   OUT1_reg_30_inst : DLH_X1 port map( G => n200, D => N407, Q => OUT1(30));
   OUT1_reg_29_inst : DLH_X1 port map( G => n200, D => N406, Q => OUT1(29));
   OUT1_reg_28_inst : DLH_X1 port map( G => n200, D => N405, Q => OUT1(28));
   OUT1_reg_27_inst : DLH_X1 port map( G => n200, D => N404, Q => OUT1(27));
   OUT1_reg_26_inst : DLH_X1 port map( G => n200, D => N403, Q => OUT1(26));
   OUT1_reg_25_inst : DLH_X1 port map( G => n200, D => N402, Q => OUT1(25));
   OUT1_reg_24_inst : DLH_X1 port map( G => n200, D => N401, Q => OUT1(24));
   OUT1_reg_23_inst : DLH_X1 port map( G => n200, D => N400, Q => OUT1(23));
   OUT1_reg_22_inst : DLH_X1 port map( G => n200, D => N399, Q => OUT1(22));
   OUT1_reg_21_inst : DLH_X1 port map( G => n201, D => N398, Q => OUT1(21));
   OUT1_reg_20_inst : DLH_X1 port map( G => n201, D => N397, Q => OUT1(20));
   OUT1_reg_19_inst : DLH_X1 port map( G => n201, D => N396, Q => OUT1(19));
   OUT1_reg_18_inst : DLH_X1 port map( G => n201, D => N395, Q => OUT1(18));
   OUT1_reg_17_inst : DLH_X1 port map( G => n201, D => N394, Q => OUT1(17));
   OUT1_reg_16_inst : DLH_X1 port map( G => n201, D => N393, Q => OUT1(16));
   OUT1_reg_15_inst : DLH_X1 port map( G => n201, D => N392, Q => OUT1(15));
   OUT1_reg_14_inst : DLH_X1 port map( G => n201, D => N391, Q => OUT1(14));
   OUT1_reg_13_inst : DLH_X1 port map( G => n201, D => N390, Q => OUT1(13));
   OUT1_reg_12_inst : DLH_X1 port map( G => n201, D => N389, Q => OUT1(12));
   OUT1_reg_11_inst : DLH_X1 port map( G => n202, D => N388, Q => OUT1(11));
   OUT1_reg_10_inst : DLH_X1 port map( G => n202, D => N387, Q => OUT1(10));
   OUT1_reg_9_inst : DLH_X1 port map( G => n202, D => N386, Q => OUT1(9));
   OUT1_reg_8_inst : DLH_X1 port map( G => n202, D => N385, Q => OUT1(8));
   OUT1_reg_7_inst : DLH_X1 port map( G => n202, D => N384, Q => OUT1(7));
   OUT1_reg_6_inst : DLH_X1 port map( G => n202, D => N383, Q => OUT1(6));
   OUT1_reg_5_inst : DLH_X1 port map( G => n202, D => N382, Q => OUT1(5));
   OUT1_reg_4_inst : DLH_X1 port map( G => n202, D => N381, Q => OUT1(4));
   OUT1_reg_3_inst : DLH_X1 port map( G => n202, D => N380, Q => OUT1(3));
   OUT1_reg_2_inst : DLH_X1 port map( G => n202, D => N379, Q => OUT1(2));
   OUT1_reg_1_inst : DLH_X1 port map( G => n203, D => N378, Q => OUT1(1));
   OUT1_reg_0_inst : DLH_X1 port map( G => n203, D => N377, Q => OUT1(0));
   OUT2_reg_31_inst : DLH_X1 port map( G => n196, D => N441, Q => OUT2(31));
   OUT2_reg_30_inst : DLH_X1 port map( G => n196, D => N440, Q => OUT2(30));
   OUT2_reg_29_inst : DLH_X1 port map( G => n196, D => N439, Q => OUT2(29));
   OUT2_reg_28_inst : DLH_X1 port map( G => n196, D => N438, Q => OUT2(28));
   OUT2_reg_27_inst : DLH_X1 port map( G => n196, D => N437, Q => OUT2(27));
   OUT2_reg_26_inst : DLH_X1 port map( G => n196, D => N436, Q => OUT2(26));
   OUT2_reg_25_inst : DLH_X1 port map( G => n196, D => N435, Q => OUT2(25));
   OUT2_reg_24_inst : DLH_X1 port map( G => n196, D => N434, Q => OUT2(24));
   OUT2_reg_23_inst : DLH_X1 port map( G => n196, D => N433, Q => OUT2(23));
   OUT2_reg_22_inst : DLH_X1 port map( G => n196, D => N432, Q => OUT2(22));
   OUT2_reg_21_inst : DLH_X1 port map( G => n197, D => N431, Q => OUT2(21));
   OUT2_reg_20_inst : DLH_X1 port map( G => n197, D => N430, Q => OUT2(20));
   OUT2_reg_19_inst : DLH_X1 port map( G => n197, D => N429, Q => OUT2(19));
   OUT2_reg_18_inst : DLH_X1 port map( G => n197, D => N428, Q => OUT2(18));
   OUT2_reg_17_inst : DLH_X1 port map( G => n197, D => N427, Q => OUT2(17));
   OUT2_reg_16_inst : DLH_X1 port map( G => n197, D => N426, Q => OUT2(16));
   OUT2_reg_15_inst : DLH_X1 port map( G => n197, D => N425, Q => OUT2(15));
   OUT2_reg_14_inst : DLH_X1 port map( G => n197, D => N424, Q => OUT2(14));
   OUT2_reg_13_inst : DLH_X1 port map( G => n197, D => N423, Q => OUT2(13));
   OUT2_reg_12_inst : DLH_X1 port map( G => n197, D => N422, Q => OUT2(12));
   OUT2_reg_11_inst : DLH_X1 port map( G => n198, D => N421, Q => OUT2(11));
   OUT2_reg_10_inst : DLH_X1 port map( G => n198, D => N420, Q => OUT2(10));
   OUT2_reg_9_inst : DLH_X1 port map( G => n198, D => N419, Q => OUT2(9));
   OUT2_reg_8_inst : DLH_X1 port map( G => n198, D => N418, Q => OUT2(8));
   OUT2_reg_7_inst : DLH_X1 port map( G => n198, D => N417, Q => OUT2(7));
   OUT2_reg_6_inst : DLH_X1 port map( G => n198, D => N416, Q => OUT2(6));
   OUT2_reg_5_inst : DLH_X1 port map( G => n198, D => N415, Q => OUT2(5));
   OUT2_reg_4_inst : DLH_X1 port map( G => n198, D => N414, Q => OUT2(4));
   OUT2_reg_3_inst : DLH_X1 port map( G => n198, D => N413, Q => OUT2(3));
   OUT2_reg_2_inst : DLH_X1 port map( G => n198, D => N412, Q => OUT2(2));
   OUT2_reg_1_inst : DLH_X1 port map( G => n199, D => N411, Q => OUT2(1));
   OUT2_reg_0_inst : DLH_X1 port map( G => n199, D => N410, Q => OUT2(0));
   U1911 : NAND3_X1 port map( A1 => n2262, A2 => n2263, A3 => WR, ZN => n1778);
   U1912 : NAND3_X1 port map( A1 => WR, A2 => n2263, A3 => ADD_WR(3), ZN => 
                           n1787);
   U1913 : NAND3_X1 port map( A1 => WR, A2 => n2262, A3 => ADD_WR(4), ZN => 
                           n1788);
   U1914 : NAND3_X1 port map( A1 => n2260, A2 => n2261, A3 => ADD_WR(0), ZN => 
                           n1779);
   U1915 : NAND3_X1 port map( A1 => n2259, A2 => n2261, A3 => ADD_WR(1), ZN => 
                           n1780);
   U1916 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n2261, A3 => ADD_WR(1), ZN
                           => n1781);
   U1917 : NAND3_X1 port map( A1 => n2259, A2 => n2260, A3 => ADD_WR(2), ZN => 
                           n1782);
   U1918 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n2260, A3 => ADD_WR(2), ZN
                           => n1783);
   U1919 : NAND3_X1 port map( A1 => ADD_WR(1), A2 => n2259, A3 => ADD_WR(2), ZN
                           => n1784);
   U1920 : NAND3_X1 port map( A1 => n2260, A2 => n2261, A3 => n2259, ZN => 
                           n1786);
   U1921 : NAND3_X1 port map( A1 => ADD_WR(3), A2 => WR, A3 => ADD_WR(4), ZN =>
                           n1789);
   U1922 : NAND3_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(0), A3 => ADD_WR(2)
                           , ZN => n1785);
   U3 : NOR2_X1 port map( A1 => n2253, A2 => ADD_RD2(1), ZN => n1130);
   U4 : NOR2_X1 port map( A1 => n2257, A2 => ADD_RD1(1), ZN => n1755);
   U5 : NOR2_X1 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(2), ZN => n1127);
   U6 : BUF_X1 port map( A => n549, Z => n154);
   U7 : BUF_X1 port map( A => n549, Z => n155);
   U8 : BUF_X1 port map( A => n1167, Z => n76);
   U9 : BUF_X1 port map( A => n1191, Z => n28);
   U10 : BUF_X1 port map( A => n1201, Z => n4);
   U11 : BUF_X1 port map( A => n1167, Z => n77);
   U12 : BUF_X1 port map( A => n1191, Z => n29);
   U13 : BUF_X1 port map( A => n1201, Z => n5);
   U14 : BUF_X1 port map( A => n1174, Z => n60);
   U15 : BUF_X1 port map( A => n542, Z => n172);
   U16 : BUF_X1 port map( A => n566, Z => n124);
   U17 : BUF_X1 port map( A => n576, Z => n100);
   U18 : BUF_X1 port map( A => n542, Z => n173);
   U19 : BUF_X1 port map( A => n566, Z => n125);
   U20 : BUF_X1 port map( A => n576, Z => n101);
   U21 : BUF_X1 port map( A => n549, Z => n156);
   U22 : BUF_X1 port map( A => n1167, Z => n78);
   U23 : BUF_X1 port map( A => n1191, Z => n30);
   U24 : BUF_X1 port map( A => n1201, Z => n6);
   U25 : BUF_X1 port map( A => n542, Z => n174);
   U26 : BUF_X1 port map( A => n566, Z => n126);
   U27 : BUF_X1 port map( A => n576, Z => n102);
   U28 : BUF_X1 port map( A => n1174, Z => n58);
   U29 : BUF_X1 port map( A => n1174, Z => n59);
   U30 : INV_X1 port map( A => n473, ZN => n462);
   U31 : INV_X1 port map( A => n473, ZN => n463);
   U32 : INV_X1 port map( A => n473, ZN => n464);
   U33 : BUF_X1 port map( A => n1161, Z => n91);
   U34 : BUF_X1 port map( A => n1166, Z => n79);
   U35 : BUF_X1 port map( A => n1171, Z => n67);
   U36 : BUF_X1 port map( A => n1176, Z => n55);
   U37 : BUF_X1 port map( A => n1185, Z => n43);
   U38 : BUF_X1 port map( A => n1190, Z => n31);
   U39 : BUF_X1 port map( A => n1195, Z => n19);
   U40 : BUF_X1 port map( A => n1200, Z => n7);
   U41 : BUF_X1 port map( A => n1161, Z => n92);
   U42 : BUF_X1 port map( A => n1166, Z => n80);
   U43 : BUF_X1 port map( A => n1171, Z => n68);
   U44 : BUF_X1 port map( A => n1176, Z => n56);
   U45 : BUF_X1 port map( A => n1185, Z => n44);
   U46 : BUF_X1 port map( A => n1190, Z => n32);
   U47 : BUF_X1 port map( A => n1195, Z => n20);
   U48 : BUF_X1 port map( A => n1200, Z => n8);
   U49 : BUF_X1 port map( A => n1158, Z => n97);
   U50 : BUF_X1 port map( A => n1182, Z => n49);
   U51 : BUF_X1 port map( A => n1192, Z => n25);
   U52 : BUF_X1 port map( A => n1168, Z => n73);
   U53 : BUF_X1 port map( A => n1163, Z => n85);
   U54 : BUF_X1 port map( A => n1187, Z => n37);
   U55 : BUF_X1 port map( A => n1197, Z => n13);
   U56 : BUF_X1 port map( A => n1173, Z => n61);
   U57 : BUF_X1 port map( A => n534, Z => n190);
   U58 : BUF_X1 port map( A => n539, Z => n178);
   U59 : BUF_X1 port map( A => n544, Z => n166);
   U60 : BUF_X1 port map( A => n558, Z => n142);
   U61 : BUF_X1 port map( A => n563, Z => n130);
   U62 : BUF_X1 port map( A => n568, Z => n118);
   U63 : BUF_X1 port map( A => n573, Z => n106);
   U64 : BUF_X1 port map( A => n534, Z => n191);
   U65 : BUF_X1 port map( A => n539, Z => n179);
   U66 : BUF_X1 port map( A => n544, Z => n167);
   U67 : BUF_X1 port map( A => n558, Z => n143);
   U68 : BUF_X1 port map( A => n563, Z => n131);
   U69 : BUF_X1 port map( A => n568, Z => n119);
   U70 : BUF_X1 port map( A => n573, Z => n107);
   U71 : BUF_X1 port map( A => n1162, Z => n88);
   U72 : BUF_X1 port map( A => n1172, Z => n64);
   U73 : BUF_X1 port map( A => n1177, Z => n52);
   U74 : BUF_X1 port map( A => n1186, Z => n40);
   U75 : BUF_X1 port map( A => n1196, Z => n16);
   U76 : BUF_X1 port map( A => n1162, Z => n89);
   U77 : BUF_X1 port map( A => n1172, Z => n65);
   U78 : BUF_X1 port map( A => n1177, Z => n53);
   U79 : BUF_X1 port map( A => n1186, Z => n41);
   U80 : BUF_X1 port map( A => n1196, Z => n17);
   U81 : BUF_X1 port map( A => n1159, Z => n96);
   U82 : BUF_X1 port map( A => n1183, Z => n48);
   U83 : BUF_X1 port map( A => n1193, Z => n24);
   U84 : BUF_X1 port map( A => n1169, Z => n72);
   U85 : BUF_X1 port map( A => n1164, Z => n84);
   U86 : BUF_X1 port map( A => n1188, Z => n36);
   U87 : BUF_X1 port map( A => n1198, Z => n12);
   U88 : BUF_X1 port map( A => n1161, Z => n93);
   U89 : BUF_X1 port map( A => n1171, Z => n69);
   U90 : BUF_X1 port map( A => n1166, Z => n81);
   U91 : BUF_X1 port map( A => n1176, Z => n57);
   U92 : BUF_X1 port map( A => n1185, Z => n45);
   U93 : BUF_X1 port map( A => n1190, Z => n33);
   U94 : BUF_X1 port map( A => n1195, Z => n21);
   U95 : BUF_X1 port map( A => n1200, Z => n9);
   U96 : BUF_X1 port map( A => n1158, Z => n99);
   U97 : BUF_X1 port map( A => n1182, Z => n51);
   U98 : BUF_X1 port map( A => n1192, Z => n27);
   U99 : BUF_X1 port map( A => n1168, Z => n75);
   U100 : BUF_X1 port map( A => n1163, Z => n87);
   U101 : BUF_X1 port map( A => n1187, Z => n39);
   U102 : BUF_X1 port map( A => n1197, Z => n15);
   U103 : BUF_X1 port map( A => n1173, Z => n63);
   U104 : BUF_X1 port map( A => n533, Z => n193);
   U105 : BUF_X1 port map( A => n557, Z => n145);
   U106 : BUF_X1 port map( A => n567, Z => n121);
   U107 : BUF_X1 port map( A => n533, Z => n194);
   U108 : BUF_X1 port map( A => n557, Z => n146);
   U109 : BUF_X1 port map( A => n567, Z => n122);
   U110 : BUF_X1 port map( A => n538, Z => n181);
   U111 : BUF_X1 port map( A => n562, Z => n133);
   U112 : BUF_X1 port map( A => n572, Z => n109);
   U113 : BUF_X1 port map( A => n538, Z => n182);
   U114 : BUF_X1 port map( A => n562, Z => n134);
   U115 : BUF_X1 port map( A => n572, Z => n110);
   U116 : BUF_X1 port map( A => n543, Z => n169);
   U117 : BUF_X1 port map( A => n543, Z => n170);
   U118 : BUF_X1 port map( A => n536, Z => n187);
   U119 : BUF_X1 port map( A => n541, Z => n175);
   U120 : BUF_X1 port map( A => n546, Z => n163);
   U121 : BUF_X1 port map( A => n551, Z => n151);
   U122 : BUF_X1 port map( A => n560, Z => n139);
   U123 : BUF_X1 port map( A => n565, Z => n127);
   U124 : BUF_X1 port map( A => n570, Z => n115);
   U125 : BUF_X1 port map( A => n575, Z => n103);
   U126 : BUF_X1 port map( A => n536, Z => n188);
   U127 : BUF_X1 port map( A => n541, Z => n176);
   U128 : BUF_X1 port map( A => n546, Z => n164);
   U129 : BUF_X1 port map( A => n551, Z => n152);
   U130 : BUF_X1 port map( A => n560, Z => n140);
   U131 : BUF_X1 port map( A => n565, Z => n128);
   U132 : BUF_X1 port map( A => n570, Z => n116);
   U133 : BUF_X1 port map( A => n575, Z => n104);
   U134 : BUF_X1 port map( A => n548, Z => n157);
   U135 : BUF_X1 port map( A => n548, Z => n158);
   U136 : BUF_X1 port map( A => n537, Z => n184);
   U137 : BUF_X1 port map( A => n547, Z => n160);
   U138 : BUF_X1 port map( A => n552, Z => n148);
   U139 : BUF_X1 port map( A => n561, Z => n136);
   U140 : BUF_X1 port map( A => n571, Z => n112);
   U141 : BUF_X1 port map( A => n537, Z => n185);
   U142 : BUF_X1 port map( A => n547, Z => n161);
   U143 : BUF_X1 port map( A => n552, Z => n149);
   U144 : BUF_X1 port map( A => n561, Z => n137);
   U145 : BUF_X1 port map( A => n571, Z => n113);
   U146 : BUF_X1 port map( A => n534, Z => n192);
   U147 : BUF_X1 port map( A => n539, Z => n180);
   U148 : BUF_X1 port map( A => n544, Z => n168);
   U149 : BUF_X1 port map( A => n558, Z => n144);
   U150 : BUF_X1 port map( A => n563, Z => n132);
   U151 : BUF_X1 port map( A => n568, Z => n120);
   U152 : BUF_X1 port map( A => n573, Z => n108);
   U153 : BUF_X1 port map( A => n1162, Z => n90);
   U154 : BUF_X1 port map( A => n1172, Z => n66);
   U155 : BUF_X1 port map( A => n1177, Z => n54);
   U156 : BUF_X1 port map( A => n1186, Z => n42);
   U157 : BUF_X1 port map( A => n1196, Z => n18);
   U158 : BUF_X1 port map( A => n533, Z => n195);
   U159 : BUF_X1 port map( A => n557, Z => n147);
   U160 : BUF_X1 port map( A => n567, Z => n123);
   U161 : BUF_X1 port map( A => n538, Z => n183);
   U162 : BUF_X1 port map( A => n562, Z => n135);
   U163 : BUF_X1 port map( A => n572, Z => n111);
   U164 : BUF_X1 port map( A => n543, Z => n171);
   U165 : BUF_X1 port map( A => n536, Z => n189);
   U166 : BUF_X1 port map( A => n541, Z => n177);
   U167 : BUF_X1 port map( A => n546, Z => n165);
   U168 : BUF_X1 port map( A => n551, Z => n153);
   U169 : BUF_X1 port map( A => n560, Z => n141);
   U170 : BUF_X1 port map( A => n565, Z => n129);
   U171 : BUF_X1 port map( A => n570, Z => n117);
   U172 : BUF_X1 port map( A => n575, Z => n105);
   U173 : BUF_X1 port map( A => n548, Z => n159);
   U174 : BUF_X1 port map( A => n537, Z => n186);
   U175 : BUF_X1 port map( A => n547, Z => n162);
   U176 : BUF_X1 port map( A => n552, Z => n150);
   U177 : BUF_X1 port map( A => n561, Z => n138);
   U178 : BUF_X1 port map( A => n571, Z => n114);
   U179 : BUF_X1 port map( A => n1159, Z => n94);
   U180 : BUF_X1 port map( A => n1183, Z => n46);
   U181 : BUF_X1 port map( A => n1193, Z => n22);
   U182 : BUF_X1 port map( A => n1159, Z => n95);
   U183 : BUF_X1 port map( A => n1183, Z => n47);
   U184 : BUF_X1 port map( A => n1193, Z => n23);
   U185 : BUF_X1 port map( A => n1169, Z => n70);
   U186 : BUF_X1 port map( A => n1169, Z => n71);
   U187 : BUF_X1 port map( A => n1164, Z => n82);
   U188 : BUF_X1 port map( A => n1188, Z => n34);
   U189 : BUF_X1 port map( A => n1198, Z => n10);
   U190 : BUF_X1 port map( A => n1164, Z => n83);
   U191 : BUF_X1 port map( A => n1188, Z => n35);
   U192 : BUF_X1 port map( A => n1198, Z => n11);
   U193 : BUF_X1 port map( A => n1158, Z => n98);
   U194 : BUF_X1 port map( A => n1182, Z => n50);
   U195 : BUF_X1 port map( A => n1192, Z => n26);
   U196 : BUF_X1 port map( A => n1168, Z => n74);
   U197 : BUF_X1 port map( A => n1163, Z => n86);
   U198 : BUF_X1 port map( A => n1173, Z => n62);
   U199 : BUF_X1 port map( A => n1187, Z => n38);
   U200 : BUF_X1 port map( A => n1197, Z => n14);
   U201 : NAND2_X1 port map( A1 => n1758, A2 => n1754, ZN => n1174);
   U202 : AND2_X1 port map( A1 => n1124, A2 => n1129, ZN => n542);
   U203 : AND2_X1 port map( A1 => n1142, A2 => n1129, ZN => n566);
   U204 : AND2_X1 port map( A1 => n1147, A2 => n1129, ZN => n576);
   U205 : NAND2_X1 port map( A1 => n1133, A2 => n1129, ZN => n549);
   U206 : AND2_X1 port map( A1 => n1749, A2 => n1754, ZN => n1167);
   U207 : AND2_X1 port map( A1 => n1767, A2 => n1754, ZN => n1191);
   U208 : AND2_X1 port map( A1 => n1772, A2 => n1754, ZN => n1201);
   U209 : NOR2_X1 port map( A1 => n2253, A2 => n2252, ZN => n1129);
   U210 : NOR2_X1 port map( A1 => n2257, A2 => n2256, ZN => n1754);
   U211 : NAND2_X1 port map( A1 => n1752, A2 => n1758, ZN => n1169);
   U212 : NAND2_X1 port map( A1 => n1752, A2 => n1759, ZN => n1168);
   U213 : NAND2_X1 port map( A1 => n1749, A2 => n1752, ZN => n1159);
   U214 : NAND2_X1 port map( A1 => n1767, A2 => n1752, ZN => n1183);
   U215 : NAND2_X1 port map( A1 => n1772, A2 => n1752, ZN => n1193);
   U216 : NAND2_X1 port map( A1 => n1751, A2 => n1752, ZN => n1158);
   U217 : NAND2_X1 port map( A1 => n1768, A2 => n1752, ZN => n1182);
   U218 : NAND2_X1 port map( A1 => n1773, A2 => n1752, ZN => n1192);
   U219 : NAND2_X1 port map( A1 => n1127, A2 => n1134, ZN => n543);
   U220 : NAND2_X1 port map( A1 => n1127, A2 => n1133, ZN => n544);
   U221 : NAND2_X1 port map( A1 => n1129, A2 => n1134, ZN => n548);
   U222 : NAND2_X1 port map( A1 => n1126, A2 => n1127, ZN => n533);
   U223 : NAND2_X1 port map( A1 => n1143, A2 => n1127, ZN => n557);
   U224 : NAND2_X1 port map( A1 => n1148, A2 => n1127, ZN => n567);
   U225 : NAND2_X1 port map( A1 => n1754, A2 => n1759, ZN => n1173);
   U226 : NAND2_X1 port map( A1 => n1126, A2 => n1130, ZN => n538);
   U227 : NAND2_X1 port map( A1 => n1143, A2 => n1130, ZN => n562);
   U228 : NAND2_X1 port map( A1 => n1148, A2 => n1130, ZN => n572);
   U229 : NAND2_X1 port map( A1 => n1749, A2 => n1755, ZN => n1164);
   U230 : NAND2_X1 port map( A1 => n1767, A2 => n1755, ZN => n1188);
   U231 : NAND2_X1 port map( A1 => n1772, A2 => n1755, ZN => n1198);
   U232 : NAND2_X1 port map( A1 => n1751, A2 => n1755, ZN => n1163);
   U233 : NAND2_X1 port map( A1 => n1768, A2 => n1755, ZN => n1187);
   U234 : NAND2_X1 port map( A1 => n1773, A2 => n1755, ZN => n1197);
   U235 : BUF_X1 port map( A => n461, Z => n473);
   U236 : NAND2_X1 port map( A1 => n1124, A2 => n1127, ZN => n534);
   U237 : NAND2_X1 port map( A1 => n1142, A2 => n1127, ZN => n558);
   U238 : NAND2_X1 port map( A1 => n1147, A2 => n1127, ZN => n568);
   U239 : AND2_X1 port map( A1 => n1136, A2 => n2251, ZN => n1133);
   U240 : AND2_X1 port map( A1 => n1761, A2 => n2255, ZN => n1758);
   U241 : AND2_X1 port map( A1 => n1145, A2 => n2251, ZN => n1142);
   U242 : AND2_X1 port map( A1 => n1150, A2 => n2251, ZN => n1147);
   U243 : AND2_X1 port map( A1 => n1770, A2 => n2255, ZN => n1767);
   U244 : AND2_X1 port map( A1 => n1775, A2 => n2255, ZN => n1772);
   U245 : AND2_X1 port map( A1 => n1131, A2 => n2251, ZN => n1124);
   U246 : AND2_X1 port map( A1 => n1756, A2 => n2255, ZN => n1749);
   U247 : NAND2_X1 port map( A1 => n1124, A2 => n1130, ZN => n539);
   U248 : NAND2_X1 port map( A1 => n1142, A2 => n1130, ZN => n563);
   U249 : NAND2_X1 port map( A1 => n1147, A2 => n1130, ZN => n573);
   U250 : AND2_X1 port map( A1 => n1130, A2 => n1134, ZN => n551);
   U251 : AND2_X1 port map( A1 => n1130, A2 => n1133, ZN => n552);
   U252 : AND2_X1 port map( A1 => n1125, A2 => n1134, ZN => n546);
   U253 : AND2_X1 port map( A1 => n1125, A2 => n1133, ZN => n547);
   U254 : AND2_X1 port map( A1 => n1126, A2 => n1129, ZN => n541);
   U255 : AND2_X1 port map( A1 => n1143, A2 => n1129, ZN => n565);
   U256 : AND2_X1 port map( A1 => n1148, A2 => n1129, ZN => n575);
   U257 : AND2_X1 port map( A1 => n1126, A2 => n1125, ZN => n536);
   U258 : AND2_X1 port map( A1 => n1124, A2 => n1125, ZN => n537);
   U259 : AND2_X1 port map( A1 => n1143, A2 => n1125, ZN => n560);
   U260 : AND2_X1 port map( A1 => n1142, A2 => n1125, ZN => n561);
   U261 : AND2_X1 port map( A1 => n1148, A2 => n1125, ZN => n570);
   U262 : AND2_X1 port map( A1 => n1147, A2 => n1125, ZN => n571);
   U263 : BUF_X1 port map( A => n461, Z => n471);
   U264 : BUF_X1 port map( A => n461, Z => n470);
   U265 : BUF_X1 port map( A => n460, Z => n469);
   U266 : BUF_X1 port map( A => n460, Z => n468);
   U267 : BUF_X1 port map( A => n460, Z => n467);
   U268 : BUF_X1 port map( A => n460, Z => n466);
   U269 : BUF_X1 port map( A => n460, Z => n465);
   U270 : BUF_X1 port map( A => n461, Z => n472);
   U271 : BUF_X1 port map( A => n461, Z => n474);
   U272 : AND2_X1 port map( A1 => n1750, A2 => n1759, ZN => n1171);
   U273 : AND2_X1 port map( A1 => n1750, A2 => n1758, ZN => n1172);
   U274 : AND2_X1 port map( A1 => n1755, A2 => n1759, ZN => n1176);
   U275 : AND2_X1 port map( A1 => n1755, A2 => n1758, ZN => n1177);
   U276 : AND2_X1 port map( A1 => n1751, A2 => n1750, ZN => n1161);
   U277 : AND2_X1 port map( A1 => n1749, A2 => n1750, ZN => n1162);
   U278 : AND2_X1 port map( A1 => n1768, A2 => n1750, ZN => n1185);
   U279 : AND2_X1 port map( A1 => n1767, A2 => n1750, ZN => n1186);
   U280 : AND2_X1 port map( A1 => n1773, A2 => n1750, ZN => n1195);
   U281 : AND2_X1 port map( A1 => n1772, A2 => n1750, ZN => n1196);
   U282 : AND2_X1 port map( A1 => n1751, A2 => n1754, ZN => n1166);
   U283 : AND2_X1 port map( A1 => n1768, A2 => n1754, ZN => n1190);
   U284 : AND2_X1 port map( A1 => n1773, A2 => n1754, ZN => n1200);
   U285 : NAND2_X1 port map( A1 => n472, A2 => n1151, ZN => N409);
   U286 : NAND2_X1 port map( A1 => RD2, A2 => ENABLE, ZN => n1151);
   U287 : NAND2_X1 port map( A1 => n473, A2 => n1776, ZN => N376);
   U288 : NAND2_X1 port map( A1 => RD1, A2 => ENABLE, ZN => n1776);
   U289 : NOR2_X1 port map( A1 => n2252, A2 => ADD_RD2(2), ZN => n1125);
   U290 : INV_X1 port map( A => ADD_RD2(0), ZN => n2251);
   U291 : BUF_X1 port map( A => n1790, Z => n2);
   U292 : BUF_X1 port map( A => n1790, Z => n1);
   U293 : INV_X1 port map( A => ADD_RD2(1), ZN => n2252);
   U294 : INV_X1 port map( A => ADD_RD2(2), ZN => n2253);
   U295 : BUF_X1 port map( A => n1790, Z => n3);
   U296 : NOR2_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), ZN => n1145);
   U297 : NOR2_X1 port map( A1 => n2254, A2 => ADD_RD2(4), ZN => n1150);
   U298 : INV_X1 port map( A => ADD_RD1(0), ZN => n2255);
   U299 : AND2_X1 port map( A1 => ADD_RD2(0), A2 => n1136, ZN => n1134);
   U300 : INV_X1 port map( A => ADD_RD2(3), ZN => n2254);
   U301 : AND2_X1 port map( A1 => ADD_RD1(0), A2 => n1761, ZN => n1759);
   U302 : AND2_X1 port map( A1 => n1131, A2 => ADD_RD2(0), ZN => n1126);
   U303 : AND2_X1 port map( A1 => n1145, A2 => ADD_RD2(0), ZN => n1143);
   U304 : AND2_X1 port map( A1 => n1150, A2 => ADD_RD2(0), ZN => n1148);
   U305 : AND2_X1 port map( A1 => n1756, A2 => ADD_RD1(0), ZN => n1751);
   U306 : AND2_X1 port map( A1 => n1770, A2 => ADD_RD1(0), ZN => n1768);
   U307 : AND2_X1 port map( A1 => n1775, A2 => ADD_RD1(0), ZN => n1773);
   U308 : NOR2_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), ZN => n1770);
   U309 : NOR2_X1 port map( A1 => n2258, A2 => ADD_RD1(4), ZN => n1775);
   U310 : INV_X1 port map( A => ADD_RD1(1), ZN => n2256);
   U311 : BUF_X1 port map( A => N313, Z => n454);
   U312 : BUF_X1 port map( A => N314, Z => n450);
   U313 : BUF_X1 port map( A => N315, Z => n446);
   U314 : BUF_X1 port map( A => N316, Z => n442);
   U315 : BUF_X1 port map( A => N317, Z => n438_port);
   U316 : BUF_X1 port map( A => N318, Z => n434_port);
   U317 : BUF_X1 port map( A => N319, Z => n430_port);
   U318 : BUF_X1 port map( A => N320, Z => n426_port);
   U319 : BUF_X1 port map( A => N321, Z => n422_port);
   U320 : BUF_X1 port map( A => N322, Z => n418_port);
   U321 : BUF_X1 port map( A => N323, Z => n414_port);
   U322 : BUF_X1 port map( A => N324, Z => n410_port);
   U323 : BUF_X1 port map( A => N325, Z => n406_port);
   U324 : BUF_X1 port map( A => N326, Z => n402_port);
   U325 : BUF_X1 port map( A => N327, Z => n398_port);
   U326 : BUF_X1 port map( A => N328, Z => n394_port);
   U327 : BUF_X1 port map( A => N329, Z => n390_port);
   U328 : BUF_X1 port map( A => N330, Z => n386_port);
   U329 : BUF_X1 port map( A => N331, Z => n382_port);
   U330 : BUF_X1 port map( A => N332, Z => n378_port);
   U331 : BUF_X1 port map( A => N333, Z => n374_port);
   U332 : BUF_X1 port map( A => N334, Z => n370_port);
   U333 : BUF_X1 port map( A => N335, Z => n366_port);
   U334 : BUF_X1 port map( A => N336, Z => n362_port);
   U335 : BUF_X1 port map( A => N337, Z => n358_port);
   U336 : BUF_X1 port map( A => N338, Z => n354_port);
   U337 : BUF_X1 port map( A => N339, Z => n350_port);
   U338 : BUF_X1 port map( A => N340, Z => n346_port);
   U339 : BUF_X1 port map( A => N341, Z => n342_port);
   U340 : BUF_X1 port map( A => N342, Z => n338_port);
   U341 : BUF_X1 port map( A => N343, Z => n334_port);
   U342 : BUF_X1 port map( A => N344, Z => n330_port);
   U343 : BUF_X1 port map( A => N313, Z => n453);
   U344 : BUF_X1 port map( A => N314, Z => n449);
   U345 : BUF_X1 port map( A => N315, Z => n445);
   U346 : BUF_X1 port map( A => N316, Z => n441_port);
   U347 : BUF_X1 port map( A => N317, Z => n437_port);
   U348 : BUF_X1 port map( A => N318, Z => n433_port);
   U349 : BUF_X1 port map( A => N319, Z => n429_port);
   U350 : BUF_X1 port map( A => N320, Z => n425_port);
   U351 : BUF_X1 port map( A => N321, Z => n421_port);
   U352 : BUF_X1 port map( A => N322, Z => n417_port);
   U353 : BUF_X1 port map( A => N323, Z => n413_port);
   U354 : BUF_X1 port map( A => N324, Z => n409_port);
   U355 : BUF_X1 port map( A => N325, Z => n405_port);
   U356 : BUF_X1 port map( A => N326, Z => n401_port);
   U357 : BUF_X1 port map( A => N327, Z => n397_port);
   U358 : BUF_X1 port map( A => N328, Z => n393_port);
   U359 : BUF_X1 port map( A => N329, Z => n389_port);
   U360 : BUF_X1 port map( A => N330, Z => n385_port);
   U361 : BUF_X1 port map( A => N331, Z => n381_port);
   U362 : BUF_X1 port map( A => N332, Z => n377_port);
   U363 : BUF_X1 port map( A => N333, Z => n373_port);
   U364 : BUF_X1 port map( A => N334, Z => n369_port);
   U365 : BUF_X1 port map( A => N335, Z => n365_port);
   U366 : BUF_X1 port map( A => N336, Z => n361_port);
   U367 : BUF_X1 port map( A => N337, Z => n357_port);
   U368 : BUF_X1 port map( A => N338, Z => n353_port);
   U369 : BUF_X1 port map( A => N339, Z => n349_port);
   U370 : BUF_X1 port map( A => N340, Z => n345_port);
   U371 : BUF_X1 port map( A => N341, Z => n341_port);
   U372 : BUF_X1 port map( A => N342, Z => n337_port);
   U373 : BUF_X1 port map( A => N343, Z => n333_port);
   U374 : BUF_X1 port map( A => N344, Z => n329_port);
   U375 : BUF_X1 port map( A => N313, Z => n452);
   U376 : BUF_X1 port map( A => N314, Z => n448);
   U377 : BUF_X1 port map( A => N315, Z => n444);
   U378 : BUF_X1 port map( A => N316, Z => n440_port);
   U379 : BUF_X1 port map( A => N317, Z => n436_port);
   U380 : BUF_X1 port map( A => N318, Z => n432_port);
   U381 : BUF_X1 port map( A => N319, Z => n428_port);
   U382 : BUF_X1 port map( A => N320, Z => n424_port);
   U383 : BUF_X1 port map( A => N321, Z => n420_port);
   U384 : BUF_X1 port map( A => N322, Z => n416_port);
   U385 : BUF_X1 port map( A => N323, Z => n412_port);
   U386 : BUF_X1 port map( A => N324, Z => n408_port);
   U387 : BUF_X1 port map( A => N325, Z => n404_port);
   U388 : BUF_X1 port map( A => N326, Z => n400_port);
   U389 : BUF_X1 port map( A => N327, Z => n396_port);
   U390 : BUF_X1 port map( A => N328, Z => n392_port);
   U391 : BUF_X1 port map( A => N329, Z => n388_port);
   U392 : BUF_X1 port map( A => N330, Z => n384_port);
   U393 : BUF_X1 port map( A => N331, Z => n380_port);
   U394 : BUF_X1 port map( A => N332, Z => n376_port);
   U395 : BUF_X1 port map( A => N333, Z => n372_port);
   U396 : BUF_X1 port map( A => N334, Z => n368_port);
   U397 : BUF_X1 port map( A => N335, Z => n364_port);
   U398 : BUF_X1 port map( A => N336, Z => n360_port);
   U399 : BUF_X1 port map( A => N337, Z => n356_port);
   U400 : BUF_X1 port map( A => N338, Z => n352_port);
   U401 : BUF_X1 port map( A => N339, Z => n348_port);
   U402 : BUF_X1 port map( A => N340, Z => n344_port);
   U403 : BUF_X1 port map( A => N341, Z => n340_port);
   U404 : BUF_X1 port map( A => N342, Z => n336_port);
   U405 : BUF_X1 port map( A => N343, Z => n332_port);
   U406 : BUF_X1 port map( A => N344, Z => n328_port);
   U407 : INV_X1 port map( A => ADD_RD1(3), ZN => n2258);
   U408 : AND2_X1 port map( A1 => ADD_RD2(4), A2 => ADD_RD2(3), ZN => n1136);
   U409 : AND2_X1 port map( A1 => ADD_RD2(4), A2 => n2254, ZN => n1131);
   U410 : AND2_X1 port map( A1 => ADD_RD1(4), A2 => ADD_RD1(3), ZN => n1761);
   U411 : AND2_X1 port map( A1 => ADD_RD1(4), A2 => n2258, ZN => n1756);
   U412 : BUF_X1 port map( A => RESET, Z => n460);
   U413 : BUF_X1 port map( A => RESET, Z => n461);
   U414 : OAI21_X1 port map( B1 => n1778, B2 => n1785, A => n466, ZN => N368);
   U415 : OAI21_X1 port map( B1 => n1778, B2 => n1784, A => n466, ZN => N369);
   U416 : OAI21_X1 port map( B1 => n1778, B2 => n1783, A => n466, ZN => N370);
   U417 : OAI21_X1 port map( B1 => n1778, B2 => n1782, A => n465, ZN => N371);
   U418 : OAI21_X1 port map( B1 => n1778, B2 => n1781, A => n465, ZN => N372);
   U419 : OAI21_X1 port map( B1 => n1778, B2 => n1780, A => n465, ZN => N373);
   U420 : OAI21_X1 port map( B1 => n1778, B2 => n1779, A => n465, ZN => N374);
   U421 : OAI21_X1 port map( B1 => n1785, B2 => n1789, A => n472, ZN => N312);
   U422 : OAI21_X1 port map( B1 => n1784, B2 => n1789, A => n470, ZN => N345);
   U423 : OAI21_X1 port map( B1 => n1783, B2 => n1789, A => n472, ZN => N346);
   U424 : OAI21_X1 port map( B1 => n1782, B2 => n1789, A => n472, ZN => N347);
   U425 : OAI21_X1 port map( B1 => n1781, B2 => n1789, A => n471, ZN => N348);
   U426 : OAI21_X1 port map( B1 => n1780, B2 => n1789, A => n471, ZN => N349);
   U427 : OAI21_X1 port map( B1 => n1779, B2 => n1789, A => n471, ZN => N350);
   U428 : OAI21_X1 port map( B1 => n1786, B2 => n1789, A => n471, ZN => N351);
   U429 : OAI21_X1 port map( B1 => n1785, B2 => n1787, A => n468, ZN => N360);
   U430 : OAI21_X1 port map( B1 => n1784, B2 => n1787, A => n468, ZN => N361);
   U431 : OAI21_X1 port map( B1 => n1783, B2 => n1787, A => n468, ZN => N362);
   U432 : OAI21_X1 port map( B1 => n1782, B2 => n1787, A => n467, ZN => N363);
   U433 : OAI21_X1 port map( B1 => n1781, B2 => n1787, A => n467, ZN => N364);
   U434 : OAI21_X1 port map( B1 => n1780, B2 => n1787, A => n467, ZN => N365);
   U435 : OAI21_X1 port map( B1 => n1779, B2 => n1787, A => n467, ZN => N366);
   U436 : OAI21_X1 port map( B1 => n1786, B2 => n1787, A => n466, ZN => N367);
   U437 : OAI21_X1 port map( B1 => n1785, B2 => n1788, A => n470, ZN => N352);
   U438 : OAI21_X1 port map( B1 => n1784, B2 => n1788, A => n470, ZN => N353);
   U439 : OAI21_X1 port map( B1 => n1783, B2 => n1788, A => n470, ZN => N354);
   U440 : OAI21_X1 port map( B1 => n1782, B2 => n1788, A => n469, ZN => N355);
   U441 : OAI21_X1 port map( B1 => n1781, B2 => n1788, A => n469, ZN => N356);
   U442 : OAI21_X1 port map( B1 => n1780, B2 => n1788, A => n469, ZN => N357);
   U443 : OAI21_X1 port map( B1 => n1779, B2 => n1788, A => n469, ZN => N358);
   U444 : OAI21_X1 port map( B1 => n1786, B2 => n1788, A => n468, ZN => N359);
   U445 : AOI21_X1 port map( B1 => n1117, B2 => n1118, A => n464, ZN => N410);
   U446 : NOR4_X1 port map( A1 => n1137, A2 => n1138, A3 => n1139, A4 => n1140,
                           ZN => n1117);
   U447 : NOR4_X1 port map( A1 => n1119, A2 => n1120, A3 => n1121, A4 => n1122,
                           ZN => n1118);
   U448 : OAI221_X1 port map( B1 => n109, B2 => n1994, C1 => n106, C2 => n1962,
                           A => n1149, ZN => n1137);
   U449 : AOI21_X1 port map( B1 => n1742, B2 => n1743, A => n462, ZN => N377);
   U450 : NOR4_X1 port map( A1 => n1762, A2 => n1763, A3 => n1764, A4 => n1765,
                           ZN => n1742);
   U451 : NOR4_X1 port map( A1 => n1744, A2 => n1745, A3 => n1746, A4 => n1747,
                           ZN => n1743);
   U452 : OAI221_X1 port map( B1 => n1994, B2 => n13, C1 => n1962, C2 => n10, A
                           => n1774, ZN => n1762);
   U453 : AOI21_X1 port map( B1 => n1724, B2 => n1725, A => n462, ZN => N378);
   U454 : NOR4_X1 port map( A1 => n1734, A2 => n1735, A3 => n1736, A4 => n1737,
                           ZN => n1724);
   U455 : NOR4_X1 port map( A1 => n1726, A2 => n1727, A3 => n1728, A4 => n1729,
                           ZN => n1725);
   U456 : OAI221_X1 port map( B1 => n1993, B2 => n13, C1 => n1961, C2 => n10, A
                           => n1741, ZN => n1734);
   U457 : AOI21_X1 port map( B1 => n1706, B2 => n1707, A => n462, ZN => N379);
   U458 : NOR4_X1 port map( A1 => n1716, A2 => n1717, A3 => n1718, A4 => n1719,
                           ZN => n1706);
   U459 : NOR4_X1 port map( A1 => n1708, A2 => n1709, A3 => n1710, A4 => n1711,
                           ZN => n1707);
   U460 : OAI221_X1 port map( B1 => n1992, B2 => n13, C1 => n1960, C2 => n10, A
                           => n1723, ZN => n1716);
   U461 : AOI21_X1 port map( B1 => n1688, B2 => n1689, A => n462, ZN => N380);
   U462 : NOR4_X1 port map( A1 => n1698, A2 => n1699, A3 => n1700, A4 => n1701,
                           ZN => n1688);
   U463 : NOR4_X1 port map( A1 => n1690, A2 => n1691, A3 => n1692, A4 => n1693,
                           ZN => n1689);
   U464 : OAI221_X1 port map( B1 => n1991, B2 => n13, C1 => n1959, C2 => n10, A
                           => n1705, ZN => n1698);
   U465 : AOI21_X1 port map( B1 => n1670, B2 => n1671, A => n462, ZN => N381);
   U466 : NOR4_X1 port map( A1 => n1680, A2 => n1681, A3 => n1682, A4 => n1683,
                           ZN => n1670);
   U467 : NOR4_X1 port map( A1 => n1672, A2 => n1673, A3 => n1674, A4 => n1675,
                           ZN => n1671);
   U468 : OAI221_X1 port map( B1 => n1990, B2 => n13, C1 => n1958, C2 => n10, A
                           => n1687, ZN => n1680);
   U469 : AOI21_X1 port map( B1 => n1652, B2 => n1653, A => n462, ZN => N382);
   U470 : NOR4_X1 port map( A1 => n1662, A2 => n1663, A3 => n1664, A4 => n1665,
                           ZN => n1652);
   U471 : NOR4_X1 port map( A1 => n1654, A2 => n1655, A3 => n1656, A4 => n1657,
                           ZN => n1653);
   U472 : OAI221_X1 port map( B1 => n1989, B2 => n13, C1 => n1957, C2 => n10, A
                           => n1669, ZN => n1662);
   U473 : AOI21_X1 port map( B1 => n1634, B2 => n1635, A => n462, ZN => N383);
   U474 : NOR4_X1 port map( A1 => n1644, A2 => n1645, A3 => n1646, A4 => n1647,
                           ZN => n1634);
   U475 : NOR4_X1 port map( A1 => n1636, A2 => n1637, A3 => n1638, A4 => n1639,
                           ZN => n1635);
   U476 : OAI221_X1 port map( B1 => n1988, B2 => n13, C1 => n1956, C2 => n10, A
                           => n1651, ZN => n1644);
   U477 : AOI21_X1 port map( B1 => n1616, B2 => n1617, A => n462, ZN => N384);
   U478 : NOR4_X1 port map( A1 => n1626, A2 => n1627, A3 => n1628, A4 => n1629,
                           ZN => n1616);
   U479 : NOR4_X1 port map( A1 => n1618, A2 => n1619, A3 => n1620, A4 => n1621,
                           ZN => n1617);
   U480 : OAI221_X1 port map( B1 => n1987, B2 => n13, C1 => n1955, C2 => n10, A
                           => n1633, ZN => n1626);
   U481 : AOI21_X1 port map( B1 => n1598, B2 => n1599, A => n462, ZN => N385);
   U482 : NOR4_X1 port map( A1 => n1608, A2 => n1609, A3 => n1610, A4 => n1611,
                           ZN => n1598);
   U483 : NOR4_X1 port map( A1 => n1600, A2 => n1601, A3 => n1602, A4 => n1603,
                           ZN => n1599);
   U484 : OAI221_X1 port map( B1 => n1986, B2 => n13, C1 => n1954, C2 => n10, A
                           => n1615, ZN => n1608);
   U485 : AOI21_X1 port map( B1 => n1580, B2 => n1581, A => n462, ZN => N386);
   U486 : NOR4_X1 port map( A1 => n1590, A2 => n1591, A3 => n1592, A4 => n1593,
                           ZN => n1580);
   U487 : NOR4_X1 port map( A1 => n1582, A2 => n1583, A3 => n1584, A4 => n1585,
                           ZN => n1581);
   U488 : OAI221_X1 port map( B1 => n1985, B2 => n13, C1 => n1953, C2 => n10, A
                           => n1597, ZN => n1590);
   U489 : AOI21_X1 port map( B1 => n1562, B2 => n1563, A => n462, ZN => N387);
   U490 : NOR4_X1 port map( A1 => n1572, A2 => n1573, A3 => n1574, A4 => n1575,
                           ZN => n1562);
   U491 : NOR4_X1 port map( A1 => n1564, A2 => n1565, A3 => n1566, A4 => n1567,
                           ZN => n1563);
   U492 : OAI221_X1 port map( B1 => n1984, B2 => n13, C1 => n1952, C2 => n10, A
                           => n1579, ZN => n1572);
   U493 : AOI21_X1 port map( B1 => n1544, B2 => n1545, A => n463, ZN => N388);
   U494 : NOR4_X1 port map( A1 => n1554, A2 => n1555, A3 => n1556, A4 => n1557,
                           ZN => n1544);
   U495 : NOR4_X1 port map( A1 => n1546, A2 => n1547, A3 => n1548, A4 => n1549,
                           ZN => n1545);
   U496 : OAI221_X1 port map( B1 => n1983, B2 => n14, C1 => n1951, C2 => n11, A
                           => n1561, ZN => n1554);
   U497 : AOI21_X1 port map( B1 => n1526, B2 => n1527, A => n463, ZN => N389);
   U498 : NOR4_X1 port map( A1 => n1536, A2 => n1537, A3 => n1538, A4 => n1539,
                           ZN => n1526);
   U499 : NOR4_X1 port map( A1 => n1528, A2 => n1529, A3 => n1530, A4 => n1531,
                           ZN => n1527);
   U500 : OAI221_X1 port map( B1 => n1982, B2 => n14, C1 => n1950, C2 => n11, A
                           => n1543, ZN => n1536);
   U501 : AOI21_X1 port map( B1 => n1508, B2 => n1509, A => n463, ZN => N390);
   U502 : NOR4_X1 port map( A1 => n1518, A2 => n1519, A3 => n1520, A4 => n1521,
                           ZN => n1508);
   U503 : NOR4_X1 port map( A1 => n1510, A2 => n1511, A3 => n1512, A4 => n1513,
                           ZN => n1509);
   U504 : OAI221_X1 port map( B1 => n1981, B2 => n14, C1 => n1949, C2 => n11, A
                           => n1525, ZN => n1518);
   U505 : AOI21_X1 port map( B1 => n1490, B2 => n1491, A => n463, ZN => N391);
   U506 : NOR4_X1 port map( A1 => n1500, A2 => n1501, A3 => n1502, A4 => n1503,
                           ZN => n1490);
   U507 : NOR4_X1 port map( A1 => n1492, A2 => n1493, A3 => n1494, A4 => n1495,
                           ZN => n1491);
   U508 : OAI221_X1 port map( B1 => n1980, B2 => n14, C1 => n1948, C2 => n11, A
                           => n1507, ZN => n1500);
   U509 : AOI21_X1 port map( B1 => n1472, B2 => n1473, A => n463, ZN => N392);
   U510 : NOR4_X1 port map( A1 => n1482, A2 => n1483, A3 => n1484, A4 => n1485,
                           ZN => n1472);
   U511 : NOR4_X1 port map( A1 => n1474, A2 => n1475, A3 => n1476, A4 => n1477,
                           ZN => n1473);
   U512 : OAI221_X1 port map( B1 => n1979, B2 => n14, C1 => n1947, C2 => n11, A
                           => n1489, ZN => n1482);
   U513 : AOI21_X1 port map( B1 => n1454, B2 => n1455, A => n463, ZN => N393);
   U514 : NOR4_X1 port map( A1 => n1464, A2 => n1465, A3 => n1466, A4 => n1467,
                           ZN => n1454);
   U515 : NOR4_X1 port map( A1 => n1456, A2 => n1457, A3 => n1458, A4 => n1459,
                           ZN => n1455);
   U516 : OAI221_X1 port map( B1 => n1978, B2 => n14, C1 => n1946, C2 => n11, A
                           => n1471, ZN => n1464);
   U517 : AOI21_X1 port map( B1 => n1436, B2 => n1437, A => n463, ZN => N394);
   U518 : NOR4_X1 port map( A1 => n1446, A2 => n1447, A3 => n1448, A4 => n1449,
                           ZN => n1436);
   U519 : NOR4_X1 port map( A1 => n1438, A2 => n1439, A3 => n1440, A4 => n1441,
                           ZN => n1437);
   U520 : OAI221_X1 port map( B1 => n1977, B2 => n14, C1 => n1945, C2 => n11, A
                           => n1453, ZN => n1446);
   U521 : AOI21_X1 port map( B1 => n1418, B2 => n1419, A => n463, ZN => N395);
   U522 : NOR4_X1 port map( A1 => n1428, A2 => n1429, A3 => n1430, A4 => n1431,
                           ZN => n1418);
   U523 : NOR4_X1 port map( A1 => n1420, A2 => n1421, A3 => n1422, A4 => n1423,
                           ZN => n1419);
   U524 : OAI221_X1 port map( B1 => n1976, B2 => n14, C1 => n1944, C2 => n11, A
                           => n1435, ZN => n1428);
   U525 : AOI21_X1 port map( B1 => n1400, B2 => n1401, A => n463, ZN => N396);
   U526 : NOR4_X1 port map( A1 => n1410, A2 => n1411, A3 => n1412, A4 => n1413,
                           ZN => n1400);
   U527 : NOR4_X1 port map( A1 => n1402, A2 => n1403, A3 => n1404, A4 => n1405,
                           ZN => n1401);
   U528 : OAI221_X1 port map( B1 => n1975, B2 => n14, C1 => n1943, C2 => n11, A
                           => n1417, ZN => n1410);
   U529 : AOI21_X1 port map( B1 => n1382, B2 => n1383, A => n463, ZN => N397);
   U530 : NOR4_X1 port map( A1 => n1392, A2 => n1393, A3 => n1394, A4 => n1395,
                           ZN => n1382);
   U531 : NOR4_X1 port map( A1 => n1384, A2 => n1385, A3 => n1386, A4 => n1387,
                           ZN => n1383);
   U532 : OAI221_X1 port map( B1 => n1974, B2 => n14, C1 => n1942, C2 => n11, A
                           => n1399, ZN => n1392);
   U533 : AOI21_X1 port map( B1 => n1364, B2 => n1365, A => n463, ZN => N398);
   U534 : NOR4_X1 port map( A1 => n1374, A2 => n1375, A3 => n1376, A4 => n1377,
                           ZN => n1364);
   U535 : NOR4_X1 port map( A1 => n1366, A2 => n1367, A3 => n1368, A4 => n1369,
                           ZN => n1365);
   U536 : OAI221_X1 port map( B1 => n1973, B2 => n14, C1 => n1941, C2 => n11, A
                           => n1381, ZN => n1374);
   U537 : AOI21_X1 port map( B1 => n1346, B2 => n1347, A => n464, ZN => N399);
   U538 : NOR4_X1 port map( A1 => n1356, A2 => n1357, A3 => n1358, A4 => n1359,
                           ZN => n1346);
   U539 : NOR4_X1 port map( A1 => n1348, A2 => n1349, A3 => n1350, A4 => n1351,
                           ZN => n1347);
   U540 : OAI221_X1 port map( B1 => n1972, B2 => n15, C1 => n1940, C2 => n12, A
                           => n1363, ZN => n1356);
   U541 : AOI21_X1 port map( B1 => n1328, B2 => n1329, A => n464, ZN => N400);
   U542 : NOR4_X1 port map( A1 => n1338, A2 => n1339, A3 => n1340, A4 => n1341,
                           ZN => n1328);
   U543 : NOR4_X1 port map( A1 => n1330, A2 => n1331, A3 => n1332, A4 => n1333,
                           ZN => n1329);
   U544 : OAI221_X1 port map( B1 => n1971, B2 => n15, C1 => n1939, C2 => n12, A
                           => n1345, ZN => n1338);
   U545 : AOI21_X1 port map( B1 => n1310, B2 => n1311, A => n464, ZN => N401);
   U546 : NOR4_X1 port map( A1 => n1320, A2 => n1321, A3 => n1322, A4 => n1323,
                           ZN => n1310);
   U547 : NOR4_X1 port map( A1 => n1312, A2 => n1313, A3 => n1314, A4 => n1315,
                           ZN => n1311);
   U548 : OAI221_X1 port map( B1 => n1970, B2 => n15, C1 => n1938, C2 => n12, A
                           => n1327, ZN => n1320);
   U549 : AOI21_X1 port map( B1 => n1292, B2 => n1293, A => n464, ZN => N402);
   U550 : NOR4_X1 port map( A1 => n1302, A2 => n1303, A3 => n1304, A4 => n1305,
                           ZN => n1292);
   U551 : NOR4_X1 port map( A1 => n1294, A2 => n1295, A3 => n1296, A4 => n1297,
                           ZN => n1293);
   U552 : OAI221_X1 port map( B1 => n1969, B2 => n15, C1 => n1937, C2 => n12, A
                           => n1309, ZN => n1302);
   U553 : AOI21_X1 port map( B1 => n1274, B2 => n1275, A => n464, ZN => N403);
   U554 : NOR4_X1 port map( A1 => n1284, A2 => n1285, A3 => n1286, A4 => n1287,
                           ZN => n1274);
   U555 : NOR4_X1 port map( A1 => n1276, A2 => n1277, A3 => n1278, A4 => n1279,
                           ZN => n1275);
   U556 : OAI221_X1 port map( B1 => n1968, B2 => n15, C1 => n1936, C2 => n12, A
                           => n1291, ZN => n1284);
   U557 : AOI21_X1 port map( B1 => n1256, B2 => n1257, A => n464, ZN => N404);
   U558 : NOR4_X1 port map( A1 => n1266, A2 => n1267, A3 => n1268, A4 => n1269,
                           ZN => n1256);
   U559 : NOR4_X1 port map( A1 => n1258, A2 => n1259, A3 => n1260, A4 => n1261,
                           ZN => n1257);
   U560 : OAI221_X1 port map( B1 => n1967, B2 => n15, C1 => n1935, C2 => n12, A
                           => n1273, ZN => n1266);
   U561 : AOI21_X1 port map( B1 => n1238, B2 => n1239, A => n464, ZN => N405);
   U562 : NOR4_X1 port map( A1 => n1248, A2 => n1249, A3 => n1250, A4 => n1251,
                           ZN => n1238);
   U563 : NOR4_X1 port map( A1 => n1240, A2 => n1241, A3 => n1242, A4 => n1243,
                           ZN => n1239);
   U564 : OAI221_X1 port map( B1 => n1966, B2 => n15, C1 => n1934, C2 => n12, A
                           => n1255, ZN => n1248);
   U565 : AOI21_X1 port map( B1 => n1220, B2 => n1221, A => n464, ZN => N406);
   U566 : NOR4_X1 port map( A1 => n1230, A2 => n1231, A3 => n1232, A4 => n1233,
                           ZN => n1220);
   U567 : NOR4_X1 port map( A1 => n1222, A2 => n1223, A3 => n1224, A4 => n1225,
                           ZN => n1221);
   U568 : OAI221_X1 port map( B1 => n1965, B2 => n15, C1 => n1933, C2 => n12, A
                           => n1237, ZN => n1230);
   U569 : AOI21_X1 port map( B1 => n1202, B2 => n1203, A => n464, ZN => N407);
   U570 : NOR4_X1 port map( A1 => n1212, A2 => n1213, A3 => n1214, A4 => n1215,
                           ZN => n1202);
   U571 : NOR4_X1 port map( A1 => n1204, A2 => n1205, A3 => n1206, A4 => n1207,
                           ZN => n1203);
   U572 : OAI221_X1 port map( B1 => n1964, B2 => n15, C1 => n1932, C2 => n12, A
                           => n1219, ZN => n1212);
   U573 : AOI21_X1 port map( B1 => n1152, B2 => n1153, A => n464, ZN => N408);
   U574 : NOR4_X1 port map( A1 => n1178, A2 => n1179, A3 => n1180, A4 => n1181,
                           ZN => n1152);
   U575 : NOR4_X1 port map( A1 => n1154, A2 => n1155, A3 => n1156, A4 => n1157,
                           ZN => n1153);
   U576 : OAI221_X1 port map( B1 => n1963, B2 => n15, C1 => n1931, C2 => n12, A
                           => n1199, ZN => n1178);
   U577 : AOI21_X1 port map( B1 => n1099, B2 => n1100, A => n464, ZN => N411);
   U578 : NOR4_X1 port map( A1 => n1109, A2 => n1110, A3 => n1111, A4 => n1112,
                           ZN => n1099);
   U579 : NOR4_X1 port map( A1 => n1101, A2 => n1102, A3 => n1103, A4 => n1104,
                           ZN => n1100);
   U580 : OAI221_X1 port map( B1 => n109, B2 => n1993, C1 => n106, C2 => n1961,
                           A => n1116, ZN => n1109);
   U581 : AOI21_X1 port map( B1 => n1081, B2 => n1082, A => n462, ZN => N412);
   U582 : NOR4_X1 port map( A1 => n1091, A2 => n1092, A3 => n1093, A4 => n1094,
                           ZN => n1081);
   U583 : NOR4_X1 port map( A1 => n1083, A2 => n1084, A3 => n1085, A4 => n1086,
                           ZN => n1082);
   U584 : OAI221_X1 port map( B1 => n109, B2 => n1992, C1 => n106, C2 => n1960,
                           A => n1098, ZN => n1091);
   U585 : AOI21_X1 port map( B1 => n1063, B2 => n1064, A => n463, ZN => N413);
   U586 : NOR4_X1 port map( A1 => n1073, A2 => n1074, A3 => n1075, A4 => n1076,
                           ZN => n1063);
   U587 : NOR4_X1 port map( A1 => n1065, A2 => n1066, A3 => n1067, A4 => n1068,
                           ZN => n1064);
   U588 : OAI221_X1 port map( B1 => n109, B2 => n1991, C1 => n106, C2 => n1959,
                           A => n1080, ZN => n1073);
   U589 : AOI21_X1 port map( B1 => n1045, B2 => n1046, A => n464, ZN => N414);
   U590 : NOR4_X1 port map( A1 => n1055, A2 => n1056, A3 => n1057, A4 => n1058,
                           ZN => n1045);
   U591 : NOR4_X1 port map( A1 => n1047, A2 => n1048, A3 => n1049, A4 => n1050,
                           ZN => n1046);
   U592 : OAI221_X1 port map( B1 => n109, B2 => n1990, C1 => n106, C2 => n1958,
                           A => n1062, ZN => n1055);
   U593 : AOI21_X1 port map( B1 => n1027, B2 => n1028, A => n462, ZN => N415);
   U594 : NOR4_X1 port map( A1 => n1037, A2 => n1038, A3 => n1039, A4 => n1040,
                           ZN => n1027);
   U595 : NOR4_X1 port map( A1 => n1029, A2 => n1030, A3 => n1031, A4 => n1032,
                           ZN => n1028);
   U596 : OAI221_X1 port map( B1 => n109, B2 => n1989, C1 => n106, C2 => n1957,
                           A => n1044, ZN => n1037);
   U597 : AOI21_X1 port map( B1 => n1009, B2 => n1010, A => n463, ZN => N416);
   U598 : NOR4_X1 port map( A1 => n1019, A2 => n1020, A3 => n1021, A4 => n1022,
                           ZN => n1009);
   U599 : NOR4_X1 port map( A1 => n1011, A2 => n1012, A3 => n1013, A4 => n1014,
                           ZN => n1010);
   U600 : OAI221_X1 port map( B1 => n109, B2 => n1988, C1 => n106, C2 => n1956,
                           A => n1026, ZN => n1019);
   U601 : AOI21_X1 port map( B1 => n991, B2 => n992, A => n464, ZN => N417);
   U602 : NOR4_X1 port map( A1 => n1001, A2 => n1002, A3 => n1003, A4 => n1004,
                           ZN => n991);
   U603 : NOR4_X1 port map( A1 => n993, A2 => n994, A3 => n995, A4 => n996, ZN 
                           => n992);
   U604 : OAI221_X1 port map( B1 => n109, B2 => n1987, C1 => n106, C2 => n1955,
                           A => n1008, ZN => n1001);
   U605 : AOI21_X1 port map( B1 => n973, B2 => n974, A => n462, ZN => N418);
   U606 : NOR4_X1 port map( A1 => n983, A2 => n984, A3 => n985, A4 => n986, ZN 
                           => n973);
   U607 : NOR4_X1 port map( A1 => n975, A2 => n976, A3 => n977, A4 => n978, ZN 
                           => n974);
   U608 : OAI221_X1 port map( B1 => n109, B2 => n1986, C1 => n106, C2 => n1954,
                           A => n990, ZN => n983);
   U609 : AOI21_X1 port map( B1 => n955, B2 => n956, A => n463, ZN => N419);
   U610 : NOR4_X1 port map( A1 => n965, A2 => n966, A3 => n967, A4 => n968, ZN 
                           => n955);
   U611 : NOR4_X1 port map( A1 => n957, A2 => n958, A3 => n959, A4 => n960, ZN 
                           => n956);
   U612 : OAI221_X1 port map( B1 => n109, B2 => n1985, C1 => n106, C2 => n1953,
                           A => n972, ZN => n965);
   U613 : AOI21_X1 port map( B1 => n937, B2 => n938, A => n464, ZN => N420);
   U614 : NOR4_X1 port map( A1 => n947, A2 => n948, A3 => n949, A4 => n950, ZN 
                           => n937);
   U615 : NOR4_X1 port map( A1 => n939, A2 => n940, A3 => n941, A4 => n942, ZN 
                           => n938);
   U616 : OAI221_X1 port map( B1 => n109, B2 => n1984, C1 => n106, C2 => n1952,
                           A => n954, ZN => n947);
   U617 : AOI21_X1 port map( B1 => n919, B2 => n920, A => n462, ZN => N421);
   U618 : NOR4_X1 port map( A1 => n929, A2 => n930, A3 => n931, A4 => n932, ZN 
                           => n919);
   U619 : NOR4_X1 port map( A1 => n921, A2 => n922, A3 => n923, A4 => n924, ZN 
                           => n920);
   U620 : OAI221_X1 port map( B1 => n109, B2 => n1983, C1 => n107, C2 => n1951,
                           A => n936, ZN => n929);
   U621 : AOI21_X1 port map( B1 => n901, B2 => n902, A => n463, ZN => N422);
   U622 : NOR4_X1 port map( A1 => n911, A2 => n912, A3 => n913, A4 => n914, ZN 
                           => n901);
   U623 : NOR4_X1 port map( A1 => n903, A2 => n904, A3 => n905, A4 => n906, ZN 
                           => n902);
   U624 : OAI221_X1 port map( B1 => n110, B2 => n1982, C1 => n107, C2 => n1950,
                           A => n918, ZN => n911);
   U625 : AOI21_X1 port map( B1 => n883, B2 => n884, A => n464, ZN => N423);
   U626 : NOR4_X1 port map( A1 => n893, A2 => n894, A3 => n895, A4 => n896, ZN 
                           => n883);
   U627 : NOR4_X1 port map( A1 => n885, A2 => n886, A3 => n887, A4 => n888, ZN 
                           => n884);
   U628 : OAI221_X1 port map( B1 => n110, B2 => n1981, C1 => n107, C2 => n1949,
                           A => n900, ZN => n893);
   U629 : AOI21_X1 port map( B1 => n865, B2 => n866, A => n462, ZN => N424);
   U630 : NOR4_X1 port map( A1 => n875, A2 => n876, A3 => n877, A4 => n878, ZN 
                           => n865);
   U631 : NOR4_X1 port map( A1 => n867, A2 => n868, A3 => n869, A4 => n870, ZN 
                           => n866);
   U632 : OAI221_X1 port map( B1 => n110, B2 => n1980, C1 => n107, C2 => n1948,
                           A => n882, ZN => n875);
   U633 : AOI21_X1 port map( B1 => n847, B2 => n848, A => n462, ZN => N425);
   U634 : NOR4_X1 port map( A1 => n857, A2 => n858, A3 => n859, A4 => n860, ZN 
                           => n847);
   U635 : NOR4_X1 port map( A1 => n849, A2 => n850, A3 => n851, A4 => n852, ZN 
                           => n848);
   U636 : OAI221_X1 port map( B1 => n110, B2 => n1979, C1 => n107, C2 => n1947,
                           A => n864, ZN => n857);
   U637 : AOI21_X1 port map( B1 => n829, B2 => n830, A => n463, ZN => N426);
   U638 : NOR4_X1 port map( A1 => n839, A2 => n840, A3 => n841, A4 => n842, ZN 
                           => n829);
   U639 : NOR4_X1 port map( A1 => n831, A2 => n832, A3 => n833, A4 => n834, ZN 
                           => n830);
   U640 : OAI221_X1 port map( B1 => n110, B2 => n1978, C1 => n107, C2 => n1946,
                           A => n846, ZN => n839);
   U641 : AOI21_X1 port map( B1 => n811, B2 => n812, A => n464, ZN => N427);
   U642 : NOR4_X1 port map( A1 => n821, A2 => n822, A3 => n823, A4 => n824, ZN 
                           => n811);
   U643 : NOR4_X1 port map( A1 => n813, A2 => n814, A3 => n815, A4 => n816, ZN 
                           => n812);
   U644 : OAI221_X1 port map( B1 => n110, B2 => n1977, C1 => n107, C2 => n1945,
                           A => n828, ZN => n821);
   U645 : AOI21_X1 port map( B1 => n793, B2 => n794, A => n463, ZN => N428);
   U646 : NOR4_X1 port map( A1 => n803, A2 => n804, A3 => n805, A4 => n806, ZN 
                           => n793);
   U647 : NOR4_X1 port map( A1 => n795, A2 => n796, A3 => n797, A4 => n798, ZN 
                           => n794);
   U648 : OAI221_X1 port map( B1 => n110, B2 => n1976, C1 => n107, C2 => n1944,
                           A => n810, ZN => n803);
   U649 : AOI21_X1 port map( B1 => n775, B2 => n776, A => n462, ZN => N429);
   U650 : NOR4_X1 port map( A1 => n785, A2 => n786, A3 => n787, A4 => n788, ZN 
                           => n775);
   U651 : NOR4_X1 port map( A1 => n777, A2 => n778, A3 => n779, A4 => n780, ZN 
                           => n776);
   U652 : OAI221_X1 port map( B1 => n110, B2 => n1975, C1 => n107, C2 => n1943,
                           A => n792, ZN => n785);
   U653 : AOI21_X1 port map( B1 => n757, B2 => n758, A => n463, ZN => N430);
   U654 : NOR4_X1 port map( A1 => n767, A2 => n768, A3 => n769, A4 => n770, ZN 
                           => n757);
   U655 : NOR4_X1 port map( A1 => n759, A2 => n760, A3 => n761, A4 => n762, ZN 
                           => n758);
   U656 : OAI221_X1 port map( B1 => n110, B2 => n1974, C1 => n107, C2 => n1942,
                           A => n774, ZN => n767);
   U657 : AOI21_X1 port map( B1 => n739, B2 => n740, A => n464, ZN => N431);
   U658 : NOR4_X1 port map( A1 => n749, A2 => n750, A3 => n751, A4 => n752, ZN 
                           => n739);
   U659 : NOR4_X1 port map( A1 => n741, A2 => n742, A3 => n743, A4 => n744, ZN 
                           => n740);
   U660 : OAI221_X1 port map( B1 => n110, B2 => n1973, C1 => n107, C2 => n1941,
                           A => n756, ZN => n749);
   U661 : AOI21_X1 port map( B1 => n721, B2 => n722, A => n464, ZN => N432);
   U662 : NOR4_X1 port map( A1 => n731, A2 => n732, A3 => n733, A4 => n734, ZN 
                           => n721);
   U663 : NOR4_X1 port map( A1 => n723, A2 => n724, A3 => n725, A4 => n726, ZN 
                           => n722);
   U664 : OAI221_X1 port map( B1 => n110, B2 => n1972, C1 => n108, C2 => n1940,
                           A => n738, ZN => n731);
   U665 : AOI21_X1 port map( B1 => n703, B2 => n704, A => n462, ZN => N433);
   U666 : NOR4_X1 port map( A1 => n713, A2 => n714, A3 => n715, A4 => n716, ZN 
                           => n703);
   U667 : NOR4_X1 port map( A1 => n705, A2 => n706, A3 => n707, A4 => n708, ZN 
                           => n704);
   U668 : OAI221_X1 port map( B1 => n110, B2 => n1971, C1 => n108, C2 => n1939,
                           A => n720, ZN => n713);
   U669 : AOI21_X1 port map( B1 => n685, B2 => n686, A => n463, ZN => N434);
   U670 : NOR4_X1 port map( A1 => n695, A2 => n696, A3 => n697, A4 => n698, ZN 
                           => n685);
   U671 : NOR4_X1 port map( A1 => n687, A2 => n688, A3 => n689, A4 => n690, ZN 
                           => n686);
   U672 : OAI221_X1 port map( B1 => n111, B2 => n1970, C1 => n108, C2 => n1938,
                           A => n702, ZN => n695);
   U673 : AOI21_X1 port map( B1 => n667, B2 => n668, A => n464, ZN => N435);
   U674 : NOR4_X1 port map( A1 => n677, A2 => n678, A3 => n679, A4 => n680, ZN 
                           => n667);
   U675 : NOR4_X1 port map( A1 => n669, A2 => n670, A3 => n671, A4 => n672, ZN 
                           => n668);
   U676 : OAI221_X1 port map( B1 => n111, B2 => n1969, C1 => n108, C2 => n1937,
                           A => n684, ZN => n677);
   U677 : AOI21_X1 port map( B1 => n649, B2 => n650, A => n462, ZN => N436);
   U678 : NOR4_X1 port map( A1 => n659, A2 => n660, A3 => n661, A4 => n662, ZN 
                           => n649);
   U679 : NOR4_X1 port map( A1 => n651, A2 => n652, A3 => n653, A4 => n654, ZN 
                           => n650);
   U680 : OAI221_X1 port map( B1 => n111, B2 => n1968, C1 => n108, C2 => n1936,
                           A => n666, ZN => n659);
   U681 : AOI21_X1 port map( B1 => n631, B2 => n632, A => n462, ZN => N437);
   U682 : NOR4_X1 port map( A1 => n641, A2 => n642, A3 => n643, A4 => n644, ZN 
                           => n631);
   U683 : NOR4_X1 port map( A1 => n633, A2 => n634, A3 => n635, A4 => n636, ZN 
                           => n632);
   U684 : OAI221_X1 port map( B1 => n111, B2 => n1967, C1 => n108, C2 => n1935,
                           A => n648, ZN => n641);
   U685 : AOI21_X1 port map( B1 => n613, B2 => n614, A => n462, ZN => N438);
   U686 : NOR4_X1 port map( A1 => n623, A2 => n624, A3 => n625, A4 => n626, ZN 
                           => n613);
   U687 : NOR4_X1 port map( A1 => n615, A2 => n616, A3 => n617, A4 => n618, ZN 
                           => n614);
   U688 : OAI221_X1 port map( B1 => n111, B2 => n1966, C1 => n108, C2 => n1934,
                           A => n630, ZN => n623);
   U689 : AOI21_X1 port map( B1 => n595, B2 => n596, A => n463, ZN => N439);
   U690 : NOR4_X1 port map( A1 => n605, A2 => n606, A3 => n607, A4 => n608, ZN 
                           => n595);
   U691 : NOR4_X1 port map( A1 => n597, A2 => n598, A3 => n599, A4 => n600, ZN 
                           => n596);
   U692 : OAI221_X1 port map( B1 => n111, B2 => n1965, C1 => n108, C2 => n1933,
                           A => n612, ZN => n605);
   U693 : AOI21_X1 port map( B1 => n577, B2 => n578, A => n464, ZN => N440);
   U694 : NOR4_X1 port map( A1 => n587, A2 => n588, A3 => n589, A4 => n590, ZN 
                           => n577);
   U695 : NOR4_X1 port map( A1 => n579, A2 => n580, A3 => n581, A4 => n582, ZN 
                           => n578);
   U696 : OAI221_X1 port map( B1 => n111, B2 => n1964, C1 => n108, C2 => n1932,
                           A => n594, ZN => n587);
   U697 : AOI21_X1 port map( B1 => n527, B2 => n528, A => n463, ZN => N441);
   U698 : NOR4_X1 port map( A1 => n553, A2 => n554, A3 => n555, A4 => n556, ZN 
                           => n527);
   U699 : NOR4_X1 port map( A1 => n529, A2 => n530, A3 => n531, A4 => n532, ZN 
                           => n528);
   U700 : OAI221_X1 port map( B1 => n111, B2 => n1963, C1 => n108, C2 => n1931,
                           A => n574, ZN => n553);
   U701 : AND2_X1 port map( A1 => DATAIN(10), A2 => n2, ZN => N323);
   U702 : AND2_X1 port map( A1 => DATAIN(11), A2 => n2, ZN => N324);
   U703 : AND2_X1 port map( A1 => DATAIN(12), A2 => n2, ZN => N325);
   U704 : AND2_X1 port map( A1 => DATAIN(13), A2 => n2, ZN => N326);
   U705 : AND2_X1 port map( A1 => DATAIN(14), A2 => n2, ZN => N327);
   U706 : AND2_X1 port map( A1 => DATAIN(15), A2 => n2, ZN => N328);
   U707 : AND2_X1 port map( A1 => DATAIN(16), A2 => n2, ZN => N329);
   U708 : AND2_X1 port map( A1 => DATAIN(17), A2 => n2, ZN => N330);
   U709 : AND2_X1 port map( A1 => DATAIN(18), A2 => n2, ZN => N331);
   U710 : AND2_X1 port map( A1 => DATAIN(19), A2 => n2, ZN => N332);
   U711 : AND2_X1 port map( A1 => DATAIN(20), A2 => n2, ZN => N333);
   U712 : AND2_X1 port map( A1 => DATAIN(21), A2 => n1, ZN => N334);
   U713 : AND2_X1 port map( A1 => DATAIN(22), A2 => n1, ZN => N335);
   U714 : AND2_X1 port map( A1 => DATAIN(23), A2 => n1, ZN => N336);
   U715 : AND2_X1 port map( A1 => DATAIN(24), A2 => n1, ZN => N337);
   U716 : AND2_X1 port map( A1 => DATAIN(25), A2 => n1, ZN => N338);
   U717 : AND2_X1 port map( A1 => DATAIN(26), A2 => n1, ZN => N339);
   U718 : AND2_X1 port map( A1 => DATAIN(27), A2 => n1, ZN => N340);
   U719 : AND2_X1 port map( A1 => DATAIN(28), A2 => n1, ZN => N341);
   U720 : AND2_X1 port map( A1 => DATAIN(29), A2 => n1, ZN => N342);
   U721 : AND2_X1 port map( A1 => DATAIN(30), A2 => n1, ZN => N343);
   U722 : AND2_X1 port map( A1 => DATAIN(31), A2 => n1, ZN => N344);
   U723 : AND2_X1 port map( A1 => DATAIN(0), A2 => n3, ZN => N313);
   U724 : AND2_X1 port map( A1 => DATAIN(1), A2 => n3, ZN => N314);
   U725 : AND2_X1 port map( A1 => DATAIN(2), A2 => n3, ZN => N315);
   U726 : AND2_X1 port map( A1 => DATAIN(3), A2 => n3, ZN => N316);
   U727 : AND2_X1 port map( A1 => DATAIN(4), A2 => n3, ZN => N317);
   U728 : AND2_X1 port map( A1 => DATAIN(5), A2 => n3, ZN => N318);
   U729 : AND2_X1 port map( A1 => DATAIN(6), A2 => n3, ZN => N319);
   U730 : AND2_X1 port map( A1 => DATAIN(7), A2 => n3, ZN => N320);
   U731 : AND2_X1 port map( A1 => DATAIN(8), A2 => n3, ZN => N321);
   U732 : AND2_X1 port map( A1 => DATAIN(9), A2 => n3, ZN => N322);
   U733 : NAND2_X1 port map( A1 => n473, A2 => n1777, ZN => N375);
   U734 : AND2_X1 port map( A1 => n474, A2 => n1777, ZN => n1790);
   U735 : OAI221_X1 port map( B1 => n195, B2 => n2034, C1 => n192, C2 => n2002,
                           A => n691, ZN => n690);
   U736 : AOI22_X1 port map( A1 => REGISTERS_19_24_port, A2 => n189, B1 => 
                           REGISTERS_18_24_port, B2 => n186, ZN => n691);
   U737 : OAI221_X1 port map( B1 => n147, B2 => n514, C1 => n144, C2 => n482, A
                           => n699, ZN => n698);
   U738 : AOI22_X1 port map( A1 => REGISTERS_3_24_port, A2 => n141, B1 => 
                           REGISTERS_2_24_port, B2 => n138, ZN => n699);
   U739 : OAI221_X1 port map( B1 => n195, B2 => n2033, C1 => n192, C2 => n2001,
                           A => n673, ZN => n672);
   U740 : AOI22_X1 port map( A1 => REGISTERS_19_25_port, A2 => n189, B1 => 
                           REGISTERS_18_25_port, B2 => n186, ZN => n673);
   U741 : OAI221_X1 port map( B1 => n147, B2 => n513, C1 => n144, C2 => n481, A
                           => n681, ZN => n680);
   U742 : AOI22_X1 port map( A1 => REGISTERS_3_25_port, A2 => n141, B1 => 
                           REGISTERS_2_25_port, B2 => n138, ZN => n681);
   U743 : OAI221_X1 port map( B1 => n195, B2 => n2032, C1 => n192, C2 => n2000,
                           A => n655, ZN => n654);
   U744 : AOI22_X1 port map( A1 => REGISTERS_19_26_port, A2 => n189, B1 => 
                           REGISTERS_18_26_port, B2 => n186, ZN => n655);
   U745 : OAI221_X1 port map( B1 => n147, B2 => n512, C1 => n144, C2 => n480, A
                           => n663, ZN => n662);
   U746 : AOI22_X1 port map( A1 => REGISTERS_3_26_port, A2 => n141, B1 => 
                           REGISTERS_2_26_port, B2 => n138, ZN => n663);
   U747 : OAI221_X1 port map( B1 => n195, B2 => n2031, C1 => n192, C2 => n1999,
                           A => n637, ZN => n636);
   U748 : AOI22_X1 port map( A1 => REGISTERS_19_27_port, A2 => n189, B1 => 
                           REGISTERS_18_27_port, B2 => n186, ZN => n637);
   U749 : OAI221_X1 port map( B1 => n147, B2 => n511, C1 => n144, C2 => n479, A
                           => n645, ZN => n644);
   U750 : AOI22_X1 port map( A1 => REGISTERS_3_27_port, A2 => n141, B1 => 
                           REGISTERS_2_27_port, B2 => n138, ZN => n645);
   U751 : OAI221_X1 port map( B1 => n195, B2 => n2030, C1 => n192, C2 => n1998,
                           A => n619, ZN => n618);
   U752 : AOI22_X1 port map( A1 => REGISTERS_19_28_port, A2 => n189, B1 => 
                           REGISTERS_18_28_port, B2 => n186, ZN => n619);
   U753 : OAI221_X1 port map( B1 => n147, B2 => n510, C1 => n144, C2 => n478, A
                           => n627, ZN => n626);
   U754 : AOI22_X1 port map( A1 => REGISTERS_3_28_port, A2 => n141, B1 => 
                           REGISTERS_2_28_port, B2 => n138, ZN => n627);
   U755 : OAI221_X1 port map( B1 => n195, B2 => n2029, C1 => n192, C2 => n1997,
                           A => n601, ZN => n600);
   U756 : AOI22_X1 port map( A1 => REGISTERS_19_29_port, A2 => n189, B1 => 
                           REGISTERS_18_29_port, B2 => n186, ZN => n601);
   U757 : OAI221_X1 port map( B1 => n147, B2 => n509, C1 => n144, C2 => n477, A
                           => n609, ZN => n608);
   U758 : AOI22_X1 port map( A1 => REGISTERS_3_29_port, A2 => n141, B1 => 
                           REGISTERS_2_29_port, B2 => n138, ZN => n609);
   U759 : OAI221_X1 port map( B1 => n195, B2 => n2028, C1 => n192, C2 => n1996,
                           A => n583, ZN => n582);
   U760 : AOI22_X1 port map( A1 => REGISTERS_19_30_port, A2 => n189, B1 => 
                           REGISTERS_18_30_port, B2 => n186, ZN => n583);
   U761 : OAI221_X1 port map( B1 => n147, B2 => n508, C1 => n144, C2 => n476, A
                           => n591, ZN => n590);
   U762 : AOI22_X1 port map( A1 => REGISTERS_3_30_port, A2 => n141, B1 => 
                           REGISTERS_2_30_port, B2 => n138, ZN => n591);
   U763 : OAI221_X1 port map( B1 => n195, B2 => n2027, C1 => n192, C2 => n1995,
                           A => n535, ZN => n532);
   U764 : AOI22_X1 port map( A1 => REGISTERS_19_31_port, A2 => n189, B1 => 
                           REGISTERS_18_31_port, B2 => n186, ZN => n535);
   U765 : OAI221_X1 port map( B1 => n147, B2 => n507, C1 => n144, C2 => n475, A
                           => n559, ZN => n556);
   U766 : AOI22_X1 port map( A1 => REGISTERS_3_31_port, A2 => n141, B1 => 
                           REGISTERS_2_31_port, B2 => n138, ZN => n559);
   U767 : OAI221_X1 port map( B1 => n2058, B2 => n97, C1 => n2026, C2 => n94, A
                           => n1748, ZN => n1747);
   U768 : AOI22_X1 port map( A1 => n91, A2 => REGISTERS_19_0_port, B1 => n88, 
                           B2 => REGISTERS_18_0_port, ZN => n1748);
   U769 : OAI221_X1 port map( B1 => n1802, B2 => n49, C1 => n506, C2 => n46, A 
                           => n1766, ZN => n1765);
   U770 : AOI22_X1 port map( A1 => n43, A2 => REGISTERS_3_0_port, B1 => n40, B2
                           => REGISTERS_2_0_port, ZN => n1766);
   U771 : OAI221_X1 port map( B1 => n2057, B2 => n97, C1 => n2025, C2 => n94, A
                           => n1730, ZN => n1729);
   U772 : AOI22_X1 port map( A1 => n91, A2 => REGISTERS_19_1_port, B1 => n88, 
                           B2 => REGISTERS_18_1_port, ZN => n1730);
   U773 : OAI221_X1 port map( B1 => n1801, B2 => n49, C1 => n505, C2 => n46, A 
                           => n1738, ZN => n1737);
   U774 : AOI22_X1 port map( A1 => n43, A2 => REGISTERS_3_1_port, B1 => n40, B2
                           => REGISTERS_2_1_port, ZN => n1738);
   U775 : OAI221_X1 port map( B1 => n2056, B2 => n97, C1 => n2024, C2 => n94, A
                           => n1712, ZN => n1711);
   U776 : AOI22_X1 port map( A1 => n91, A2 => REGISTERS_19_2_port, B1 => n88, 
                           B2 => REGISTERS_18_2_port, ZN => n1712);
   U777 : OAI221_X1 port map( B1 => n1800, B2 => n49, C1 => n504, C2 => n46, A 
                           => n1720, ZN => n1719);
   U778 : AOI22_X1 port map( A1 => n43, A2 => REGISTERS_3_2_port, B1 => n40, B2
                           => REGISTERS_2_2_port, ZN => n1720);
   U779 : OAI221_X1 port map( B1 => n2055, B2 => n97, C1 => n2023, C2 => n94, A
                           => n1694, ZN => n1693);
   U780 : AOI22_X1 port map( A1 => n91, A2 => REGISTERS_19_3_port, B1 => n88, 
                           B2 => REGISTERS_18_3_port, ZN => n1694);
   U781 : OAI221_X1 port map( B1 => n1799, B2 => n49, C1 => n503, C2 => n46, A 
                           => n1702, ZN => n1701);
   U782 : AOI22_X1 port map( A1 => n43, A2 => REGISTERS_3_3_port, B1 => n40, B2
                           => REGISTERS_2_3_port, ZN => n1702);
   U783 : OAI221_X1 port map( B1 => n2054, B2 => n97, C1 => n2022, C2 => n94, A
                           => n1676, ZN => n1675);
   U784 : AOI22_X1 port map( A1 => n91, A2 => REGISTERS_19_4_port, B1 => n88, 
                           B2 => REGISTERS_18_4_port, ZN => n1676);
   U785 : OAI221_X1 port map( B1 => n1798, B2 => n49, C1 => n502, C2 => n46, A 
                           => n1684, ZN => n1683);
   U786 : AOI22_X1 port map( A1 => n43, A2 => REGISTERS_3_4_port, B1 => n40, B2
                           => REGISTERS_2_4_port, ZN => n1684);
   U787 : OAI221_X1 port map( B1 => n2053, B2 => n97, C1 => n2021, C2 => n94, A
                           => n1658, ZN => n1657);
   U788 : AOI22_X1 port map( A1 => n91, A2 => REGISTERS_19_5_port, B1 => n88, 
                           B2 => REGISTERS_18_5_port, ZN => n1658);
   U789 : OAI221_X1 port map( B1 => n1797, B2 => n49, C1 => n501, C2 => n46, A 
                           => n1666, ZN => n1665);
   U790 : AOI22_X1 port map( A1 => n43, A2 => REGISTERS_3_5_port, B1 => n40, B2
                           => REGISTERS_2_5_port, ZN => n1666);
   U791 : OAI221_X1 port map( B1 => n2052, B2 => n97, C1 => n2020, C2 => n94, A
                           => n1640, ZN => n1639);
   U792 : AOI22_X1 port map( A1 => n91, A2 => REGISTERS_19_6_port, B1 => n88, 
                           B2 => REGISTERS_18_6_port, ZN => n1640);
   U793 : OAI221_X1 port map( B1 => n1796, B2 => n49, C1 => n500, C2 => n46, A 
                           => n1648, ZN => n1647);
   U794 : AOI22_X1 port map( A1 => n43, A2 => REGISTERS_3_6_port, B1 => n40, B2
                           => REGISTERS_2_6_port, ZN => n1648);
   U795 : OAI221_X1 port map( B1 => n2051, B2 => n97, C1 => n2019, C2 => n94, A
                           => n1622, ZN => n1621);
   U796 : AOI22_X1 port map( A1 => n91, A2 => REGISTERS_19_7_port, B1 => n88, 
                           B2 => REGISTERS_18_7_port, ZN => n1622);
   U797 : OAI221_X1 port map( B1 => n1795, B2 => n49, C1 => n499, C2 => n46, A 
                           => n1630, ZN => n1629);
   U798 : AOI22_X1 port map( A1 => n43, A2 => REGISTERS_3_7_port, B1 => n40, B2
                           => REGISTERS_2_7_port, ZN => n1630);
   U799 : OAI221_X1 port map( B1 => n2050, B2 => n97, C1 => n2018, C2 => n94, A
                           => n1604, ZN => n1603);
   U800 : AOI22_X1 port map( A1 => n91, A2 => REGISTERS_19_8_port, B1 => n88, 
                           B2 => REGISTERS_18_8_port, ZN => n1604);
   U801 : OAI221_X1 port map( B1 => n1794, B2 => n49, C1 => n498, C2 => n46, A 
                           => n1612, ZN => n1611);
   U802 : AOI22_X1 port map( A1 => n43, A2 => REGISTERS_3_8_port, B1 => n40, B2
                           => REGISTERS_2_8_port, ZN => n1612);
   U803 : OAI221_X1 port map( B1 => n2049, B2 => n97, C1 => n2017, C2 => n94, A
                           => n1586, ZN => n1585);
   U804 : AOI22_X1 port map( A1 => n91, A2 => REGISTERS_19_9_port, B1 => n88, 
                           B2 => REGISTERS_18_9_port, ZN => n1586);
   U805 : OAI221_X1 port map( B1 => n1793, B2 => n49, C1 => n497, C2 => n46, A 
                           => n1594, ZN => n1593);
   U806 : AOI22_X1 port map( A1 => n43, A2 => REGISTERS_3_9_port, B1 => n40, B2
                           => REGISTERS_2_9_port, ZN => n1594);
   U807 : OAI221_X1 port map( B1 => n2048, B2 => n97, C1 => n2016, C2 => n94, A
                           => n1568, ZN => n1567);
   U808 : AOI22_X1 port map( A1 => n91, A2 => REGISTERS_19_10_port, B1 => n88, 
                           B2 => REGISTERS_18_10_port, ZN => n1568);
   U809 : OAI221_X1 port map( B1 => n1792, B2 => n49, C1 => n496, C2 => n46, A 
                           => n1576, ZN => n1575);
   U810 : AOI22_X1 port map( A1 => n43, A2 => REGISTERS_3_10_port, B1 => n40, 
                           B2 => REGISTERS_2_10_port, ZN => n1576);
   U811 : OAI221_X1 port map( B1 => n2036, B2 => n99, C1 => n2004, C2 => n96, A
                           => n1352, ZN => n1351);
   U812 : AOI22_X1 port map( A1 => n93, A2 => REGISTERS_19_22_port, B1 => n90, 
                           B2 => REGISTERS_18_22_port, ZN => n1352);
   U813 : OAI221_X1 port map( B1 => n516, B2 => n51, C1 => n484, C2 => n48, A 
                           => n1360, ZN => n1359);
   U814 : AOI22_X1 port map( A1 => n45, A2 => REGISTERS_3_22_port, B1 => n42, 
                           B2 => REGISTERS_2_22_port, ZN => n1360);
   U815 : OAI221_X1 port map( B1 => n2035, B2 => n99, C1 => n2003, C2 => n96, A
                           => n1334, ZN => n1333);
   U816 : AOI22_X1 port map( A1 => n93, A2 => REGISTERS_19_23_port, B1 => n90, 
                           B2 => REGISTERS_18_23_port, ZN => n1334);
   U817 : OAI221_X1 port map( B1 => n515, B2 => n51, C1 => n483, C2 => n48, A 
                           => n1342, ZN => n1341);
   U818 : AOI22_X1 port map( A1 => n45, A2 => REGISTERS_3_23_port, B1 => n42, 
                           B2 => REGISTERS_2_23_port, ZN => n1342);
   U819 : OAI221_X1 port map( B1 => n2034, B2 => n99, C1 => n2002, C2 => n96, A
                           => n1316, ZN => n1315);
   U820 : AOI22_X1 port map( A1 => n93, A2 => REGISTERS_19_24_port, B1 => n90, 
                           B2 => REGISTERS_18_24_port, ZN => n1316);
   U821 : OAI221_X1 port map( B1 => n514, B2 => n51, C1 => n482, C2 => n48, A 
                           => n1324, ZN => n1323);
   U822 : AOI22_X1 port map( A1 => n45, A2 => REGISTERS_3_24_port, B1 => n42, 
                           B2 => REGISTERS_2_24_port, ZN => n1324);
   U823 : OAI221_X1 port map( B1 => n2033, B2 => n99, C1 => n2001, C2 => n96, A
                           => n1298, ZN => n1297);
   U824 : AOI22_X1 port map( A1 => n93, A2 => REGISTERS_19_25_port, B1 => n90, 
                           B2 => REGISTERS_18_25_port, ZN => n1298);
   U825 : OAI221_X1 port map( B1 => n513, B2 => n51, C1 => n481, C2 => n48, A 
                           => n1306, ZN => n1305);
   U826 : AOI22_X1 port map( A1 => n45, A2 => REGISTERS_3_25_port, B1 => n42, 
                           B2 => REGISTERS_2_25_port, ZN => n1306);
   U827 : OAI221_X1 port map( B1 => n2032, B2 => n99, C1 => n2000, C2 => n96, A
                           => n1280, ZN => n1279);
   U828 : AOI22_X1 port map( A1 => n93, A2 => REGISTERS_19_26_port, B1 => n90, 
                           B2 => REGISTERS_18_26_port, ZN => n1280);
   U829 : OAI221_X1 port map( B1 => n512, B2 => n51, C1 => n480, C2 => n48, A 
                           => n1288, ZN => n1287);
   U830 : AOI22_X1 port map( A1 => n45, A2 => REGISTERS_3_26_port, B1 => n42, 
                           B2 => REGISTERS_2_26_port, ZN => n1288);
   U831 : OAI221_X1 port map( B1 => n2031, B2 => n99, C1 => n1999, C2 => n96, A
                           => n1262, ZN => n1261);
   U832 : AOI22_X1 port map( A1 => n93, A2 => REGISTERS_19_27_port, B1 => n90, 
                           B2 => REGISTERS_18_27_port, ZN => n1262);
   U833 : OAI221_X1 port map( B1 => n511, B2 => n51, C1 => n479, C2 => n48, A 
                           => n1270, ZN => n1269);
   U834 : AOI22_X1 port map( A1 => n45, A2 => REGISTERS_3_27_port, B1 => n42, 
                           B2 => REGISTERS_2_27_port, ZN => n1270);
   U835 : OAI221_X1 port map( B1 => n2030, B2 => n99, C1 => n1998, C2 => n96, A
                           => n1244, ZN => n1243);
   U836 : AOI22_X1 port map( A1 => n93, A2 => REGISTERS_19_28_port, B1 => n90, 
                           B2 => REGISTERS_18_28_port, ZN => n1244);
   U837 : OAI221_X1 port map( B1 => n510, B2 => n51, C1 => n478, C2 => n48, A 
                           => n1252, ZN => n1251);
   U838 : AOI22_X1 port map( A1 => n45, A2 => REGISTERS_3_28_port, B1 => n42, 
                           B2 => REGISTERS_2_28_port, ZN => n1252);
   U839 : OAI221_X1 port map( B1 => n2029, B2 => n99, C1 => n1997, C2 => n96, A
                           => n1226, ZN => n1225);
   U840 : AOI22_X1 port map( A1 => n93, A2 => REGISTERS_19_29_port, B1 => n90, 
                           B2 => REGISTERS_18_29_port, ZN => n1226);
   U841 : OAI221_X1 port map( B1 => n509, B2 => n51, C1 => n477, C2 => n48, A 
                           => n1234, ZN => n1233);
   U842 : AOI22_X1 port map( A1 => n45, A2 => REGISTERS_3_29_port, B1 => n42, 
                           B2 => REGISTERS_2_29_port, ZN => n1234);
   U843 : OAI221_X1 port map( B1 => n2028, B2 => n99, C1 => n1996, C2 => n96, A
                           => n1208, ZN => n1207);
   U844 : AOI22_X1 port map( A1 => n93, A2 => REGISTERS_19_30_port, B1 => n90, 
                           B2 => REGISTERS_18_30_port, ZN => n1208);
   U845 : OAI221_X1 port map( B1 => n508, B2 => n51, C1 => n476, C2 => n48, A 
                           => n1216, ZN => n1215);
   U846 : AOI22_X1 port map( A1 => n45, A2 => REGISTERS_3_30_port, B1 => n42, 
                           B2 => REGISTERS_2_30_port, ZN => n1216);
   U847 : OAI221_X1 port map( B1 => n2027, B2 => n99, C1 => n1995, C2 => n96, A
                           => n1160, ZN => n1157);
   U848 : AOI22_X1 port map( A1 => n93, A2 => REGISTERS_19_31_port, B1 => n90, 
                           B2 => REGISTERS_18_31_port, ZN => n1160);
   U849 : OAI221_X1 port map( B1 => n507, B2 => n51, C1 => n475, C2 => n48, A 
                           => n1184, ZN => n1181);
   U850 : AOI22_X1 port map( A1 => n45, A2 => REGISTERS_3_31_port, B1 => n42, 
                           B2 => REGISTERS_2_31_port, ZN => n1184);
   U851 : OAI221_X1 port map( B1 => n183, B2 => n2098, C1 => n180, C2 => n2066,
                           A => n692, ZN => n689);
   U852 : AOI22_X1 port map( A1 => REGISTERS_23_24_port, A2 => n177, B1 => 
                           REGISTERS_22_24_port, B2 => n174, ZN => n692);
   U853 : OAI221_X1 port map( B1 => n135, B2 => n1842, C1 => n132, C2 => n1810,
                           A => n700, ZN => n697);
   U854 : AOI22_X1 port map( A1 => REGISTERS_7_24_port, A2 => n129, B1 => 
                           REGISTERS_6_24_port, B2 => n126, ZN => n700);
   U855 : OAI221_X1 port map( B1 => n183, B2 => n2097, C1 => n180, C2 => n2065,
                           A => n674, ZN => n671);
   U856 : AOI22_X1 port map( A1 => REGISTERS_23_25_port, A2 => n177, B1 => 
                           REGISTERS_22_25_port, B2 => n174, ZN => n674);
   U857 : OAI221_X1 port map( B1 => n135, B2 => n1841, C1 => n132, C2 => n1809,
                           A => n682, ZN => n679);
   U858 : AOI22_X1 port map( A1 => REGISTERS_7_25_port, A2 => n129, B1 => 
                           REGISTERS_6_25_port, B2 => n126, ZN => n682);
   U859 : OAI221_X1 port map( B1 => n183, B2 => n2096, C1 => n180, C2 => n2064,
                           A => n656, ZN => n653);
   U860 : AOI22_X1 port map( A1 => REGISTERS_23_26_port, A2 => n177, B1 => 
                           REGISTERS_22_26_port, B2 => n174, ZN => n656);
   U861 : OAI221_X1 port map( B1 => n135, B2 => n1840, C1 => n132, C2 => n1808,
                           A => n664, ZN => n661);
   U862 : AOI22_X1 port map( A1 => REGISTERS_7_26_port, A2 => n129, B1 => 
                           REGISTERS_6_26_port, B2 => n126, ZN => n664);
   U863 : OAI221_X1 port map( B1 => n183, B2 => n2095, C1 => n180, C2 => n2063,
                           A => n638, ZN => n635);
   U864 : AOI22_X1 port map( A1 => REGISTERS_23_27_port, A2 => n177, B1 => 
                           REGISTERS_22_27_port, B2 => n174, ZN => n638);
   U865 : OAI221_X1 port map( B1 => n135, B2 => n1839, C1 => n132, C2 => n1807,
                           A => n646, ZN => n643);
   U866 : AOI22_X1 port map( A1 => REGISTERS_7_27_port, A2 => n129, B1 => 
                           REGISTERS_6_27_port, B2 => n126, ZN => n646);
   U867 : OAI221_X1 port map( B1 => n183, B2 => n2094, C1 => n180, C2 => n2062,
                           A => n620, ZN => n617);
   U868 : AOI22_X1 port map( A1 => REGISTERS_23_28_port, A2 => n177, B1 => 
                           REGISTERS_22_28_port, B2 => n174, ZN => n620);
   U869 : OAI221_X1 port map( B1 => n135, B2 => n1838, C1 => n132, C2 => n1806,
                           A => n628, ZN => n625);
   U870 : AOI22_X1 port map( A1 => REGISTERS_7_28_port, A2 => n129, B1 => 
                           REGISTERS_6_28_port, B2 => n126, ZN => n628);
   U871 : OAI221_X1 port map( B1 => n183, B2 => n2093, C1 => n180, C2 => n2061,
                           A => n602, ZN => n599);
   U872 : AOI22_X1 port map( A1 => REGISTERS_23_29_port, A2 => n177, B1 => 
                           REGISTERS_22_29_port, B2 => n174, ZN => n602);
   U873 : OAI221_X1 port map( B1 => n135, B2 => n1837, C1 => n132, C2 => n1805,
                           A => n610, ZN => n607);
   U874 : AOI22_X1 port map( A1 => REGISTERS_7_29_port, A2 => n129, B1 => 
                           REGISTERS_6_29_port, B2 => n126, ZN => n610);
   U875 : OAI221_X1 port map( B1 => n183, B2 => n2092, C1 => n180, C2 => n2060,
                           A => n584, ZN => n581);
   U876 : AOI22_X1 port map( A1 => REGISTERS_23_30_port, A2 => n177, B1 => 
                           REGISTERS_22_30_port, B2 => n174, ZN => n584);
   U877 : OAI221_X1 port map( B1 => n135, B2 => n1836, C1 => n132, C2 => n1804,
                           A => n592, ZN => n589);
   U878 : AOI22_X1 port map( A1 => REGISTERS_7_30_port, A2 => n129, B1 => 
                           REGISTERS_6_30_port, B2 => n126, ZN => n592);
   U879 : OAI221_X1 port map( B1 => n183, B2 => n2091, C1 => n180, C2 => n2059,
                           A => n540, ZN => n531);
   U880 : AOI22_X1 port map( A1 => REGISTERS_23_31_port, A2 => n177, B1 => 
                           REGISTERS_22_31_port, B2 => n174, ZN => n540);
   U881 : OAI221_X1 port map( B1 => n135, B2 => n1835, C1 => n132, C2 => n1803,
                           A => n564, ZN => n555);
   U882 : AOI22_X1 port map( A1 => REGISTERS_7_31_port, A2 => n129, B1 => 
                           REGISTERS_6_31_port, B2 => n126, ZN => n564);
   U883 : OAI221_X1 port map( B1 => n193, B2 => n2058, C1 => n190, C2 => n2026,
                           A => n1123, ZN => n1122);
   U884 : AOI22_X1 port map( A1 => REGISTERS_19_0_port, A2 => n187, B1 => 
                           REGISTERS_18_0_port, B2 => n184, ZN => n1123);
   U885 : OAI221_X1 port map( B1 => n145, B2 => n1802, C1 => n142, C2 => n506, 
                           A => n1141, ZN => n1140);
   U886 : AOI22_X1 port map( A1 => REGISTERS_3_0_port, A2 => n139, B1 => 
                           REGISTERS_2_0_port, B2 => n136, ZN => n1141);
   U887 : OAI221_X1 port map( B1 => n193, B2 => n2057, C1 => n190, C2 => n2025,
                           A => n1105, ZN => n1104);
   U888 : AOI22_X1 port map( A1 => REGISTERS_19_1_port, A2 => n187, B1 => 
                           REGISTERS_18_1_port, B2 => n184, ZN => n1105);
   U889 : OAI221_X1 port map( B1 => n145, B2 => n1801, C1 => n142, C2 => n505, 
                           A => n1113, ZN => n1112);
   U890 : AOI22_X1 port map( A1 => REGISTERS_3_1_port, A2 => n139, B1 => 
                           REGISTERS_2_1_port, B2 => n136, ZN => n1113);
   U891 : OAI221_X1 port map( B1 => n193, B2 => n2056, C1 => n190, C2 => n2024,
                           A => n1087, ZN => n1086);
   U892 : AOI22_X1 port map( A1 => REGISTERS_19_2_port, A2 => n187, B1 => 
                           REGISTERS_18_2_port, B2 => n184, ZN => n1087);
   U893 : OAI221_X1 port map( B1 => n145, B2 => n1800, C1 => n142, C2 => n504, 
                           A => n1095, ZN => n1094);
   U894 : AOI22_X1 port map( A1 => REGISTERS_3_2_port, A2 => n139, B1 => 
                           REGISTERS_2_2_port, B2 => n136, ZN => n1095);
   U895 : OAI221_X1 port map( B1 => n193, B2 => n2055, C1 => n190, C2 => n2023,
                           A => n1069, ZN => n1068);
   U896 : AOI22_X1 port map( A1 => REGISTERS_19_3_port, A2 => n187, B1 => 
                           REGISTERS_18_3_port, B2 => n184, ZN => n1069);
   U897 : OAI221_X1 port map( B1 => n145, B2 => n1799, C1 => n142, C2 => n503, 
                           A => n1077, ZN => n1076);
   U898 : AOI22_X1 port map( A1 => REGISTERS_3_3_port, A2 => n139, B1 => 
                           REGISTERS_2_3_port, B2 => n136, ZN => n1077);
   U899 : OAI221_X1 port map( B1 => n193, B2 => n2054, C1 => n190, C2 => n2022,
                           A => n1051, ZN => n1050);
   U900 : AOI22_X1 port map( A1 => REGISTERS_19_4_port, A2 => n187, B1 => 
                           REGISTERS_18_4_port, B2 => n184, ZN => n1051);
   U901 : OAI221_X1 port map( B1 => n145, B2 => n1798, C1 => n142, C2 => n502, 
                           A => n1059, ZN => n1058);
   U902 : AOI22_X1 port map( A1 => REGISTERS_3_4_port, A2 => n139, B1 => 
                           REGISTERS_2_4_port, B2 => n136, ZN => n1059);
   U903 : OAI221_X1 port map( B1 => n193, B2 => n2053, C1 => n190, C2 => n2021,
                           A => n1033, ZN => n1032);
   U904 : AOI22_X1 port map( A1 => REGISTERS_19_5_port, A2 => n187, B1 => 
                           REGISTERS_18_5_port, B2 => n184, ZN => n1033);
   U905 : OAI221_X1 port map( B1 => n145, B2 => n1797, C1 => n142, C2 => n501, 
                           A => n1041, ZN => n1040);
   U906 : AOI22_X1 port map( A1 => REGISTERS_3_5_port, A2 => n139, B1 => 
                           REGISTERS_2_5_port, B2 => n136, ZN => n1041);
   U907 : OAI221_X1 port map( B1 => n193, B2 => n2052, C1 => n190, C2 => n2020,
                           A => n1015, ZN => n1014);
   U908 : AOI22_X1 port map( A1 => REGISTERS_19_6_port, A2 => n187, B1 => 
                           REGISTERS_18_6_port, B2 => n184, ZN => n1015);
   U909 : OAI221_X1 port map( B1 => n145, B2 => n1796, C1 => n142, C2 => n500, 
                           A => n1023, ZN => n1022);
   U910 : AOI22_X1 port map( A1 => REGISTERS_3_6_port, A2 => n139, B1 => 
                           REGISTERS_2_6_port, B2 => n136, ZN => n1023);
   U911 : OAI221_X1 port map( B1 => n193, B2 => n2051, C1 => n190, C2 => n2019,
                           A => n997, ZN => n996);
   U912 : AOI22_X1 port map( A1 => REGISTERS_19_7_port, A2 => n187, B1 => 
                           REGISTERS_18_7_port, B2 => n184, ZN => n997);
   U913 : OAI221_X1 port map( B1 => n145, B2 => n1795, C1 => n142, C2 => n499, 
                           A => n1005, ZN => n1004);
   U914 : AOI22_X1 port map( A1 => REGISTERS_3_7_port, A2 => n139, B1 => 
                           REGISTERS_2_7_port, B2 => n136, ZN => n1005);
   U915 : OAI221_X1 port map( B1 => n193, B2 => n2050, C1 => n190, C2 => n2018,
                           A => n979, ZN => n978);
   U916 : AOI22_X1 port map( A1 => REGISTERS_19_8_port, A2 => n187, B1 => 
                           REGISTERS_18_8_port, B2 => n184, ZN => n979);
   U917 : OAI221_X1 port map( B1 => n145, B2 => n1794, C1 => n142, C2 => n498, 
                           A => n987, ZN => n986);
   U918 : AOI22_X1 port map( A1 => REGISTERS_3_8_port, A2 => n139, B1 => 
                           REGISTERS_2_8_port, B2 => n136, ZN => n987);
   U919 : OAI221_X1 port map( B1 => n193, B2 => n2049, C1 => n190, C2 => n2017,
                           A => n961, ZN => n960);
   U920 : AOI22_X1 port map( A1 => REGISTERS_19_9_port, A2 => n187, B1 => 
                           REGISTERS_18_9_port, B2 => n184, ZN => n961);
   U921 : OAI221_X1 port map( B1 => n145, B2 => n1793, C1 => n142, C2 => n497, 
                           A => n969, ZN => n968);
   U922 : AOI22_X1 port map( A1 => REGISTERS_3_9_port, A2 => n139, B1 => 
                           REGISTERS_2_9_port, B2 => n136, ZN => n969);
   U923 : OAI221_X1 port map( B1 => n193, B2 => n2048, C1 => n190, C2 => n2016,
                           A => n943, ZN => n942);
   U924 : AOI22_X1 port map( A1 => REGISTERS_19_10_port, A2 => n187, B1 => 
                           REGISTERS_18_10_port, B2 => n184, ZN => n943);
   U925 : OAI221_X1 port map( B1 => n145, B2 => n1792, C1 => n142, C2 => n496, 
                           A => n951, ZN => n950);
   U926 : AOI22_X1 port map( A1 => REGISTERS_3_10_port, A2 => n139, B1 => 
                           REGISTERS_2_10_port, B2 => n136, ZN => n951);
   U927 : OAI221_X1 port map( B1 => n193, B2 => n2047, C1 => n191, C2 => n2015,
                           A => n925, ZN => n924);
   U928 : AOI22_X1 port map( A1 => REGISTERS_19_11_port, A2 => n187, B1 => 
                           REGISTERS_18_11_port, B2 => n184, ZN => n925);
   U929 : OAI221_X1 port map( B1 => n145, B2 => n1791, C1 => n143, C2 => n495, 
                           A => n933, ZN => n932);
   U930 : AOI22_X1 port map( A1 => REGISTERS_3_11_port, A2 => n139, B1 => 
                           REGISTERS_2_11_port, B2 => n136, ZN => n933);
   U931 : OAI221_X1 port map( B1 => n194, B2 => n2046, C1 => n191, C2 => n2014,
                           A => n907, ZN => n906);
   U932 : AOI22_X1 port map( A1 => REGISTERS_19_12_port, A2 => n188, B1 => 
                           REGISTERS_18_12_port, B2 => n185, ZN => n907);
   U933 : OAI221_X1 port map( B1 => n146, B2 => n526, C1 => n143, C2 => n494, A
                           => n915, ZN => n914);
   U934 : AOI22_X1 port map( A1 => REGISTERS_3_12_port, A2 => n140, B1 => 
                           REGISTERS_2_12_port, B2 => n137, ZN => n915);
   U935 : OAI221_X1 port map( B1 => n194, B2 => n2045, C1 => n191, C2 => n2013,
                           A => n889, ZN => n888);
   U936 : AOI22_X1 port map( A1 => REGISTERS_19_13_port, A2 => n188, B1 => 
                           REGISTERS_18_13_port, B2 => n185, ZN => n889);
   U937 : OAI221_X1 port map( B1 => n146, B2 => n525, C1 => n143, C2 => n493, A
                           => n897, ZN => n896);
   U938 : AOI22_X1 port map( A1 => REGISTERS_3_13_port, A2 => n140, B1 => 
                           REGISTERS_2_13_port, B2 => n137, ZN => n897);
   U939 : OAI221_X1 port map( B1 => n194, B2 => n2044, C1 => n191, C2 => n2012,
                           A => n871, ZN => n870);
   U940 : AOI22_X1 port map( A1 => REGISTERS_19_14_port, A2 => n188, B1 => 
                           REGISTERS_18_14_port, B2 => n185, ZN => n871);
   U941 : OAI221_X1 port map( B1 => n146, B2 => n524, C1 => n143, C2 => n492, A
                           => n879, ZN => n878);
   U942 : AOI22_X1 port map( A1 => REGISTERS_3_14_port, A2 => n140, B1 => 
                           REGISTERS_2_14_port, B2 => n137, ZN => n879);
   U943 : OAI221_X1 port map( B1 => n194, B2 => n2043, C1 => n191, C2 => n2011,
                           A => n853, ZN => n852);
   U944 : AOI22_X1 port map( A1 => REGISTERS_19_15_port, A2 => n188, B1 => 
                           REGISTERS_18_15_port, B2 => n185, ZN => n853);
   U945 : OAI221_X1 port map( B1 => n146, B2 => n523, C1 => n143, C2 => n491, A
                           => n861, ZN => n860);
   U946 : AOI22_X1 port map( A1 => REGISTERS_3_15_port, A2 => n140, B1 => 
                           REGISTERS_2_15_port, B2 => n137, ZN => n861);
   U947 : OAI221_X1 port map( B1 => n194, B2 => n2042, C1 => n191, C2 => n2010,
                           A => n835, ZN => n834);
   U948 : AOI22_X1 port map( A1 => REGISTERS_19_16_port, A2 => n188, B1 => 
                           REGISTERS_18_16_port, B2 => n185, ZN => n835);
   U949 : OAI221_X1 port map( B1 => n146, B2 => n522, C1 => n143, C2 => n490, A
                           => n843, ZN => n842);
   U950 : AOI22_X1 port map( A1 => REGISTERS_3_16_port, A2 => n140, B1 => 
                           REGISTERS_2_16_port, B2 => n137, ZN => n843);
   U951 : OAI221_X1 port map( B1 => n194, B2 => n2041, C1 => n191, C2 => n2009,
                           A => n817, ZN => n816);
   U952 : AOI22_X1 port map( A1 => REGISTERS_19_17_port, A2 => n188, B1 => 
                           REGISTERS_18_17_port, B2 => n185, ZN => n817);
   U953 : OAI221_X1 port map( B1 => n146, B2 => n521, C1 => n143, C2 => n489, A
                           => n825, ZN => n824);
   U954 : AOI22_X1 port map( A1 => REGISTERS_3_17_port, A2 => n140, B1 => 
                           REGISTERS_2_17_port, B2 => n137, ZN => n825);
   U955 : OAI221_X1 port map( B1 => n194, B2 => n2040, C1 => n191, C2 => n2008,
                           A => n799, ZN => n798);
   U956 : AOI22_X1 port map( A1 => REGISTERS_19_18_port, A2 => n188, B1 => 
                           REGISTERS_18_18_port, B2 => n185, ZN => n799);
   U957 : OAI221_X1 port map( B1 => n146, B2 => n520, C1 => n143, C2 => n488, A
                           => n807, ZN => n806);
   U958 : AOI22_X1 port map( A1 => REGISTERS_3_18_port, A2 => n140, B1 => 
                           REGISTERS_2_18_port, B2 => n137, ZN => n807);
   U959 : OAI221_X1 port map( B1 => n194, B2 => n2039, C1 => n191, C2 => n2007,
                           A => n781, ZN => n780);
   U960 : AOI22_X1 port map( A1 => REGISTERS_19_19_port, A2 => n188, B1 => 
                           REGISTERS_18_19_port, B2 => n185, ZN => n781);
   U961 : OAI221_X1 port map( B1 => n146, B2 => n519, C1 => n143, C2 => n487, A
                           => n789, ZN => n788);
   U962 : AOI22_X1 port map( A1 => REGISTERS_3_19_port, A2 => n140, B1 => 
                           REGISTERS_2_19_port, B2 => n137, ZN => n789);
   U963 : OAI221_X1 port map( B1 => n194, B2 => n2038, C1 => n191, C2 => n2006,
                           A => n763, ZN => n762);
   U964 : AOI22_X1 port map( A1 => REGISTERS_19_20_port, A2 => n188, B1 => 
                           REGISTERS_18_20_port, B2 => n185, ZN => n763);
   U965 : OAI221_X1 port map( B1 => n146, B2 => n518, C1 => n143, C2 => n486, A
                           => n771, ZN => n770);
   U966 : AOI22_X1 port map( A1 => REGISTERS_3_20_port, A2 => n140, B1 => 
                           REGISTERS_2_20_port, B2 => n137, ZN => n771);
   U967 : OAI221_X1 port map( B1 => n194, B2 => n2037, C1 => n191, C2 => n2005,
                           A => n745, ZN => n744);
   U968 : AOI22_X1 port map( A1 => REGISTERS_19_21_port, A2 => n188, B1 => 
                           REGISTERS_18_21_port, B2 => n185, ZN => n745);
   U969 : OAI221_X1 port map( B1 => n146, B2 => n517, C1 => n143, C2 => n485, A
                           => n753, ZN => n752);
   U970 : AOI22_X1 port map( A1 => REGISTERS_3_21_port, A2 => n140, B1 => 
                           REGISTERS_2_21_port, B2 => n137, ZN => n753);
   U971 : OAI221_X1 port map( B1 => n194, B2 => n2036, C1 => n192, C2 => n2004,
                           A => n727, ZN => n726);
   U972 : AOI22_X1 port map( A1 => REGISTERS_19_22_port, A2 => n188, B1 => 
                           REGISTERS_18_22_port, B2 => n185, ZN => n727);
   U973 : OAI221_X1 port map( B1 => n146, B2 => n516, C1 => n144, C2 => n484, A
                           => n735, ZN => n734);
   U974 : AOI22_X1 port map( A1 => REGISTERS_3_22_port, A2 => n140, B1 => 
                           REGISTERS_2_22_port, B2 => n137, ZN => n735);
   U975 : OAI221_X1 port map( B1 => n194, B2 => n2035, C1 => n192, C2 => n2003,
                           A => n709, ZN => n708);
   U976 : AOI22_X1 port map( A1 => REGISTERS_19_23_port, A2 => n188, B1 => 
                           REGISTERS_18_23_port, B2 => n185, ZN => n709);
   U977 : OAI221_X1 port map( B1 => n146, B2 => n515, C1 => n144, C2 => n483, A
                           => n717, ZN => n716);
   U978 : AOI22_X1 port map( A1 => REGISTERS_3_23_port, A2 => n140, B1 => 
                           REGISTERS_2_23_port, B2 => n137, ZN => n717);
   U979 : OAI221_X1 port map( B1 => n2047, B2 => n98, C1 => n2015, C2 => n95, A
                           => n1550, ZN => n1549);
   U980 : AOI22_X1 port map( A1 => n92, A2 => REGISTERS_19_11_port, B1 => n89, 
                           B2 => REGISTERS_18_11_port, ZN => n1550);
   U981 : OAI221_X1 port map( B1 => n1791, B2 => n50, C1 => n495, C2 => n47, A 
                           => n1558, ZN => n1557);
   U982 : AOI22_X1 port map( A1 => n44, A2 => REGISTERS_3_11_port, B1 => n41, 
                           B2 => REGISTERS_2_11_port, ZN => n1558);
   U983 : OAI221_X1 port map( B1 => n2046, B2 => n98, C1 => n2014, C2 => n95, A
                           => n1532, ZN => n1531);
   U984 : AOI22_X1 port map( A1 => n92, A2 => REGISTERS_19_12_port, B1 => n89, 
                           B2 => REGISTERS_18_12_port, ZN => n1532);
   U985 : OAI221_X1 port map( B1 => n526, B2 => n50, C1 => n494, C2 => n47, A 
                           => n1540, ZN => n1539);
   U986 : AOI22_X1 port map( A1 => n44, A2 => REGISTERS_3_12_port, B1 => n41, 
                           B2 => REGISTERS_2_12_port, ZN => n1540);
   U987 : OAI221_X1 port map( B1 => n2045, B2 => n98, C1 => n2013, C2 => n95, A
                           => n1514, ZN => n1513);
   U988 : AOI22_X1 port map( A1 => n92, A2 => REGISTERS_19_13_port, B1 => n89, 
                           B2 => REGISTERS_18_13_port, ZN => n1514);
   U989 : OAI221_X1 port map( B1 => n525, B2 => n50, C1 => n493, C2 => n47, A 
                           => n1522, ZN => n1521);
   U990 : AOI22_X1 port map( A1 => n44, A2 => REGISTERS_3_13_port, B1 => n41, 
                           B2 => REGISTERS_2_13_port, ZN => n1522);
   U991 : OAI221_X1 port map( B1 => n2044, B2 => n98, C1 => n2012, C2 => n95, A
                           => n1496, ZN => n1495);
   U992 : AOI22_X1 port map( A1 => n92, A2 => REGISTERS_19_14_port, B1 => n89, 
                           B2 => REGISTERS_18_14_port, ZN => n1496);
   U993 : OAI221_X1 port map( B1 => n524, B2 => n50, C1 => n492, C2 => n47, A 
                           => n1504, ZN => n1503);
   U994 : AOI22_X1 port map( A1 => n44, A2 => REGISTERS_3_14_port, B1 => n41, 
                           B2 => REGISTERS_2_14_port, ZN => n1504);
   U995 : OAI221_X1 port map( B1 => n2043, B2 => n98, C1 => n2011, C2 => n95, A
                           => n1478, ZN => n1477);
   U996 : AOI22_X1 port map( A1 => n92, A2 => REGISTERS_19_15_port, B1 => n89, 
                           B2 => REGISTERS_18_15_port, ZN => n1478);
   U997 : OAI221_X1 port map( B1 => n523, B2 => n50, C1 => n491, C2 => n47, A 
                           => n1486, ZN => n1485);
   U998 : AOI22_X1 port map( A1 => n44, A2 => REGISTERS_3_15_port, B1 => n41, 
                           B2 => REGISTERS_2_15_port, ZN => n1486);
   U999 : OAI221_X1 port map( B1 => n2042, B2 => n98, C1 => n2010, C2 => n95, A
                           => n1460, ZN => n1459);
   U1000 : AOI22_X1 port map( A1 => n92, A2 => REGISTERS_19_16_port, B1 => n89,
                           B2 => REGISTERS_18_16_port, ZN => n1460);
   U1001 : OAI221_X1 port map( B1 => n522, B2 => n50, C1 => n490, C2 => n47, A 
                           => n1468, ZN => n1467);
   U1002 : AOI22_X1 port map( A1 => n44, A2 => REGISTERS_3_16_port, B1 => n41, 
                           B2 => REGISTERS_2_16_port, ZN => n1468);
   U1003 : OAI221_X1 port map( B1 => n2041, B2 => n98, C1 => n2009, C2 => n95, 
                           A => n1442, ZN => n1441);
   U1004 : AOI22_X1 port map( A1 => n92, A2 => REGISTERS_19_17_port, B1 => n89,
                           B2 => REGISTERS_18_17_port, ZN => n1442);
   U1005 : OAI221_X1 port map( B1 => n521, B2 => n50, C1 => n489, C2 => n47, A 
                           => n1450, ZN => n1449);
   U1006 : AOI22_X1 port map( A1 => n44, A2 => REGISTERS_3_17_port, B1 => n41, 
                           B2 => REGISTERS_2_17_port, ZN => n1450);
   U1007 : OAI221_X1 port map( B1 => n2040, B2 => n98, C1 => n2008, C2 => n95, 
                           A => n1424, ZN => n1423);
   U1008 : AOI22_X1 port map( A1 => n92, A2 => REGISTERS_19_18_port, B1 => n89,
                           B2 => REGISTERS_18_18_port, ZN => n1424);
   U1009 : OAI221_X1 port map( B1 => n520, B2 => n50, C1 => n488, C2 => n47, A 
                           => n1432, ZN => n1431);
   U1010 : AOI22_X1 port map( A1 => n44, A2 => REGISTERS_3_18_port, B1 => n41, 
                           B2 => REGISTERS_2_18_port, ZN => n1432);
   U1011 : OAI221_X1 port map( B1 => n2039, B2 => n98, C1 => n2007, C2 => n95, 
                           A => n1406, ZN => n1405);
   U1012 : AOI22_X1 port map( A1 => n92, A2 => REGISTERS_19_19_port, B1 => n89,
                           B2 => REGISTERS_18_19_port, ZN => n1406);
   U1013 : OAI221_X1 port map( B1 => n519, B2 => n50, C1 => n487, C2 => n47, A 
                           => n1414, ZN => n1413);
   U1014 : AOI22_X1 port map( A1 => n44, A2 => REGISTERS_3_19_port, B1 => n41, 
                           B2 => REGISTERS_2_19_port, ZN => n1414);
   U1015 : OAI221_X1 port map( B1 => n2038, B2 => n98, C1 => n2006, C2 => n95, 
                           A => n1388, ZN => n1387);
   U1016 : AOI22_X1 port map( A1 => n92, A2 => REGISTERS_19_20_port, B1 => n89,
                           B2 => REGISTERS_18_20_port, ZN => n1388);
   U1017 : OAI221_X1 port map( B1 => n518, B2 => n50, C1 => n486, C2 => n47, A 
                           => n1396, ZN => n1395);
   U1018 : AOI22_X1 port map( A1 => n44, A2 => REGISTERS_3_20_port, B1 => n41, 
                           B2 => REGISTERS_2_20_port, ZN => n1396);
   U1019 : OAI221_X1 port map( B1 => n2037, B2 => n98, C1 => n2005, C2 => n95, 
                           A => n1370, ZN => n1369);
   U1020 : AOI22_X1 port map( A1 => n92, A2 => REGISTERS_19_21_port, B1 => n89,
                           B2 => REGISTERS_18_21_port, ZN => n1370);
   U1021 : OAI221_X1 port map( B1 => n517, B2 => n50, C1 => n485, C2 => n47, A 
                           => n1378, ZN => n1377);
   U1022 : AOI22_X1 port map( A1 => n44, A2 => REGISTERS_3_21_port, B1 => n41, 
                           B2 => REGISTERS_2_21_port, ZN => n1378);
   U1023 : OAI221_X1 port map( B1 => n2122, B2 => n85, C1 => n2090, C2 => n82, 
                           A => n1753, ZN => n1746);
   U1024 : AOI22_X1 port map( A1 => n79, A2 => REGISTERS_23_0_port, B1 => n76, 
                           B2 => REGISTERS_22_0_port, ZN => n1753);
   U1025 : OAI221_X1 port map( B1 => n1866, B2 => n37, C1 => n1834, C2 => n34, 
                           A => n1769, ZN => n1764);
   U1026 : AOI22_X1 port map( A1 => n31, A2 => REGISTERS_7_0_port, B1 => n28, 
                           B2 => REGISTERS_6_0_port, ZN => n1769);
   U1027 : OAI221_X1 port map( B1 => n2121, B2 => n85, C1 => n2089, C2 => n82, 
                           A => n1731, ZN => n1728);
   U1028 : AOI22_X1 port map( A1 => n79, A2 => REGISTERS_23_1_port, B1 => n76, 
                           B2 => REGISTERS_22_1_port, ZN => n1731);
   U1029 : OAI221_X1 port map( B1 => n1865, B2 => n37, C1 => n1833, C2 => n34, 
                           A => n1739, ZN => n1736);
   U1030 : AOI22_X1 port map( A1 => n31, A2 => REGISTERS_7_1_port, B1 => n28, 
                           B2 => REGISTERS_6_1_port, ZN => n1739);
   U1031 : OAI221_X1 port map( B1 => n2120, B2 => n85, C1 => n2088, C2 => n82, 
                           A => n1713, ZN => n1710);
   U1032 : AOI22_X1 port map( A1 => n79, A2 => REGISTERS_23_2_port, B1 => n76, 
                           B2 => REGISTERS_22_2_port, ZN => n1713);
   U1033 : OAI221_X1 port map( B1 => n1864, B2 => n37, C1 => n1832, C2 => n34, 
                           A => n1721, ZN => n1718);
   U1034 : AOI22_X1 port map( A1 => n31, A2 => REGISTERS_7_2_port, B1 => n28, 
                           B2 => REGISTERS_6_2_port, ZN => n1721);
   U1035 : OAI221_X1 port map( B1 => n2119, B2 => n85, C1 => n2087, C2 => n82, 
                           A => n1695, ZN => n1692);
   U1036 : AOI22_X1 port map( A1 => n79, A2 => REGISTERS_23_3_port, B1 => n76, 
                           B2 => REGISTERS_22_3_port, ZN => n1695);
   U1037 : OAI221_X1 port map( B1 => n1863, B2 => n37, C1 => n1831, C2 => n34, 
                           A => n1703, ZN => n1700);
   U1038 : AOI22_X1 port map( A1 => n31, A2 => REGISTERS_7_3_port, B1 => n28, 
                           B2 => REGISTERS_6_3_port, ZN => n1703);
   U1039 : OAI221_X1 port map( B1 => n2118, B2 => n85, C1 => n2086, C2 => n82, 
                           A => n1677, ZN => n1674);
   U1040 : AOI22_X1 port map( A1 => n79, A2 => REGISTERS_23_4_port, B1 => n76, 
                           B2 => REGISTERS_22_4_port, ZN => n1677);
   U1041 : OAI221_X1 port map( B1 => n1862, B2 => n37, C1 => n1830, C2 => n34, 
                           A => n1685, ZN => n1682);
   U1042 : AOI22_X1 port map( A1 => n31, A2 => REGISTERS_7_4_port, B1 => n28, 
                           B2 => REGISTERS_6_4_port, ZN => n1685);
   U1043 : OAI221_X1 port map( B1 => n2117, B2 => n85, C1 => n2085, C2 => n82, 
                           A => n1659, ZN => n1656);
   U1044 : AOI22_X1 port map( A1 => n79, A2 => REGISTERS_23_5_port, B1 => n76, 
                           B2 => REGISTERS_22_5_port, ZN => n1659);
   U1045 : OAI221_X1 port map( B1 => n1861, B2 => n37, C1 => n1829, C2 => n34, 
                           A => n1667, ZN => n1664);
   U1046 : AOI22_X1 port map( A1 => n31, A2 => REGISTERS_7_5_port, B1 => n28, 
                           B2 => REGISTERS_6_5_port, ZN => n1667);
   U1047 : OAI221_X1 port map( B1 => n2116, B2 => n85, C1 => n2084, C2 => n82, 
                           A => n1641, ZN => n1638);
   U1048 : AOI22_X1 port map( A1 => n79, A2 => REGISTERS_23_6_port, B1 => n76, 
                           B2 => REGISTERS_22_6_port, ZN => n1641);
   U1049 : OAI221_X1 port map( B1 => n1860, B2 => n37, C1 => n1828, C2 => n34, 
                           A => n1649, ZN => n1646);
   U1050 : AOI22_X1 port map( A1 => n31, A2 => REGISTERS_7_6_port, B1 => n28, 
                           B2 => REGISTERS_6_6_port, ZN => n1649);
   U1051 : OAI221_X1 port map( B1 => n2115, B2 => n85, C1 => n2083, C2 => n82, 
                           A => n1623, ZN => n1620);
   U1052 : AOI22_X1 port map( A1 => n79, A2 => REGISTERS_23_7_port, B1 => n76, 
                           B2 => REGISTERS_22_7_port, ZN => n1623);
   U1053 : OAI221_X1 port map( B1 => n1859, B2 => n37, C1 => n1827, C2 => n34, 
                           A => n1631, ZN => n1628);
   U1054 : AOI22_X1 port map( A1 => n31, A2 => REGISTERS_7_7_port, B1 => n28, 
                           B2 => REGISTERS_6_7_port, ZN => n1631);
   U1055 : OAI221_X1 port map( B1 => n2114, B2 => n85, C1 => n2082, C2 => n82, 
                           A => n1605, ZN => n1602);
   U1056 : AOI22_X1 port map( A1 => n79, A2 => REGISTERS_23_8_port, B1 => n76, 
                           B2 => REGISTERS_22_8_port, ZN => n1605);
   U1057 : OAI221_X1 port map( B1 => n1858, B2 => n37, C1 => n1826, C2 => n34, 
                           A => n1613, ZN => n1610);
   U1058 : AOI22_X1 port map( A1 => n31, A2 => REGISTERS_7_8_port, B1 => n28, 
                           B2 => REGISTERS_6_8_port, ZN => n1613);
   U1059 : OAI221_X1 port map( B1 => n2113, B2 => n85, C1 => n2081, C2 => n82, 
                           A => n1587, ZN => n1584);
   U1060 : AOI22_X1 port map( A1 => n79, A2 => REGISTERS_23_9_port, B1 => n76, 
                           B2 => REGISTERS_22_9_port, ZN => n1587);
   U1061 : OAI221_X1 port map( B1 => n1857, B2 => n37, C1 => n1825, C2 => n34, 
                           A => n1595, ZN => n1592);
   U1062 : AOI22_X1 port map( A1 => n31, A2 => REGISTERS_7_9_port, B1 => n28, 
                           B2 => REGISTERS_6_9_port, ZN => n1595);
   U1063 : OAI221_X1 port map( B1 => n2112, B2 => n85, C1 => n2080, C2 => n82, 
                           A => n1569, ZN => n1566);
   U1064 : AOI22_X1 port map( A1 => n79, A2 => REGISTERS_23_10_port, B1 => n76,
                           B2 => REGISTERS_22_10_port, ZN => n1569);
   U1065 : OAI221_X1 port map( B1 => n1856, B2 => n37, C1 => n1824, C2 => n34, 
                           A => n1577, ZN => n1574);
   U1066 : AOI22_X1 port map( A1 => n31, A2 => REGISTERS_7_10_port, B1 => n28, 
                           B2 => REGISTERS_6_10_port, ZN => n1577);
   U1067 : OAI221_X1 port map( B1 => n2100, B2 => n87, C1 => n2068, C2 => n84, 
                           A => n1353, ZN => n1350);
   U1068 : AOI22_X1 port map( A1 => n81, A2 => REGISTERS_23_22_port, B1 => n78,
                           B2 => REGISTERS_22_22_port, ZN => n1353);
   U1069 : OAI221_X1 port map( B1 => n1844, B2 => n39, C1 => n1812, C2 => n36, 
                           A => n1361, ZN => n1358);
   U1070 : AOI22_X1 port map( A1 => n33, A2 => REGISTERS_7_22_port, B1 => n30, 
                           B2 => REGISTERS_6_22_port, ZN => n1361);
   U1071 : OAI221_X1 port map( B1 => n2099, B2 => n87, C1 => n2067, C2 => n84, 
                           A => n1335, ZN => n1332);
   U1072 : AOI22_X1 port map( A1 => n81, A2 => REGISTERS_23_23_port, B1 => n78,
                           B2 => REGISTERS_22_23_port, ZN => n1335);
   U1073 : OAI221_X1 port map( B1 => n1843, B2 => n39, C1 => n1811, C2 => n36, 
                           A => n1343, ZN => n1340);
   U1074 : AOI22_X1 port map( A1 => n33, A2 => REGISTERS_7_23_port, B1 => n30, 
                           B2 => REGISTERS_6_23_port, ZN => n1343);
   U1075 : OAI221_X1 port map( B1 => n2098, B2 => n87, C1 => n2066, C2 => n84, 
                           A => n1317, ZN => n1314);
   U1076 : AOI22_X1 port map( A1 => n81, A2 => REGISTERS_23_24_port, B1 => n78,
                           B2 => REGISTERS_22_24_port, ZN => n1317);
   U1077 : OAI221_X1 port map( B1 => n1842, B2 => n39, C1 => n1810, C2 => n36, 
                           A => n1325, ZN => n1322);
   U1078 : AOI22_X1 port map( A1 => n33, A2 => REGISTERS_7_24_port, B1 => n30, 
                           B2 => REGISTERS_6_24_port, ZN => n1325);
   U1079 : OAI221_X1 port map( B1 => n2097, B2 => n87, C1 => n2065, C2 => n84, 
                           A => n1299, ZN => n1296);
   U1080 : AOI22_X1 port map( A1 => n81, A2 => REGISTERS_23_25_port, B1 => n78,
                           B2 => REGISTERS_22_25_port, ZN => n1299);
   U1081 : OAI221_X1 port map( B1 => n1841, B2 => n39, C1 => n1809, C2 => n36, 
                           A => n1307, ZN => n1304);
   U1082 : AOI22_X1 port map( A1 => n33, A2 => REGISTERS_7_25_port, B1 => n30, 
                           B2 => REGISTERS_6_25_port, ZN => n1307);
   U1083 : OAI221_X1 port map( B1 => n2096, B2 => n87, C1 => n2064, C2 => n84, 
                           A => n1281, ZN => n1278);
   U1084 : AOI22_X1 port map( A1 => n81, A2 => REGISTERS_23_26_port, B1 => n78,
                           B2 => REGISTERS_22_26_port, ZN => n1281);
   U1085 : OAI221_X1 port map( B1 => n1840, B2 => n39, C1 => n1808, C2 => n36, 
                           A => n1289, ZN => n1286);
   U1086 : AOI22_X1 port map( A1 => n33, A2 => REGISTERS_7_26_port, B1 => n30, 
                           B2 => REGISTERS_6_26_port, ZN => n1289);
   U1087 : OAI221_X1 port map( B1 => n2095, B2 => n87, C1 => n2063, C2 => n84, 
                           A => n1263, ZN => n1260);
   U1088 : AOI22_X1 port map( A1 => n81, A2 => REGISTERS_23_27_port, B1 => n78,
                           B2 => REGISTERS_22_27_port, ZN => n1263);
   U1089 : OAI221_X1 port map( B1 => n1839, B2 => n39, C1 => n1807, C2 => n36, 
                           A => n1271, ZN => n1268);
   U1090 : AOI22_X1 port map( A1 => n33, A2 => REGISTERS_7_27_port, B1 => n30, 
                           B2 => REGISTERS_6_27_port, ZN => n1271);
   U1091 : OAI221_X1 port map( B1 => n2094, B2 => n87, C1 => n2062, C2 => n84, 
                           A => n1245, ZN => n1242);
   U1092 : AOI22_X1 port map( A1 => n81, A2 => REGISTERS_23_28_port, B1 => n78,
                           B2 => REGISTERS_22_28_port, ZN => n1245);
   U1093 : OAI221_X1 port map( B1 => n1838, B2 => n39, C1 => n1806, C2 => n36, 
                           A => n1253, ZN => n1250);
   U1094 : AOI22_X1 port map( A1 => n33, A2 => REGISTERS_7_28_port, B1 => n30, 
                           B2 => REGISTERS_6_28_port, ZN => n1253);
   U1095 : OAI221_X1 port map( B1 => n2093, B2 => n87, C1 => n2061, C2 => n84, 
                           A => n1227, ZN => n1224);
   U1096 : AOI22_X1 port map( A1 => n81, A2 => REGISTERS_23_29_port, B1 => n78,
                           B2 => REGISTERS_22_29_port, ZN => n1227);
   U1097 : OAI221_X1 port map( B1 => n1837, B2 => n39, C1 => n1805, C2 => n36, 
                           A => n1235, ZN => n1232);
   U1098 : AOI22_X1 port map( A1 => n33, A2 => REGISTERS_7_29_port, B1 => n30, 
                           B2 => REGISTERS_6_29_port, ZN => n1235);
   U1099 : OAI221_X1 port map( B1 => n2092, B2 => n87, C1 => n2060, C2 => n84, 
                           A => n1209, ZN => n1206);
   U1100 : AOI22_X1 port map( A1 => n81, A2 => REGISTERS_23_30_port, B1 => n78,
                           B2 => REGISTERS_22_30_port, ZN => n1209);
   U1101 : OAI221_X1 port map( B1 => n1836, B2 => n39, C1 => n1804, C2 => n36, 
                           A => n1217, ZN => n1214);
   U1102 : AOI22_X1 port map( A1 => n33, A2 => REGISTERS_7_30_port, B1 => n30, 
                           B2 => REGISTERS_6_30_port, ZN => n1217);
   U1103 : OAI221_X1 port map( B1 => n2091, B2 => n87, C1 => n2059, C2 => n84, 
                           A => n1165, ZN => n1156);
   U1104 : AOI22_X1 port map( A1 => n81, A2 => REGISTERS_23_31_port, B1 => n78,
                           B2 => REGISTERS_22_31_port, ZN => n1165);
   U1105 : OAI221_X1 port map( B1 => n1835, B2 => n39, C1 => n1803, C2 => n36, 
                           A => n1189, ZN => n1180);
   U1106 : AOI22_X1 port map( A1 => n33, A2 => REGISTERS_7_31_port, B1 => n30, 
                           B2 => REGISTERS_6_31_port, ZN => n1189);
   U1107 : OAI221_X1 port map( B1 => n181, B2 => n2122, C1 => n178, C2 => n2090
                           , A => n1128, ZN => n1121);
   U1108 : AOI22_X1 port map( A1 => REGISTERS_23_0_port, A2 => n175, B1 => 
                           REGISTERS_22_0_port, B2 => n172, ZN => n1128);
   U1109 : OAI221_X1 port map( B1 => n133, B2 => n1866, C1 => n130, C2 => n1834
                           , A => n1144, ZN => n1139);
   U1110 : AOI22_X1 port map( A1 => REGISTERS_7_0_port, A2 => n127, B1 => 
                           REGISTERS_6_0_port, B2 => n124, ZN => n1144);
   U1111 : OAI221_X1 port map( B1 => n181, B2 => n2121, C1 => n178, C2 => n2089
                           , A => n1106, ZN => n1103);
   U1112 : AOI22_X1 port map( A1 => REGISTERS_23_1_port, A2 => n175, B1 => 
                           REGISTERS_22_1_port, B2 => n172, ZN => n1106);
   U1113 : OAI221_X1 port map( B1 => n133, B2 => n1865, C1 => n130, C2 => n1833
                           , A => n1114, ZN => n1111);
   U1114 : AOI22_X1 port map( A1 => REGISTERS_7_1_port, A2 => n127, B1 => 
                           REGISTERS_6_1_port, B2 => n124, ZN => n1114);
   U1115 : OAI221_X1 port map( B1 => n181, B2 => n2120, C1 => n178, C2 => n2088
                           , A => n1088, ZN => n1085);
   U1116 : AOI22_X1 port map( A1 => REGISTERS_23_2_port, A2 => n175, B1 => 
                           REGISTERS_22_2_port, B2 => n172, ZN => n1088);
   U1117 : OAI221_X1 port map( B1 => n133, B2 => n1864, C1 => n130, C2 => n1832
                           , A => n1096, ZN => n1093);
   U1118 : AOI22_X1 port map( A1 => REGISTERS_7_2_port, A2 => n127, B1 => 
                           REGISTERS_6_2_port, B2 => n124, ZN => n1096);
   U1119 : OAI221_X1 port map( B1 => n181, B2 => n2119, C1 => n178, C2 => n2087
                           , A => n1070, ZN => n1067);
   U1120 : AOI22_X1 port map( A1 => REGISTERS_23_3_port, A2 => n175, B1 => 
                           REGISTERS_22_3_port, B2 => n172, ZN => n1070);
   U1121 : OAI221_X1 port map( B1 => n133, B2 => n1863, C1 => n130, C2 => n1831
                           , A => n1078, ZN => n1075);
   U1122 : AOI22_X1 port map( A1 => REGISTERS_7_3_port, A2 => n127, B1 => 
                           REGISTERS_6_3_port, B2 => n124, ZN => n1078);
   U1123 : OAI221_X1 port map( B1 => n181, B2 => n2118, C1 => n178, C2 => n2086
                           , A => n1052, ZN => n1049);
   U1124 : AOI22_X1 port map( A1 => REGISTERS_23_4_port, A2 => n175, B1 => 
                           REGISTERS_22_4_port, B2 => n172, ZN => n1052);
   U1125 : OAI221_X1 port map( B1 => n133, B2 => n1862, C1 => n130, C2 => n1830
                           , A => n1060, ZN => n1057);
   U1126 : AOI22_X1 port map( A1 => REGISTERS_7_4_port, A2 => n127, B1 => 
                           REGISTERS_6_4_port, B2 => n124, ZN => n1060);
   U1127 : OAI221_X1 port map( B1 => n181, B2 => n2117, C1 => n178, C2 => n2085
                           , A => n1034, ZN => n1031);
   U1128 : AOI22_X1 port map( A1 => REGISTERS_23_5_port, A2 => n175, B1 => 
                           REGISTERS_22_5_port, B2 => n172, ZN => n1034);
   U1129 : OAI221_X1 port map( B1 => n133, B2 => n1861, C1 => n130, C2 => n1829
                           , A => n1042, ZN => n1039);
   U1130 : AOI22_X1 port map( A1 => REGISTERS_7_5_port, A2 => n127, B1 => 
                           REGISTERS_6_5_port, B2 => n124, ZN => n1042);
   U1131 : OAI221_X1 port map( B1 => n181, B2 => n2116, C1 => n178, C2 => n2084
                           , A => n1016, ZN => n1013);
   U1132 : AOI22_X1 port map( A1 => REGISTERS_23_6_port, A2 => n175, B1 => 
                           REGISTERS_22_6_port, B2 => n172, ZN => n1016);
   U1133 : OAI221_X1 port map( B1 => n133, B2 => n1860, C1 => n130, C2 => n1828
                           , A => n1024, ZN => n1021);
   U1134 : AOI22_X1 port map( A1 => REGISTERS_7_6_port, A2 => n127, B1 => 
                           REGISTERS_6_6_port, B2 => n124, ZN => n1024);
   U1135 : OAI221_X1 port map( B1 => n181, B2 => n2115, C1 => n178, C2 => n2083
                           , A => n998, ZN => n995);
   U1136 : AOI22_X1 port map( A1 => REGISTERS_23_7_port, A2 => n175, B1 => 
                           REGISTERS_22_7_port, B2 => n172, ZN => n998);
   U1137 : OAI221_X1 port map( B1 => n133, B2 => n1859, C1 => n130, C2 => n1827
                           , A => n1006, ZN => n1003);
   U1138 : AOI22_X1 port map( A1 => REGISTERS_7_7_port, A2 => n127, B1 => 
                           REGISTERS_6_7_port, B2 => n124, ZN => n1006);
   U1139 : OAI221_X1 port map( B1 => n181, B2 => n2114, C1 => n178, C2 => n2082
                           , A => n980, ZN => n977);
   U1140 : AOI22_X1 port map( A1 => REGISTERS_23_8_port, A2 => n175, B1 => 
                           REGISTERS_22_8_port, B2 => n172, ZN => n980);
   U1141 : OAI221_X1 port map( B1 => n133, B2 => n1858, C1 => n130, C2 => n1826
                           , A => n988, ZN => n985);
   U1142 : AOI22_X1 port map( A1 => REGISTERS_7_8_port, A2 => n127, B1 => 
                           REGISTERS_6_8_port, B2 => n124, ZN => n988);
   U1143 : OAI221_X1 port map( B1 => n181, B2 => n2113, C1 => n178, C2 => n2081
                           , A => n962, ZN => n959);
   U1144 : AOI22_X1 port map( A1 => REGISTERS_23_9_port, A2 => n175, B1 => 
                           REGISTERS_22_9_port, B2 => n172, ZN => n962);
   U1145 : OAI221_X1 port map( B1 => n133, B2 => n1857, C1 => n130, C2 => n1825
                           , A => n970, ZN => n967);
   U1146 : AOI22_X1 port map( A1 => REGISTERS_7_9_port, A2 => n127, B1 => 
                           REGISTERS_6_9_port, B2 => n124, ZN => n970);
   U1147 : OAI221_X1 port map( B1 => n181, B2 => n2112, C1 => n178, C2 => n2080
                           , A => n944, ZN => n941);
   U1148 : AOI22_X1 port map( A1 => REGISTERS_23_10_port, A2 => n175, B1 => 
                           REGISTERS_22_10_port, B2 => n172, ZN => n944);
   U1149 : OAI221_X1 port map( B1 => n133, B2 => n1856, C1 => n130, C2 => n1824
                           , A => n952, ZN => n949);
   U1150 : AOI22_X1 port map( A1 => REGISTERS_7_10_port, A2 => n127, B1 => 
                           REGISTERS_6_10_port, B2 => n124, ZN => n952);
   U1151 : OAI221_X1 port map( B1 => n181, B2 => n2111, C1 => n179, C2 => n2079
                           , A => n926, ZN => n923);
   U1152 : AOI22_X1 port map( A1 => REGISTERS_23_11_port, A2 => n175, B1 => 
                           REGISTERS_22_11_port, B2 => n172, ZN => n926);
   U1153 : OAI221_X1 port map( B1 => n133, B2 => n1855, C1 => n131, C2 => n1823
                           , A => n934, ZN => n931);
   U1154 : AOI22_X1 port map( A1 => REGISTERS_7_11_port, A2 => n127, B1 => 
                           REGISTERS_6_11_port, B2 => n124, ZN => n934);
   U1155 : OAI221_X1 port map( B1 => n182, B2 => n2110, C1 => n179, C2 => n2078
                           , A => n908, ZN => n905);
   U1156 : AOI22_X1 port map( A1 => REGISTERS_23_12_port, A2 => n176, B1 => 
                           REGISTERS_22_12_port, B2 => n173, ZN => n908);
   U1157 : OAI221_X1 port map( B1 => n134, B2 => n1854, C1 => n131, C2 => n1822
                           , A => n916, ZN => n913);
   U1158 : AOI22_X1 port map( A1 => REGISTERS_7_12_port, A2 => n128, B1 => 
                           REGISTERS_6_12_port, B2 => n125, ZN => n916);
   U1159 : OAI221_X1 port map( B1 => n182, B2 => n2109, C1 => n179, C2 => n2077
                           , A => n890, ZN => n887);
   U1160 : AOI22_X1 port map( A1 => REGISTERS_23_13_port, A2 => n176, B1 => 
                           REGISTERS_22_13_port, B2 => n173, ZN => n890);
   U1161 : OAI221_X1 port map( B1 => n134, B2 => n1853, C1 => n131, C2 => n1821
                           , A => n898, ZN => n895);
   U1162 : AOI22_X1 port map( A1 => REGISTERS_7_13_port, A2 => n128, B1 => 
                           REGISTERS_6_13_port, B2 => n125, ZN => n898);
   U1163 : OAI221_X1 port map( B1 => n182, B2 => n2108, C1 => n179, C2 => n2076
                           , A => n872, ZN => n869);
   U1164 : AOI22_X1 port map( A1 => REGISTERS_23_14_port, A2 => n176, B1 => 
                           REGISTERS_22_14_port, B2 => n173, ZN => n872);
   U1165 : OAI221_X1 port map( B1 => n134, B2 => n1852, C1 => n131, C2 => n1820
                           , A => n880, ZN => n877);
   U1166 : AOI22_X1 port map( A1 => REGISTERS_7_14_port, A2 => n128, B1 => 
                           REGISTERS_6_14_port, B2 => n125, ZN => n880);
   U1167 : OAI221_X1 port map( B1 => n182, B2 => n2107, C1 => n179, C2 => n2075
                           , A => n854, ZN => n851);
   U1168 : AOI22_X1 port map( A1 => REGISTERS_23_15_port, A2 => n176, B1 => 
                           REGISTERS_22_15_port, B2 => n173, ZN => n854);
   U1169 : OAI221_X1 port map( B1 => n134, B2 => n1851, C1 => n131, C2 => n1819
                           , A => n862, ZN => n859);
   U1170 : AOI22_X1 port map( A1 => REGISTERS_7_15_port, A2 => n128, B1 => 
                           REGISTERS_6_15_port, B2 => n125, ZN => n862);
   U1171 : OAI221_X1 port map( B1 => n182, B2 => n2106, C1 => n179, C2 => n2074
                           , A => n836, ZN => n833);
   U1172 : AOI22_X1 port map( A1 => REGISTERS_23_16_port, A2 => n176, B1 => 
                           REGISTERS_22_16_port, B2 => n173, ZN => n836);
   U1173 : OAI221_X1 port map( B1 => n134, B2 => n1850, C1 => n131, C2 => n1818
                           , A => n844, ZN => n841);
   U1174 : AOI22_X1 port map( A1 => REGISTERS_7_16_port, A2 => n128, B1 => 
                           REGISTERS_6_16_port, B2 => n125, ZN => n844);
   U1175 : OAI221_X1 port map( B1 => n182, B2 => n2105, C1 => n179, C2 => n2073
                           , A => n818, ZN => n815);
   U1176 : AOI22_X1 port map( A1 => REGISTERS_23_17_port, A2 => n176, B1 => 
                           REGISTERS_22_17_port, B2 => n173, ZN => n818);
   U1177 : OAI221_X1 port map( B1 => n134, B2 => n1849, C1 => n131, C2 => n1817
                           , A => n826, ZN => n823);
   U1178 : AOI22_X1 port map( A1 => REGISTERS_7_17_port, A2 => n128, B1 => 
                           REGISTERS_6_17_port, B2 => n125, ZN => n826);
   U1179 : OAI221_X1 port map( B1 => n182, B2 => n2104, C1 => n179, C2 => n2072
                           , A => n800, ZN => n797);
   U1180 : AOI22_X1 port map( A1 => REGISTERS_23_18_port, A2 => n176, B1 => 
                           REGISTERS_22_18_port, B2 => n173, ZN => n800);
   U1181 : OAI221_X1 port map( B1 => n134, B2 => n1848, C1 => n131, C2 => n1816
                           , A => n808, ZN => n805);
   U1182 : AOI22_X1 port map( A1 => REGISTERS_7_18_port, A2 => n128, B1 => 
                           REGISTERS_6_18_port, B2 => n125, ZN => n808);
   U1183 : OAI221_X1 port map( B1 => n182, B2 => n2103, C1 => n179, C2 => n2071
                           , A => n782, ZN => n779);
   U1184 : AOI22_X1 port map( A1 => REGISTERS_23_19_port, A2 => n176, B1 => 
                           REGISTERS_22_19_port, B2 => n173, ZN => n782);
   U1185 : OAI221_X1 port map( B1 => n134, B2 => n1847, C1 => n131, C2 => n1815
                           , A => n790, ZN => n787);
   U1186 : AOI22_X1 port map( A1 => REGISTERS_7_19_port, A2 => n128, B1 => 
                           REGISTERS_6_19_port, B2 => n125, ZN => n790);
   U1187 : OAI221_X1 port map( B1 => n182, B2 => n2102, C1 => n179, C2 => n2070
                           , A => n764, ZN => n761);
   U1188 : AOI22_X1 port map( A1 => REGISTERS_23_20_port, A2 => n176, B1 => 
                           REGISTERS_22_20_port, B2 => n173, ZN => n764);
   U1189 : OAI221_X1 port map( B1 => n134, B2 => n1846, C1 => n131, C2 => n1814
                           , A => n772, ZN => n769);
   U1190 : AOI22_X1 port map( A1 => REGISTERS_7_20_port, A2 => n128, B1 => 
                           REGISTERS_6_20_port, B2 => n125, ZN => n772);
   U1191 : OAI221_X1 port map( B1 => n182, B2 => n2101, C1 => n179, C2 => n2069
                           , A => n746, ZN => n743);
   U1192 : AOI22_X1 port map( A1 => REGISTERS_23_21_port, A2 => n176, B1 => 
                           REGISTERS_22_21_port, B2 => n173, ZN => n746);
   U1193 : OAI221_X1 port map( B1 => n134, B2 => n1845, C1 => n131, C2 => n1813
                           , A => n754, ZN => n751);
   U1194 : AOI22_X1 port map( A1 => REGISTERS_7_21_port, A2 => n128, B1 => 
                           REGISTERS_6_21_port, B2 => n125, ZN => n754);
   U1195 : OAI221_X1 port map( B1 => n182, B2 => n2100, C1 => n180, C2 => n2068
                           , A => n728, ZN => n725);
   U1196 : AOI22_X1 port map( A1 => REGISTERS_23_22_port, A2 => n176, B1 => 
                           REGISTERS_22_22_port, B2 => n173, ZN => n728);
   U1197 : OAI221_X1 port map( B1 => n134, B2 => n1844, C1 => n132, C2 => n1812
                           , A => n736, ZN => n733);
   U1198 : AOI22_X1 port map( A1 => REGISTERS_7_22_port, A2 => n128, B1 => 
                           REGISTERS_6_22_port, B2 => n125, ZN => n736);
   U1199 : OAI221_X1 port map( B1 => n182, B2 => n2099, C1 => n180, C2 => n2067
                           , A => n710, ZN => n707);
   U1200 : AOI22_X1 port map( A1 => REGISTERS_23_23_port, A2 => n176, B1 => 
                           REGISTERS_22_23_port, B2 => n173, ZN => n710);
   U1201 : OAI221_X1 port map( B1 => n134, B2 => n1843, C1 => n132, C2 => n1811
                           , A => n718, ZN => n715);
   U1202 : AOI22_X1 port map( A1 => REGISTERS_7_23_port, A2 => n128, B1 => 
                           REGISTERS_6_23_port, B2 => n125, ZN => n718);
   U1203 : OAI221_X1 port map( B1 => n2111, B2 => n86, C1 => n2079, C2 => n83, 
                           A => n1551, ZN => n1548);
   U1204 : AOI22_X1 port map( A1 => n80, A2 => REGISTERS_23_11_port, B1 => n77,
                           B2 => REGISTERS_22_11_port, ZN => n1551);
   U1205 : OAI221_X1 port map( B1 => n1855, B2 => n38, C1 => n1823, C2 => n35, 
                           A => n1559, ZN => n1556);
   U1206 : AOI22_X1 port map( A1 => n32, A2 => REGISTERS_7_11_port, B1 => n29, 
                           B2 => REGISTERS_6_11_port, ZN => n1559);
   U1207 : OAI221_X1 port map( B1 => n2110, B2 => n86, C1 => n2078, C2 => n83, 
                           A => n1533, ZN => n1530);
   U1208 : AOI22_X1 port map( A1 => n80, A2 => REGISTERS_23_12_port, B1 => n77,
                           B2 => REGISTERS_22_12_port, ZN => n1533);
   U1209 : OAI221_X1 port map( B1 => n1854, B2 => n38, C1 => n1822, C2 => n35, 
                           A => n1541, ZN => n1538);
   U1210 : AOI22_X1 port map( A1 => n32, A2 => REGISTERS_7_12_port, B1 => n29, 
                           B2 => REGISTERS_6_12_port, ZN => n1541);
   U1211 : OAI221_X1 port map( B1 => n2109, B2 => n86, C1 => n2077, C2 => n83, 
                           A => n1515, ZN => n1512);
   U1212 : AOI22_X1 port map( A1 => n80, A2 => REGISTERS_23_13_port, B1 => n77,
                           B2 => REGISTERS_22_13_port, ZN => n1515);
   U1213 : OAI221_X1 port map( B1 => n1853, B2 => n38, C1 => n1821, C2 => n35, 
                           A => n1523, ZN => n1520);
   U1214 : AOI22_X1 port map( A1 => n32, A2 => REGISTERS_7_13_port, B1 => n29, 
                           B2 => REGISTERS_6_13_port, ZN => n1523);
   U1215 : OAI221_X1 port map( B1 => n2108, B2 => n86, C1 => n2076, C2 => n83, 
                           A => n1497, ZN => n1494);
   U1216 : AOI22_X1 port map( A1 => n80, A2 => REGISTERS_23_14_port, B1 => n77,
                           B2 => REGISTERS_22_14_port, ZN => n1497);
   U1217 : OAI221_X1 port map( B1 => n1852, B2 => n38, C1 => n1820, C2 => n35, 
                           A => n1505, ZN => n1502);
   U1218 : AOI22_X1 port map( A1 => n32, A2 => REGISTERS_7_14_port, B1 => n29, 
                           B2 => REGISTERS_6_14_port, ZN => n1505);
   U1219 : OAI221_X1 port map( B1 => n2107, B2 => n86, C1 => n2075, C2 => n83, 
                           A => n1479, ZN => n1476);
   U1220 : AOI22_X1 port map( A1 => n80, A2 => REGISTERS_23_15_port, B1 => n77,
                           B2 => REGISTERS_22_15_port, ZN => n1479);
   U1221 : OAI221_X1 port map( B1 => n1851, B2 => n38, C1 => n1819, C2 => n35, 
                           A => n1487, ZN => n1484);
   U1222 : AOI22_X1 port map( A1 => n32, A2 => REGISTERS_7_15_port, B1 => n29, 
                           B2 => REGISTERS_6_15_port, ZN => n1487);
   U1223 : OAI221_X1 port map( B1 => n2106, B2 => n86, C1 => n2074, C2 => n83, 
                           A => n1461, ZN => n1458);
   U1224 : AOI22_X1 port map( A1 => n80, A2 => REGISTERS_23_16_port, B1 => n77,
                           B2 => REGISTERS_22_16_port, ZN => n1461);
   U1225 : OAI221_X1 port map( B1 => n1850, B2 => n38, C1 => n1818, C2 => n35, 
                           A => n1469, ZN => n1466);
   U1226 : AOI22_X1 port map( A1 => n32, A2 => REGISTERS_7_16_port, B1 => n29, 
                           B2 => REGISTERS_6_16_port, ZN => n1469);
   U1227 : OAI221_X1 port map( B1 => n2105, B2 => n86, C1 => n2073, C2 => n83, 
                           A => n1443, ZN => n1440);
   U1228 : AOI22_X1 port map( A1 => n80, A2 => REGISTERS_23_17_port, B1 => n77,
                           B2 => REGISTERS_22_17_port, ZN => n1443);
   U1229 : OAI221_X1 port map( B1 => n1849, B2 => n38, C1 => n1817, C2 => n35, 
                           A => n1451, ZN => n1448);
   U1230 : AOI22_X1 port map( A1 => n32, A2 => REGISTERS_7_17_port, B1 => n29, 
                           B2 => REGISTERS_6_17_port, ZN => n1451);
   U1231 : OAI221_X1 port map( B1 => n2104, B2 => n86, C1 => n2072, C2 => n83, 
                           A => n1425, ZN => n1422);
   U1232 : AOI22_X1 port map( A1 => n80, A2 => REGISTERS_23_18_port, B1 => n77,
                           B2 => REGISTERS_22_18_port, ZN => n1425);
   U1233 : OAI221_X1 port map( B1 => n1848, B2 => n38, C1 => n1816, C2 => n35, 
                           A => n1433, ZN => n1430);
   U1234 : AOI22_X1 port map( A1 => n32, A2 => REGISTERS_7_18_port, B1 => n29, 
                           B2 => REGISTERS_6_18_port, ZN => n1433);
   U1235 : OAI221_X1 port map( B1 => n2103, B2 => n86, C1 => n2071, C2 => n83, 
                           A => n1407, ZN => n1404);
   U1236 : AOI22_X1 port map( A1 => n80, A2 => REGISTERS_23_19_port, B1 => n77,
                           B2 => REGISTERS_22_19_port, ZN => n1407);
   U1237 : OAI221_X1 port map( B1 => n1847, B2 => n38, C1 => n1815, C2 => n35, 
                           A => n1415, ZN => n1412);
   U1238 : AOI22_X1 port map( A1 => n32, A2 => REGISTERS_7_19_port, B1 => n29, 
                           B2 => REGISTERS_6_19_port, ZN => n1415);
   U1239 : OAI221_X1 port map( B1 => n2102, B2 => n86, C1 => n2070, C2 => n83, 
                           A => n1389, ZN => n1386);
   U1240 : AOI22_X1 port map( A1 => n80, A2 => REGISTERS_23_20_port, B1 => n77,
                           B2 => REGISTERS_22_20_port, ZN => n1389);
   U1241 : OAI221_X1 port map( B1 => n1846, B2 => n38, C1 => n1814, C2 => n35, 
                           A => n1397, ZN => n1394);
   U1242 : AOI22_X1 port map( A1 => n32, A2 => REGISTERS_7_20_port, B1 => n29, 
                           B2 => REGISTERS_6_20_port, ZN => n1397);
   U1243 : OAI221_X1 port map( B1 => n2101, B2 => n86, C1 => n2069, C2 => n83, 
                           A => n1371, ZN => n1368);
   U1244 : AOI22_X1 port map( A1 => n80, A2 => REGISTERS_23_21_port, B1 => n77,
                           B2 => REGISTERS_22_21_port, ZN => n1371);
   U1245 : OAI221_X1 port map( B1 => n1845, B2 => n38, C1 => n1813, C2 => n35, 
                           A => n1379, ZN => n1376);
   U1246 : AOI22_X1 port map( A1 => n32, A2 => REGISTERS_7_21_port, B1 => n29, 
                           B2 => REGISTERS_6_21_port, ZN => n1379);
   U1247 : OAI221_X1 port map( B1 => n171, B2 => n2162, C1 => n168, C2 => n2130
                           , A => n693, ZN => n688);
   U1248 : AOI22_X1 port map( A1 => REGISTERS_27_24_port, A2 => n165, B1 => 
                           REGISTERS_26_24_port, B2 => n162, ZN => n693);
   U1249 : OAI221_X1 port map( B1 => n171, B2 => n2161, C1 => n168, C2 => n2129
                           , A => n675, ZN => n670);
   U1250 : AOI22_X1 port map( A1 => REGISTERS_27_25_port, A2 => n165, B1 => 
                           REGISTERS_26_25_port, B2 => n162, ZN => n675);
   U1251 : OAI221_X1 port map( B1 => n171, B2 => n2160, C1 => n168, C2 => n2128
                           , A => n657, ZN => n652);
   U1252 : AOI22_X1 port map( A1 => REGISTERS_27_26_port, A2 => n165, B1 => 
                           REGISTERS_26_26_port, B2 => n162, ZN => n657);
   U1253 : OAI221_X1 port map( B1 => n171, B2 => n2159, C1 => n168, C2 => n2127
                           , A => n639, ZN => n634);
   U1254 : AOI22_X1 port map( A1 => REGISTERS_27_27_port, A2 => n165, B1 => 
                           REGISTERS_26_27_port, B2 => n162, ZN => n639);
   U1255 : OAI221_X1 port map( B1 => n171, B2 => n2158, C1 => n168, C2 => n2126
                           , A => n621, ZN => n616);
   U1256 : AOI22_X1 port map( A1 => REGISTERS_27_28_port, A2 => n165, B1 => 
                           REGISTERS_26_28_port, B2 => n162, ZN => n621);
   U1257 : OAI221_X1 port map( B1 => n171, B2 => n2157, C1 => n168, C2 => n2125
                           , A => n603, ZN => n598);
   U1258 : AOI22_X1 port map( A1 => REGISTERS_27_29_port, A2 => n165, B1 => 
                           REGISTERS_26_29_port, B2 => n162, ZN => n603);
   U1259 : OAI221_X1 port map( B1 => n171, B2 => n2156, C1 => n168, C2 => n2124
                           , A => n585, ZN => n580);
   U1260 : AOI22_X1 port map( A1 => REGISTERS_27_30_port, A2 => n165, B1 => 
                           REGISTERS_26_30_port, B2 => n162, ZN => n585);
   U1261 : OAI221_X1 port map( B1 => n171, B2 => n2155, C1 => n168, C2 => n2123
                           , A => n545, ZN => n530);
   U1262 : AOI22_X1 port map( A1 => REGISTERS_27_31_port, A2 => n165, B1 => 
                           REGISTERS_26_31_port, B2 => n162, ZN => n545);
   U1263 : OAI221_X1 port map( B1 => n123, B2 => n1906, C1 => n120, C2 => n1874
                           , A => n701, ZN => n696);
   U1264 : AOI22_X1 port map( A1 => REGISTERS_11_24_port, A2 => n117, B1 => 
                           REGISTERS_10_24_port, B2 => n114, ZN => n701);
   U1265 : OAI221_X1 port map( B1 => n123, B2 => n1905, C1 => n120, C2 => n1873
                           , A => n683, ZN => n678);
   U1266 : AOI22_X1 port map( A1 => REGISTERS_11_25_port, A2 => n117, B1 => 
                           REGISTERS_10_25_port, B2 => n114, ZN => n683);
   U1267 : OAI221_X1 port map( B1 => n123, B2 => n1904, C1 => n120, C2 => n1872
                           , A => n665, ZN => n660);
   U1268 : AOI22_X1 port map( A1 => REGISTERS_11_26_port, A2 => n117, B1 => 
                           REGISTERS_10_26_port, B2 => n114, ZN => n665);
   U1269 : OAI221_X1 port map( B1 => n123, B2 => n1903, C1 => n120, C2 => n1871
                           , A => n647, ZN => n642);
   U1270 : AOI22_X1 port map( A1 => REGISTERS_11_27_port, A2 => n117, B1 => 
                           REGISTERS_10_27_port, B2 => n114, ZN => n647);
   U1271 : OAI221_X1 port map( B1 => n123, B2 => n1902, C1 => n120, C2 => n1870
                           , A => n629, ZN => n624);
   U1272 : AOI22_X1 port map( A1 => REGISTERS_11_28_port, A2 => n117, B1 => 
                           REGISTERS_10_28_port, B2 => n114, ZN => n629);
   U1273 : OAI221_X1 port map( B1 => n123, B2 => n1901, C1 => n120, C2 => n1869
                           , A => n611, ZN => n606);
   U1274 : AOI22_X1 port map( A1 => REGISTERS_11_29_port, A2 => n117, B1 => 
                           REGISTERS_10_29_port, B2 => n114, ZN => n611);
   U1275 : OAI221_X1 port map( B1 => n123, B2 => n1900, C1 => n120, C2 => n1868
                           , A => n593, ZN => n588);
   U1276 : AOI22_X1 port map( A1 => REGISTERS_11_30_port, A2 => n117, B1 => 
                           REGISTERS_10_30_port, B2 => n114, ZN => n593);
   U1277 : OAI221_X1 port map( B1 => n123, B2 => n1899, C1 => n120, C2 => n1867
                           , A => n569, ZN => n554);
   U1278 : AOI22_X1 port map( A1 => REGISTERS_11_31_port, A2 => n117, B1 => 
                           REGISTERS_10_31_port, B2 => n114, ZN => n569);
   U1279 : OAI221_X1 port map( B1 => n2186, B2 => n73, C1 => n2154, C2 => n70, 
                           A => n1757, ZN => n1745);
   U1280 : AOI22_X1 port map( A1 => n67, A2 => REGISTERS_27_0_port, B1 => n64, 
                           B2 => REGISTERS_26_0_port, ZN => n1757);
   U1281 : OAI221_X1 port map( B1 => n1930, B2 => n25, C1 => n1898, C2 => n22, 
                           A => n1771, ZN => n1763);
   U1282 : AOI22_X1 port map( A1 => n19, A2 => REGISTERS_11_0_port, B1 => n16, 
                           B2 => REGISTERS_10_0_port, ZN => n1771);
   U1283 : OAI221_X1 port map( B1 => n2185, B2 => n73, C1 => n2153, C2 => n70, 
                           A => n1732, ZN => n1727);
   U1284 : AOI22_X1 port map( A1 => n67, A2 => REGISTERS_27_1_port, B1 => n64, 
                           B2 => REGISTERS_26_1_port, ZN => n1732);
   U1285 : OAI221_X1 port map( B1 => n1929, B2 => n25, C1 => n1897, C2 => n22, 
                           A => n1740, ZN => n1735);
   U1286 : AOI22_X1 port map( A1 => n19, A2 => REGISTERS_11_1_port, B1 => n16, 
                           B2 => REGISTERS_10_1_port, ZN => n1740);
   U1287 : OAI221_X1 port map( B1 => n2184, B2 => n73, C1 => n2152, C2 => n70, 
                           A => n1714, ZN => n1709);
   U1288 : AOI22_X1 port map( A1 => n67, A2 => REGISTERS_27_2_port, B1 => n64, 
                           B2 => REGISTERS_26_2_port, ZN => n1714);
   U1289 : OAI221_X1 port map( B1 => n1928, B2 => n25, C1 => n1896, C2 => n22, 
                           A => n1722, ZN => n1717);
   U1290 : AOI22_X1 port map( A1 => n19, A2 => REGISTERS_11_2_port, B1 => n16, 
                           B2 => REGISTERS_10_2_port, ZN => n1722);
   U1291 : OAI221_X1 port map( B1 => n2183, B2 => n73, C1 => n2151, C2 => n70, 
                           A => n1696, ZN => n1691);
   U1292 : AOI22_X1 port map( A1 => n67, A2 => REGISTERS_27_3_port, B1 => n64, 
                           B2 => REGISTERS_26_3_port, ZN => n1696);
   U1293 : OAI221_X1 port map( B1 => n1927, B2 => n25, C1 => n1895, C2 => n22, 
                           A => n1704, ZN => n1699);
   U1294 : AOI22_X1 port map( A1 => n19, A2 => REGISTERS_11_3_port, B1 => n16, 
                           B2 => REGISTERS_10_3_port, ZN => n1704);
   U1295 : OAI221_X1 port map( B1 => n2182, B2 => n73, C1 => n2150, C2 => n70, 
                           A => n1678, ZN => n1673);
   U1296 : AOI22_X1 port map( A1 => n67, A2 => REGISTERS_27_4_port, B1 => n64, 
                           B2 => REGISTERS_26_4_port, ZN => n1678);
   U1297 : OAI221_X1 port map( B1 => n1926, B2 => n25, C1 => n1894, C2 => n22, 
                           A => n1686, ZN => n1681);
   U1298 : AOI22_X1 port map( A1 => n19, A2 => REGISTERS_11_4_port, B1 => n16, 
                           B2 => REGISTERS_10_4_port, ZN => n1686);
   U1299 : OAI221_X1 port map( B1 => n2181, B2 => n73, C1 => n2149, C2 => n70, 
                           A => n1660, ZN => n1655);
   U1300 : AOI22_X1 port map( A1 => n67, A2 => REGISTERS_27_5_port, B1 => n64, 
                           B2 => REGISTERS_26_5_port, ZN => n1660);
   U1301 : OAI221_X1 port map( B1 => n1925, B2 => n25, C1 => n1893, C2 => n22, 
                           A => n1668, ZN => n1663);
   U1302 : AOI22_X1 port map( A1 => n19, A2 => REGISTERS_11_5_port, B1 => n16, 
                           B2 => REGISTERS_10_5_port, ZN => n1668);
   U1303 : OAI221_X1 port map( B1 => n2180, B2 => n73, C1 => n2148, C2 => n70, 
                           A => n1642, ZN => n1637);
   U1304 : AOI22_X1 port map( A1 => n67, A2 => REGISTERS_27_6_port, B1 => n64, 
                           B2 => REGISTERS_26_6_port, ZN => n1642);
   U1305 : OAI221_X1 port map( B1 => n1924, B2 => n25, C1 => n1892, C2 => n22, 
                           A => n1650, ZN => n1645);
   U1306 : AOI22_X1 port map( A1 => n19, A2 => REGISTERS_11_6_port, B1 => n16, 
                           B2 => REGISTERS_10_6_port, ZN => n1650);
   U1307 : OAI221_X1 port map( B1 => n2179, B2 => n73, C1 => n2147, C2 => n70, 
                           A => n1624, ZN => n1619);
   U1308 : AOI22_X1 port map( A1 => n67, A2 => REGISTERS_27_7_port, B1 => n64, 
                           B2 => REGISTERS_26_7_port, ZN => n1624);
   U1309 : OAI221_X1 port map( B1 => n1923, B2 => n25, C1 => n1891, C2 => n22, 
                           A => n1632, ZN => n1627);
   U1310 : AOI22_X1 port map( A1 => n19, A2 => REGISTERS_11_7_port, B1 => n16, 
                           B2 => REGISTERS_10_7_port, ZN => n1632);
   U1311 : OAI221_X1 port map( B1 => n2178, B2 => n73, C1 => n2146, C2 => n70, 
                           A => n1606, ZN => n1601);
   U1312 : AOI22_X1 port map( A1 => n67, A2 => REGISTERS_27_8_port, B1 => n64, 
                           B2 => REGISTERS_26_8_port, ZN => n1606);
   U1313 : OAI221_X1 port map( B1 => n1922, B2 => n25, C1 => n1890, C2 => n22, 
                           A => n1614, ZN => n1609);
   U1314 : AOI22_X1 port map( A1 => n19, A2 => REGISTERS_11_8_port, B1 => n16, 
                           B2 => REGISTERS_10_8_port, ZN => n1614);
   U1315 : OAI221_X1 port map( B1 => n2177, B2 => n73, C1 => n2145, C2 => n70, 
                           A => n1588, ZN => n1583);
   U1316 : AOI22_X1 port map( A1 => n67, A2 => REGISTERS_27_9_port, B1 => n64, 
                           B2 => REGISTERS_26_9_port, ZN => n1588);
   U1317 : OAI221_X1 port map( B1 => n1921, B2 => n25, C1 => n1889, C2 => n22, 
                           A => n1596, ZN => n1591);
   U1318 : AOI22_X1 port map( A1 => n19, A2 => REGISTERS_11_9_port, B1 => n16, 
                           B2 => REGISTERS_10_9_port, ZN => n1596);
   U1319 : OAI221_X1 port map( B1 => n2176, B2 => n73, C1 => n2144, C2 => n70, 
                           A => n1570, ZN => n1565);
   U1320 : AOI22_X1 port map( A1 => n67, A2 => REGISTERS_27_10_port, B1 => n64,
                           B2 => REGISTERS_26_10_port, ZN => n1570);
   U1321 : OAI221_X1 port map( B1 => n1920, B2 => n25, C1 => n1888, C2 => n22, 
                           A => n1578, ZN => n1573);
   U1322 : AOI22_X1 port map( A1 => n19, A2 => REGISTERS_11_10_port, B1 => n16,
                           B2 => REGISTERS_10_10_port, ZN => n1578);
   U1323 : OAI221_X1 port map( B1 => n159, B2 => n2226, C1 => n156, C2 => n2194
                           , A => n694, ZN => n687);
   U1324 : AOI22_X1 port map( A1 => REGISTERS_29_24_port, A2 => n153, B1 => 
                           REGISTERS_28_24_port, B2 => n150, ZN => n694);
   U1325 : OAI221_X1 port map( B1 => n159, B2 => n2225, C1 => n156, C2 => n2193
                           , A => n676, ZN => n669);
   U1326 : AOI22_X1 port map( A1 => REGISTERS_29_25_port, A2 => n153, B1 => 
                           REGISTERS_28_25_port, B2 => n150, ZN => n676);
   U1327 : OAI221_X1 port map( B1 => n159, B2 => n2224, C1 => n156, C2 => n2192
                           , A => n658, ZN => n651);
   U1328 : AOI22_X1 port map( A1 => REGISTERS_29_26_port, A2 => n153, B1 => 
                           REGISTERS_28_26_port, B2 => n150, ZN => n658);
   U1329 : OAI221_X1 port map( B1 => n159, B2 => n2223, C1 => n156, C2 => n2191
                           , A => n640, ZN => n633);
   U1330 : AOI22_X1 port map( A1 => REGISTERS_29_27_port, A2 => n153, B1 => 
                           REGISTERS_28_27_port, B2 => n150, ZN => n640);
   U1331 : OAI221_X1 port map( B1 => n159, B2 => n2222, C1 => n156, C2 => n2190
                           , A => n622, ZN => n615);
   U1332 : AOI22_X1 port map( A1 => REGISTERS_29_28_port, A2 => n153, B1 => 
                           REGISTERS_28_28_port, B2 => n150, ZN => n622);
   U1333 : OAI221_X1 port map( B1 => n159, B2 => n2221, C1 => n156, C2 => n2189
                           , A => n604, ZN => n597);
   U1334 : AOI22_X1 port map( A1 => REGISTERS_29_29_port, A2 => n153, B1 => 
                           REGISTERS_28_29_port, B2 => n150, ZN => n604);
   U1335 : OAI221_X1 port map( B1 => n159, B2 => n2220, C1 => n156, C2 => n2188
                           , A => n586, ZN => n579);
   U1336 : AOI22_X1 port map( A1 => REGISTERS_29_30_port, A2 => n153, B1 => 
                           REGISTERS_28_30_port, B2 => n150, ZN => n586);
   U1337 : OAI221_X1 port map( B1 => n159, B2 => n2219, C1 => n156, C2 => n2187
                           , A => n550, ZN => n529);
   U1338 : AOI22_X1 port map( A1 => REGISTERS_29_31_port, A2 => n153, B1 => 
                           REGISTERS_28_31_port, B2 => n150, ZN => n550);
   U1339 : OAI221_X1 port map( B1 => n2164, B2 => n75, C1 => n2132, C2 => n72, 
                           A => n1354, ZN => n1349);
   U1340 : AOI22_X1 port map( A1 => n69, A2 => REGISTERS_27_22_port, B1 => n66,
                           B2 => REGISTERS_26_22_port, ZN => n1354);
   U1341 : OAI221_X1 port map( B1 => n1908, B2 => n27, C1 => n1876, C2 => n24, 
                           A => n1362, ZN => n1357);
   U1342 : AOI22_X1 port map( A1 => n21, A2 => REGISTERS_11_22_port, B1 => n18,
                           B2 => REGISTERS_10_22_port, ZN => n1362);
   U1343 : OAI221_X1 port map( B1 => n2163, B2 => n75, C1 => n2131, C2 => n72, 
                           A => n1336, ZN => n1331);
   U1344 : AOI22_X1 port map( A1 => n69, A2 => REGISTERS_27_23_port, B1 => n66,
                           B2 => REGISTERS_26_23_port, ZN => n1336);
   U1345 : OAI221_X1 port map( B1 => n1907, B2 => n27, C1 => n1875, C2 => n24, 
                           A => n1344, ZN => n1339);
   U1346 : AOI22_X1 port map( A1 => n21, A2 => REGISTERS_11_23_port, B1 => n18,
                           B2 => REGISTERS_10_23_port, ZN => n1344);
   U1347 : OAI221_X1 port map( B1 => n2162, B2 => n75, C1 => n2130, C2 => n72, 
                           A => n1318, ZN => n1313);
   U1348 : AOI22_X1 port map( A1 => n69, A2 => REGISTERS_27_24_port, B1 => n66,
                           B2 => REGISTERS_26_24_port, ZN => n1318);
   U1349 : OAI221_X1 port map( B1 => n1906, B2 => n27, C1 => n1874, C2 => n24, 
                           A => n1326, ZN => n1321);
   U1350 : AOI22_X1 port map( A1 => n21, A2 => REGISTERS_11_24_port, B1 => n18,
                           B2 => REGISTERS_10_24_port, ZN => n1326);
   U1351 : OAI221_X1 port map( B1 => n2161, B2 => n75, C1 => n2129, C2 => n72, 
                           A => n1300, ZN => n1295);
   U1352 : AOI22_X1 port map( A1 => n69, A2 => REGISTERS_27_25_port, B1 => n66,
                           B2 => REGISTERS_26_25_port, ZN => n1300);
   U1353 : OAI221_X1 port map( B1 => n1905, B2 => n27, C1 => n1873, C2 => n24, 
                           A => n1308, ZN => n1303);
   U1354 : AOI22_X1 port map( A1 => n21, A2 => REGISTERS_11_25_port, B1 => n18,
                           B2 => REGISTERS_10_25_port, ZN => n1308);
   U1355 : OAI221_X1 port map( B1 => n2160, B2 => n75, C1 => n2128, C2 => n72, 
                           A => n1282, ZN => n1277);
   U1356 : AOI22_X1 port map( A1 => n69, A2 => REGISTERS_27_26_port, B1 => n66,
                           B2 => REGISTERS_26_26_port, ZN => n1282);
   U1357 : OAI221_X1 port map( B1 => n1904, B2 => n27, C1 => n1872, C2 => n24, 
                           A => n1290, ZN => n1285);
   U1358 : AOI22_X1 port map( A1 => n21, A2 => REGISTERS_11_26_port, B1 => n18,
                           B2 => REGISTERS_10_26_port, ZN => n1290);
   U1359 : OAI221_X1 port map( B1 => n2159, B2 => n75, C1 => n2127, C2 => n72, 
                           A => n1264, ZN => n1259);
   U1360 : AOI22_X1 port map( A1 => n69, A2 => REGISTERS_27_27_port, B1 => n66,
                           B2 => REGISTERS_26_27_port, ZN => n1264);
   U1361 : OAI221_X1 port map( B1 => n1903, B2 => n27, C1 => n1871, C2 => n24, 
                           A => n1272, ZN => n1267);
   U1362 : AOI22_X1 port map( A1 => n21, A2 => REGISTERS_11_27_port, B1 => n18,
                           B2 => REGISTERS_10_27_port, ZN => n1272);
   U1363 : OAI221_X1 port map( B1 => n2158, B2 => n75, C1 => n2126, C2 => n72, 
                           A => n1246, ZN => n1241);
   U1364 : AOI22_X1 port map( A1 => n69, A2 => REGISTERS_27_28_port, B1 => n66,
                           B2 => REGISTERS_26_28_port, ZN => n1246);
   U1365 : OAI221_X1 port map( B1 => n1902, B2 => n27, C1 => n1870, C2 => n24, 
                           A => n1254, ZN => n1249);
   U1366 : AOI22_X1 port map( A1 => n21, A2 => REGISTERS_11_28_port, B1 => n18,
                           B2 => REGISTERS_10_28_port, ZN => n1254);
   U1367 : OAI221_X1 port map( B1 => n2157, B2 => n75, C1 => n2125, C2 => n72, 
                           A => n1228, ZN => n1223);
   U1368 : AOI22_X1 port map( A1 => n69, A2 => REGISTERS_27_29_port, B1 => n66,
                           B2 => REGISTERS_26_29_port, ZN => n1228);
   U1369 : OAI221_X1 port map( B1 => n1901, B2 => n27, C1 => n1869, C2 => n24, 
                           A => n1236, ZN => n1231);
   U1370 : AOI22_X1 port map( A1 => n21, A2 => REGISTERS_11_29_port, B1 => n18,
                           B2 => REGISTERS_10_29_port, ZN => n1236);
   U1371 : OAI221_X1 port map( B1 => n2156, B2 => n75, C1 => n2124, C2 => n72, 
                           A => n1210, ZN => n1205);
   U1372 : AOI22_X1 port map( A1 => n69, A2 => REGISTERS_27_30_port, B1 => n66,
                           B2 => REGISTERS_26_30_port, ZN => n1210);
   U1373 : OAI221_X1 port map( B1 => n1900, B2 => n27, C1 => n1868, C2 => n24, 
                           A => n1218, ZN => n1213);
   U1374 : AOI22_X1 port map( A1 => n21, A2 => REGISTERS_11_30_port, B1 => n18,
                           B2 => REGISTERS_10_30_port, ZN => n1218);
   U1375 : OAI221_X1 port map( B1 => n2155, B2 => n75, C1 => n2123, C2 => n72, 
                           A => n1170, ZN => n1155);
   U1376 : AOI22_X1 port map( A1 => n69, A2 => REGISTERS_27_31_port, B1 => n66,
                           B2 => REGISTERS_26_31_port, ZN => n1170);
   U1377 : OAI221_X1 port map( B1 => n1899, B2 => n27, C1 => n1867, C2 => n24, 
                           A => n1194, ZN => n1179);
   U1378 : AOI22_X1 port map( A1 => n21, A2 => REGISTERS_11_31_port, B1 => n18,
                           B2 => REGISTERS_10_31_port, ZN => n1194);
   U1379 : OAI221_X1 port map( B1 => n2250, B2 => n61, C1 => n2218, C2 => n58, 
                           A => n1760, ZN => n1744);
   U1380 : AOI22_X1 port map( A1 => n55, A2 => REGISTERS_29_0_port, B1 => n52, 
                           B2 => REGISTERS_28_0_port, ZN => n1760);
   U1381 : OAI221_X1 port map( B1 => n2249, B2 => n61, C1 => n2217, C2 => n58, 
                           A => n1733, ZN => n1726);
   U1382 : AOI22_X1 port map( A1 => n55, A2 => REGISTERS_29_1_port, B1 => n52, 
                           B2 => REGISTERS_28_1_port, ZN => n1733);
   U1383 : OAI221_X1 port map( B1 => n2248, B2 => n61, C1 => n2216, C2 => n58, 
                           A => n1715, ZN => n1708);
   U1384 : AOI22_X1 port map( A1 => n55, A2 => REGISTERS_29_2_port, B1 => n52, 
                           B2 => REGISTERS_28_2_port, ZN => n1715);
   U1385 : OAI221_X1 port map( B1 => n2247, B2 => n61, C1 => n2215, C2 => n58, 
                           A => n1697, ZN => n1690);
   U1386 : AOI22_X1 port map( A1 => n55, A2 => REGISTERS_29_3_port, B1 => n52, 
                           B2 => REGISTERS_28_3_port, ZN => n1697);
   U1387 : OAI221_X1 port map( B1 => n2246, B2 => n61, C1 => n2214, C2 => n58, 
                           A => n1679, ZN => n1672);
   U1388 : AOI22_X1 port map( A1 => n55, A2 => REGISTERS_29_4_port, B1 => n52, 
                           B2 => REGISTERS_28_4_port, ZN => n1679);
   U1389 : OAI221_X1 port map( B1 => n2245, B2 => n61, C1 => n2213, C2 => n58, 
                           A => n1661, ZN => n1654);
   U1390 : AOI22_X1 port map( A1 => n55, A2 => REGISTERS_29_5_port, B1 => n52, 
                           B2 => REGISTERS_28_5_port, ZN => n1661);
   U1391 : OAI221_X1 port map( B1 => n2244, B2 => n61, C1 => n2212, C2 => n58, 
                           A => n1643, ZN => n1636);
   U1392 : AOI22_X1 port map( A1 => n55, A2 => REGISTERS_29_6_port, B1 => n52, 
                           B2 => REGISTERS_28_6_port, ZN => n1643);
   U1393 : OAI221_X1 port map( B1 => n2243, B2 => n61, C1 => n2211, C2 => n58, 
                           A => n1625, ZN => n1618);
   U1394 : AOI22_X1 port map( A1 => n55, A2 => REGISTERS_29_7_port, B1 => n52, 
                           B2 => REGISTERS_28_7_port, ZN => n1625);
   U1395 : OAI221_X1 port map( B1 => n2242, B2 => n61, C1 => n2210, C2 => n58, 
                           A => n1607, ZN => n1600);
   U1396 : AOI22_X1 port map( A1 => n55, A2 => REGISTERS_29_8_port, B1 => n52, 
                           B2 => REGISTERS_28_8_port, ZN => n1607);
   U1397 : OAI221_X1 port map( B1 => n2241, B2 => n61, C1 => n2209, C2 => n58, 
                           A => n1589, ZN => n1582);
   U1398 : AOI22_X1 port map( A1 => n55, A2 => REGISTERS_29_9_port, B1 => n52, 
                           B2 => REGISTERS_28_9_port, ZN => n1589);
   U1399 : OAI221_X1 port map( B1 => n2240, B2 => n61, C1 => n2208, C2 => n58, 
                           A => n1571, ZN => n1564);
   U1400 : AOI22_X1 port map( A1 => n55, A2 => REGISTERS_29_10_port, B1 => n52,
                           B2 => REGISTERS_28_10_port, ZN => n1571);
   U1401 : OAI221_X1 port map( B1 => n2228, B2 => n63, C1 => n2196, C2 => n60, 
                           A => n1355, ZN => n1348);
   U1402 : AOI22_X1 port map( A1 => n57, A2 => REGISTERS_29_22_port, B1 => n54,
                           B2 => REGISTERS_28_22_port, ZN => n1355);
   U1403 : OAI221_X1 port map( B1 => n2227, B2 => n63, C1 => n2195, C2 => n60, 
                           A => n1337, ZN => n1330);
   U1404 : AOI22_X1 port map( A1 => n57, A2 => REGISTERS_29_23_port, B1 => n54,
                           B2 => REGISTERS_28_23_port, ZN => n1337);
   U1405 : OAI221_X1 port map( B1 => n2226, B2 => n63, C1 => n2194, C2 => n60, 
                           A => n1319, ZN => n1312);
   U1406 : AOI22_X1 port map( A1 => n57, A2 => REGISTERS_29_24_port, B1 => n54,
                           B2 => REGISTERS_28_24_port, ZN => n1319);
   U1407 : OAI221_X1 port map( B1 => n2225, B2 => n63, C1 => n2193, C2 => n60, 
                           A => n1301, ZN => n1294);
   U1408 : AOI22_X1 port map( A1 => n57, A2 => REGISTERS_29_25_port, B1 => n54,
                           B2 => REGISTERS_28_25_port, ZN => n1301);
   U1409 : OAI221_X1 port map( B1 => n2224, B2 => n63, C1 => n2192, C2 => n60, 
                           A => n1283, ZN => n1276);
   U1410 : AOI22_X1 port map( A1 => n57, A2 => REGISTERS_29_26_port, B1 => n54,
                           B2 => REGISTERS_28_26_port, ZN => n1283);
   U1411 : OAI221_X1 port map( B1 => n2223, B2 => n63, C1 => n2191, C2 => n60, 
                           A => n1265, ZN => n1258);
   U1412 : AOI22_X1 port map( A1 => n57, A2 => REGISTERS_29_27_port, B1 => n54,
                           B2 => REGISTERS_28_27_port, ZN => n1265);
   U1413 : OAI221_X1 port map( B1 => n2222, B2 => n63, C1 => n2190, C2 => n60, 
                           A => n1247, ZN => n1240);
   U1414 : AOI22_X1 port map( A1 => n57, A2 => REGISTERS_29_28_port, B1 => n54,
                           B2 => REGISTERS_28_28_port, ZN => n1247);
   U1415 : OAI221_X1 port map( B1 => n2221, B2 => n63, C1 => n2189, C2 => n60, 
                           A => n1229, ZN => n1222);
   U1416 : AOI22_X1 port map( A1 => n57, A2 => REGISTERS_29_29_port, B1 => n54,
                           B2 => REGISTERS_28_29_port, ZN => n1229);
   U1417 : OAI221_X1 port map( B1 => n2220, B2 => n63, C1 => n2188, C2 => n60, 
                           A => n1211, ZN => n1204);
   U1418 : AOI22_X1 port map( A1 => n57, A2 => REGISTERS_29_30_port, B1 => n54,
                           B2 => REGISTERS_28_30_port, ZN => n1211);
   U1419 : OAI221_X1 port map( B1 => n2219, B2 => n63, C1 => n2187, C2 => n60, 
                           A => n1175, ZN => n1154);
   U1420 : AOI22_X1 port map( A1 => n57, A2 => REGISTERS_29_31_port, B1 => n54,
                           B2 => REGISTERS_28_31_port, ZN => n1175);
   U1421 : OAI221_X1 port map( B1 => n169, B2 => n2186, C1 => n166, C2 => n2154
                           , A => n1132, ZN => n1120);
   U1422 : AOI22_X1 port map( A1 => REGISTERS_27_0_port, A2 => n163, B1 => 
                           REGISTERS_26_0_port, B2 => n160, ZN => n1132);
   U1423 : OAI221_X1 port map( B1 => n121, B2 => n1930, C1 => n118, C2 => n1898
                           , A => n1146, ZN => n1138);
   U1424 : AOI22_X1 port map( A1 => REGISTERS_11_0_port, A2 => n115, B1 => 
                           REGISTERS_10_0_port, B2 => n112, ZN => n1146);
   U1425 : OAI221_X1 port map( B1 => n169, B2 => n2185, C1 => n166, C2 => n2153
                           , A => n1107, ZN => n1102);
   U1426 : AOI22_X1 port map( A1 => REGISTERS_27_1_port, A2 => n163, B1 => 
                           REGISTERS_26_1_port, B2 => n160, ZN => n1107);
   U1427 : OAI221_X1 port map( B1 => n121, B2 => n1929, C1 => n118, C2 => n1897
                           , A => n1115, ZN => n1110);
   U1428 : AOI22_X1 port map( A1 => REGISTERS_11_1_port, A2 => n115, B1 => 
                           REGISTERS_10_1_port, B2 => n112, ZN => n1115);
   U1429 : OAI221_X1 port map( B1 => n169, B2 => n2184, C1 => n166, C2 => n2152
                           , A => n1089, ZN => n1084);
   U1430 : AOI22_X1 port map( A1 => REGISTERS_27_2_port, A2 => n163, B1 => 
                           REGISTERS_26_2_port, B2 => n160, ZN => n1089);
   U1431 : OAI221_X1 port map( B1 => n121, B2 => n1928, C1 => n118, C2 => n1896
                           , A => n1097, ZN => n1092);
   U1432 : AOI22_X1 port map( A1 => REGISTERS_11_2_port, A2 => n115, B1 => 
                           REGISTERS_10_2_port, B2 => n112, ZN => n1097);
   U1433 : OAI221_X1 port map( B1 => n169, B2 => n2183, C1 => n166, C2 => n2151
                           , A => n1071, ZN => n1066);
   U1434 : AOI22_X1 port map( A1 => REGISTERS_27_3_port, A2 => n163, B1 => 
                           REGISTERS_26_3_port, B2 => n160, ZN => n1071);
   U1435 : OAI221_X1 port map( B1 => n121, B2 => n1927, C1 => n118, C2 => n1895
                           , A => n1079, ZN => n1074);
   U1436 : AOI22_X1 port map( A1 => REGISTERS_11_3_port, A2 => n115, B1 => 
                           REGISTERS_10_3_port, B2 => n112, ZN => n1079);
   U1437 : OAI221_X1 port map( B1 => n169, B2 => n2182, C1 => n166, C2 => n2150
                           , A => n1053, ZN => n1048);
   U1438 : AOI22_X1 port map( A1 => REGISTERS_27_4_port, A2 => n163, B1 => 
                           REGISTERS_26_4_port, B2 => n160, ZN => n1053);
   U1439 : OAI221_X1 port map( B1 => n121, B2 => n1926, C1 => n118, C2 => n1894
                           , A => n1061, ZN => n1056);
   U1440 : AOI22_X1 port map( A1 => REGISTERS_11_4_port, A2 => n115, B1 => 
                           REGISTERS_10_4_port, B2 => n112, ZN => n1061);
   U1441 : OAI221_X1 port map( B1 => n169, B2 => n2181, C1 => n166, C2 => n2149
                           , A => n1035, ZN => n1030);
   U1442 : AOI22_X1 port map( A1 => REGISTERS_27_5_port, A2 => n163, B1 => 
                           REGISTERS_26_5_port, B2 => n160, ZN => n1035);
   U1443 : OAI221_X1 port map( B1 => n121, B2 => n1925, C1 => n118, C2 => n1893
                           , A => n1043, ZN => n1038);
   U1444 : AOI22_X1 port map( A1 => REGISTERS_11_5_port, A2 => n115, B1 => 
                           REGISTERS_10_5_port, B2 => n112, ZN => n1043);
   U1445 : OAI221_X1 port map( B1 => n169, B2 => n2180, C1 => n166, C2 => n2148
                           , A => n1017, ZN => n1012);
   U1446 : AOI22_X1 port map( A1 => REGISTERS_27_6_port, A2 => n163, B1 => 
                           REGISTERS_26_6_port, B2 => n160, ZN => n1017);
   U1447 : OAI221_X1 port map( B1 => n121, B2 => n1924, C1 => n118, C2 => n1892
                           , A => n1025, ZN => n1020);
   U1448 : AOI22_X1 port map( A1 => REGISTERS_11_6_port, A2 => n115, B1 => 
                           REGISTERS_10_6_port, B2 => n112, ZN => n1025);
   U1449 : OAI221_X1 port map( B1 => n169, B2 => n2179, C1 => n166, C2 => n2147
                           , A => n999, ZN => n994);
   U1450 : AOI22_X1 port map( A1 => REGISTERS_27_7_port, A2 => n163, B1 => 
                           REGISTERS_26_7_port, B2 => n160, ZN => n999);
   U1451 : OAI221_X1 port map( B1 => n121, B2 => n1923, C1 => n118, C2 => n1891
                           , A => n1007, ZN => n1002);
   U1452 : AOI22_X1 port map( A1 => REGISTERS_11_7_port, A2 => n115, B1 => 
                           REGISTERS_10_7_port, B2 => n112, ZN => n1007);
   U1453 : OAI221_X1 port map( B1 => n169, B2 => n2178, C1 => n166, C2 => n2146
                           , A => n981, ZN => n976);
   U1454 : AOI22_X1 port map( A1 => REGISTERS_27_8_port, A2 => n163, B1 => 
                           REGISTERS_26_8_port, B2 => n160, ZN => n981);
   U1455 : OAI221_X1 port map( B1 => n121, B2 => n1922, C1 => n118, C2 => n1890
                           , A => n989, ZN => n984);
   U1456 : AOI22_X1 port map( A1 => REGISTERS_11_8_port, A2 => n115, B1 => 
                           REGISTERS_10_8_port, B2 => n112, ZN => n989);
   U1457 : OAI221_X1 port map( B1 => n169, B2 => n2177, C1 => n166, C2 => n2145
                           , A => n963, ZN => n958);
   U1458 : AOI22_X1 port map( A1 => REGISTERS_27_9_port, A2 => n163, B1 => 
                           REGISTERS_26_9_port, B2 => n160, ZN => n963);
   U1459 : OAI221_X1 port map( B1 => n121, B2 => n1921, C1 => n118, C2 => n1889
                           , A => n971, ZN => n966);
   U1460 : AOI22_X1 port map( A1 => REGISTERS_11_9_port, A2 => n115, B1 => 
                           REGISTERS_10_9_port, B2 => n112, ZN => n971);
   U1461 : OAI221_X1 port map( B1 => n169, B2 => n2176, C1 => n166, C2 => n2144
                           , A => n945, ZN => n940);
   U1462 : AOI22_X1 port map( A1 => REGISTERS_27_10_port, A2 => n163, B1 => 
                           REGISTERS_26_10_port, B2 => n160, ZN => n945);
   U1463 : OAI221_X1 port map( B1 => n121, B2 => n1920, C1 => n118, C2 => n1888
                           , A => n953, ZN => n948);
   U1464 : AOI22_X1 port map( A1 => REGISTERS_11_10_port, A2 => n115, B1 => 
                           REGISTERS_10_10_port, B2 => n112, ZN => n953);
   U1465 : OAI221_X1 port map( B1 => n169, B2 => n2175, C1 => n167, C2 => n2143
                           , A => n927, ZN => n922);
   U1466 : AOI22_X1 port map( A1 => REGISTERS_27_11_port, A2 => n163, B1 => 
                           REGISTERS_26_11_port, B2 => n160, ZN => n927);
   U1467 : OAI221_X1 port map( B1 => n121, B2 => n1919, C1 => n119, C2 => n1887
                           , A => n935, ZN => n930);
   U1468 : AOI22_X1 port map( A1 => REGISTERS_11_11_port, A2 => n115, B1 => 
                           REGISTERS_10_11_port, B2 => n112, ZN => n935);
   U1469 : OAI221_X1 port map( B1 => n170, B2 => n2174, C1 => n167, C2 => n2142
                           , A => n909, ZN => n904);
   U1470 : AOI22_X1 port map( A1 => REGISTERS_27_12_port, A2 => n164, B1 => 
                           REGISTERS_26_12_port, B2 => n161, ZN => n909);
   U1471 : OAI221_X1 port map( B1 => n122, B2 => n1918, C1 => n119, C2 => n1886
                           , A => n917, ZN => n912);
   U1472 : AOI22_X1 port map( A1 => REGISTERS_11_12_port, A2 => n116, B1 => 
                           REGISTERS_10_12_port, B2 => n113, ZN => n917);
   U1473 : OAI221_X1 port map( B1 => n170, B2 => n2173, C1 => n167, C2 => n2141
                           , A => n891, ZN => n886);
   U1474 : AOI22_X1 port map( A1 => REGISTERS_27_13_port, A2 => n164, B1 => 
                           REGISTERS_26_13_port, B2 => n161, ZN => n891);
   U1475 : OAI221_X1 port map( B1 => n122, B2 => n1917, C1 => n119, C2 => n1885
                           , A => n899, ZN => n894);
   U1476 : AOI22_X1 port map( A1 => REGISTERS_11_13_port, A2 => n116, B1 => 
                           REGISTERS_10_13_port, B2 => n113, ZN => n899);
   U1477 : OAI221_X1 port map( B1 => n170, B2 => n2172, C1 => n167, C2 => n2140
                           , A => n873, ZN => n868);
   U1478 : AOI22_X1 port map( A1 => REGISTERS_27_14_port, A2 => n164, B1 => 
                           REGISTERS_26_14_port, B2 => n161, ZN => n873);
   U1479 : OAI221_X1 port map( B1 => n122, B2 => n1916, C1 => n119, C2 => n1884
                           , A => n881, ZN => n876);
   U1480 : AOI22_X1 port map( A1 => REGISTERS_11_14_port, A2 => n116, B1 => 
                           REGISTERS_10_14_port, B2 => n113, ZN => n881);
   U1481 : OAI221_X1 port map( B1 => n170, B2 => n2171, C1 => n167, C2 => n2139
                           , A => n855, ZN => n850);
   U1482 : AOI22_X1 port map( A1 => REGISTERS_27_15_port, A2 => n164, B1 => 
                           REGISTERS_26_15_port, B2 => n161, ZN => n855);
   U1483 : OAI221_X1 port map( B1 => n122, B2 => n1915, C1 => n119, C2 => n1883
                           , A => n863, ZN => n858);
   U1484 : AOI22_X1 port map( A1 => REGISTERS_11_15_port, A2 => n116, B1 => 
                           REGISTERS_10_15_port, B2 => n113, ZN => n863);
   U1485 : OAI221_X1 port map( B1 => n170, B2 => n2170, C1 => n167, C2 => n2138
                           , A => n837, ZN => n832);
   U1486 : AOI22_X1 port map( A1 => REGISTERS_27_16_port, A2 => n164, B1 => 
                           REGISTERS_26_16_port, B2 => n161, ZN => n837);
   U1487 : OAI221_X1 port map( B1 => n122, B2 => n1914, C1 => n119, C2 => n1882
                           , A => n845, ZN => n840);
   U1488 : AOI22_X1 port map( A1 => REGISTERS_11_16_port, A2 => n116, B1 => 
                           REGISTERS_10_16_port, B2 => n113, ZN => n845);
   U1489 : OAI221_X1 port map( B1 => n170, B2 => n2169, C1 => n167, C2 => n2137
                           , A => n819, ZN => n814);
   U1490 : AOI22_X1 port map( A1 => REGISTERS_27_17_port, A2 => n164, B1 => 
                           REGISTERS_26_17_port, B2 => n161, ZN => n819);
   U1491 : OAI221_X1 port map( B1 => n122, B2 => n1913, C1 => n119, C2 => n1881
                           , A => n827, ZN => n822);
   U1492 : AOI22_X1 port map( A1 => REGISTERS_11_17_port, A2 => n116, B1 => 
                           REGISTERS_10_17_port, B2 => n113, ZN => n827);
   U1493 : OAI221_X1 port map( B1 => n170, B2 => n2168, C1 => n167, C2 => n2136
                           , A => n801, ZN => n796);
   U1494 : AOI22_X1 port map( A1 => REGISTERS_27_18_port, A2 => n164, B1 => 
                           REGISTERS_26_18_port, B2 => n161, ZN => n801);
   U1495 : OAI221_X1 port map( B1 => n122, B2 => n1912, C1 => n119, C2 => n1880
                           , A => n809, ZN => n804);
   U1496 : AOI22_X1 port map( A1 => REGISTERS_11_18_port, A2 => n116, B1 => 
                           REGISTERS_10_18_port, B2 => n113, ZN => n809);
   U1497 : OAI221_X1 port map( B1 => n170, B2 => n2167, C1 => n167, C2 => n2135
                           , A => n783, ZN => n778);
   U1498 : AOI22_X1 port map( A1 => REGISTERS_27_19_port, A2 => n164, B1 => 
                           REGISTERS_26_19_port, B2 => n161, ZN => n783);
   U1499 : OAI221_X1 port map( B1 => n122, B2 => n1911, C1 => n119, C2 => n1879
                           , A => n791, ZN => n786);
   U1500 : AOI22_X1 port map( A1 => REGISTERS_11_19_port, A2 => n116, B1 => 
                           REGISTERS_10_19_port, B2 => n113, ZN => n791);
   U1501 : OAI221_X1 port map( B1 => n170, B2 => n2166, C1 => n167, C2 => n2134
                           , A => n765, ZN => n760);
   U1502 : AOI22_X1 port map( A1 => REGISTERS_27_20_port, A2 => n164, B1 => 
                           REGISTERS_26_20_port, B2 => n161, ZN => n765);
   U1503 : OAI221_X1 port map( B1 => n122, B2 => n1910, C1 => n119, C2 => n1878
                           , A => n773, ZN => n768);
   U1504 : AOI22_X1 port map( A1 => REGISTERS_11_20_port, A2 => n116, B1 => 
                           REGISTERS_10_20_port, B2 => n113, ZN => n773);
   U1505 : OAI221_X1 port map( B1 => n170, B2 => n2165, C1 => n167, C2 => n2133
                           , A => n747, ZN => n742);
   U1506 : AOI22_X1 port map( A1 => REGISTERS_27_21_port, A2 => n164, B1 => 
                           REGISTERS_26_21_port, B2 => n161, ZN => n747);
   U1507 : OAI221_X1 port map( B1 => n122, B2 => n1909, C1 => n119, C2 => n1877
                           , A => n755, ZN => n750);
   U1508 : AOI22_X1 port map( A1 => REGISTERS_11_21_port, A2 => n116, B1 => 
                           REGISTERS_10_21_port, B2 => n113, ZN => n755);
   U1509 : OAI221_X1 port map( B1 => n170, B2 => n2164, C1 => n168, C2 => n2132
                           , A => n729, ZN => n724);
   U1510 : AOI22_X1 port map( A1 => REGISTERS_27_22_port, A2 => n164, B1 => 
                           REGISTERS_26_22_port, B2 => n161, ZN => n729);
   U1511 : OAI221_X1 port map( B1 => n122, B2 => n1908, C1 => n120, C2 => n1876
                           , A => n737, ZN => n732);
   U1512 : AOI22_X1 port map( A1 => REGISTERS_11_22_port, A2 => n116, B1 => 
                           REGISTERS_10_22_port, B2 => n113, ZN => n737);
   U1513 : OAI221_X1 port map( B1 => n170, B2 => n2163, C1 => n168, C2 => n2131
                           , A => n711, ZN => n706);
   U1514 : AOI22_X1 port map( A1 => REGISTERS_27_23_port, A2 => n164, B1 => 
                           REGISTERS_26_23_port, B2 => n161, ZN => n711);
   U1515 : OAI221_X1 port map( B1 => n122, B2 => n1907, C1 => n120, C2 => n1875
                           , A => n719, ZN => n714);
   U1516 : AOI22_X1 port map( A1 => REGISTERS_11_23_port, A2 => n116, B1 => 
                           REGISTERS_10_23_port, B2 => n113, ZN => n719);
   U1517 : OAI221_X1 port map( B1 => n2175, B2 => n74, C1 => n2143, C2 => n71, 
                           A => n1552, ZN => n1547);
   U1518 : AOI22_X1 port map( A1 => n68, A2 => REGISTERS_27_11_port, B1 => n65,
                           B2 => REGISTERS_26_11_port, ZN => n1552);
   U1519 : OAI221_X1 port map( B1 => n1919, B2 => n26, C1 => n1887, C2 => n23, 
                           A => n1560, ZN => n1555);
   U1520 : AOI22_X1 port map( A1 => n20, A2 => REGISTERS_11_11_port, B1 => n17,
                           B2 => REGISTERS_10_11_port, ZN => n1560);
   U1521 : OAI221_X1 port map( B1 => n2174, B2 => n74, C1 => n2142, C2 => n71, 
                           A => n1534, ZN => n1529);
   U1522 : AOI22_X1 port map( A1 => n68, A2 => REGISTERS_27_12_port, B1 => n65,
                           B2 => REGISTERS_26_12_port, ZN => n1534);
   U1523 : OAI221_X1 port map( B1 => n1918, B2 => n26, C1 => n1886, C2 => n23, 
                           A => n1542, ZN => n1537);
   U1524 : AOI22_X1 port map( A1 => n20, A2 => REGISTERS_11_12_port, B1 => n17,
                           B2 => REGISTERS_10_12_port, ZN => n1542);
   U1525 : OAI221_X1 port map( B1 => n2173, B2 => n74, C1 => n2141, C2 => n71, 
                           A => n1516, ZN => n1511);
   U1526 : AOI22_X1 port map( A1 => n68, A2 => REGISTERS_27_13_port, B1 => n65,
                           B2 => REGISTERS_26_13_port, ZN => n1516);
   U1527 : OAI221_X1 port map( B1 => n1917, B2 => n26, C1 => n1885, C2 => n23, 
                           A => n1524, ZN => n1519);
   U1528 : AOI22_X1 port map( A1 => n20, A2 => REGISTERS_11_13_port, B1 => n17,
                           B2 => REGISTERS_10_13_port, ZN => n1524);
   U1529 : OAI221_X1 port map( B1 => n2172, B2 => n74, C1 => n2140, C2 => n71, 
                           A => n1498, ZN => n1493);
   U1530 : AOI22_X1 port map( A1 => n68, A2 => REGISTERS_27_14_port, B1 => n65,
                           B2 => REGISTERS_26_14_port, ZN => n1498);
   U1531 : OAI221_X1 port map( B1 => n1916, B2 => n26, C1 => n1884, C2 => n23, 
                           A => n1506, ZN => n1501);
   U1532 : AOI22_X1 port map( A1 => n20, A2 => REGISTERS_11_14_port, B1 => n17,
                           B2 => REGISTERS_10_14_port, ZN => n1506);
   U1533 : OAI221_X1 port map( B1 => n2171, B2 => n74, C1 => n2139, C2 => n71, 
                           A => n1480, ZN => n1475);
   U1534 : AOI22_X1 port map( A1 => n68, A2 => REGISTERS_27_15_port, B1 => n65,
                           B2 => REGISTERS_26_15_port, ZN => n1480);
   U1535 : OAI221_X1 port map( B1 => n1915, B2 => n26, C1 => n1883, C2 => n23, 
                           A => n1488, ZN => n1483);
   U1536 : AOI22_X1 port map( A1 => n20, A2 => REGISTERS_11_15_port, B1 => n17,
                           B2 => REGISTERS_10_15_port, ZN => n1488);
   U1537 : OAI221_X1 port map( B1 => n2170, B2 => n74, C1 => n2138, C2 => n71, 
                           A => n1462, ZN => n1457);
   U1538 : AOI22_X1 port map( A1 => n68, A2 => REGISTERS_27_16_port, B1 => n65,
                           B2 => REGISTERS_26_16_port, ZN => n1462);
   U1539 : OAI221_X1 port map( B1 => n1914, B2 => n26, C1 => n1882, C2 => n23, 
                           A => n1470, ZN => n1465);
   U1540 : AOI22_X1 port map( A1 => n20, A2 => REGISTERS_11_16_port, B1 => n17,
                           B2 => REGISTERS_10_16_port, ZN => n1470);
   U1541 : OAI221_X1 port map( B1 => n2169, B2 => n74, C1 => n2137, C2 => n71, 
                           A => n1444, ZN => n1439);
   U1542 : AOI22_X1 port map( A1 => n68, A2 => REGISTERS_27_17_port, B1 => n65,
                           B2 => REGISTERS_26_17_port, ZN => n1444);
   U1543 : OAI221_X1 port map( B1 => n1913, B2 => n26, C1 => n1881, C2 => n23, 
                           A => n1452, ZN => n1447);
   U1544 : AOI22_X1 port map( A1 => n20, A2 => REGISTERS_11_17_port, B1 => n17,
                           B2 => REGISTERS_10_17_port, ZN => n1452);
   U1545 : OAI221_X1 port map( B1 => n2168, B2 => n74, C1 => n2136, C2 => n71, 
                           A => n1426, ZN => n1421);
   U1546 : AOI22_X1 port map( A1 => n68, A2 => REGISTERS_27_18_port, B1 => n65,
                           B2 => REGISTERS_26_18_port, ZN => n1426);
   U1547 : OAI221_X1 port map( B1 => n1912, B2 => n26, C1 => n1880, C2 => n23, 
                           A => n1434, ZN => n1429);
   U1548 : AOI22_X1 port map( A1 => n20, A2 => REGISTERS_11_18_port, B1 => n17,
                           B2 => REGISTERS_10_18_port, ZN => n1434);
   U1549 : OAI221_X1 port map( B1 => n2167, B2 => n74, C1 => n2135, C2 => n71, 
                           A => n1408, ZN => n1403);
   U1550 : AOI22_X1 port map( A1 => n68, A2 => REGISTERS_27_19_port, B1 => n65,
                           B2 => REGISTERS_26_19_port, ZN => n1408);
   U1551 : OAI221_X1 port map( B1 => n1911, B2 => n26, C1 => n1879, C2 => n23, 
                           A => n1416, ZN => n1411);
   U1552 : AOI22_X1 port map( A1 => n20, A2 => REGISTERS_11_19_port, B1 => n17,
                           B2 => REGISTERS_10_19_port, ZN => n1416);
   U1553 : OAI221_X1 port map( B1 => n2166, B2 => n74, C1 => n2134, C2 => n71, 
                           A => n1390, ZN => n1385);
   U1554 : AOI22_X1 port map( A1 => n68, A2 => REGISTERS_27_20_port, B1 => n65,
                           B2 => REGISTERS_26_20_port, ZN => n1390);
   U1555 : OAI221_X1 port map( B1 => n1910, B2 => n26, C1 => n1878, C2 => n23, 
                           A => n1398, ZN => n1393);
   U1556 : AOI22_X1 port map( A1 => n20, A2 => REGISTERS_11_20_port, B1 => n17,
                           B2 => REGISTERS_10_20_port, ZN => n1398);
   U1557 : OAI221_X1 port map( B1 => n2165, B2 => n74, C1 => n2133, C2 => n71, 
                           A => n1372, ZN => n1367);
   U1558 : AOI22_X1 port map( A1 => n68, A2 => REGISTERS_27_21_port, B1 => n65,
                           B2 => REGISTERS_26_21_port, ZN => n1372);
   U1559 : OAI221_X1 port map( B1 => n1909, B2 => n26, C1 => n1877, C2 => n23, 
                           A => n1380, ZN => n1375);
   U1560 : AOI22_X1 port map( A1 => n20, A2 => REGISTERS_11_21_port, B1 => n17,
                           B2 => REGISTERS_10_21_port, ZN => n1380);
   U1561 : OAI221_X1 port map( B1 => n157, B2 => n2250, C1 => n154, C2 => n2218
                           , A => n1135, ZN => n1119);
   U1562 : AOI22_X1 port map( A1 => REGISTERS_29_0_port, A2 => n151, B1 => 
                           REGISTERS_28_0_port, B2 => n148, ZN => n1135);
   U1563 : OAI221_X1 port map( B1 => n157, B2 => n2249, C1 => n154, C2 => n2217
                           , A => n1108, ZN => n1101);
   U1564 : AOI22_X1 port map( A1 => REGISTERS_29_1_port, A2 => n151, B1 => 
                           REGISTERS_28_1_port, B2 => n148, ZN => n1108);
   U1565 : OAI221_X1 port map( B1 => n157, B2 => n2248, C1 => n154, C2 => n2216
                           , A => n1090, ZN => n1083);
   U1566 : AOI22_X1 port map( A1 => REGISTERS_29_2_port, A2 => n151, B1 => 
                           REGISTERS_28_2_port, B2 => n148, ZN => n1090);
   U1567 : OAI221_X1 port map( B1 => n157, B2 => n2247, C1 => n154, C2 => n2215
                           , A => n1072, ZN => n1065);
   U1568 : AOI22_X1 port map( A1 => REGISTERS_29_3_port, A2 => n151, B1 => 
                           REGISTERS_28_3_port, B2 => n148, ZN => n1072);
   U1569 : OAI221_X1 port map( B1 => n157, B2 => n2246, C1 => n154, C2 => n2214
                           , A => n1054, ZN => n1047);
   U1570 : AOI22_X1 port map( A1 => REGISTERS_29_4_port, A2 => n151, B1 => 
                           REGISTERS_28_4_port, B2 => n148, ZN => n1054);
   U1571 : OAI221_X1 port map( B1 => n157, B2 => n2245, C1 => n154, C2 => n2213
                           , A => n1036, ZN => n1029);
   U1572 : AOI22_X1 port map( A1 => REGISTERS_29_5_port, A2 => n151, B1 => 
                           REGISTERS_28_5_port, B2 => n148, ZN => n1036);
   U1573 : OAI221_X1 port map( B1 => n157, B2 => n2244, C1 => n154, C2 => n2212
                           , A => n1018, ZN => n1011);
   U1574 : AOI22_X1 port map( A1 => REGISTERS_29_6_port, A2 => n151, B1 => 
                           REGISTERS_28_6_port, B2 => n148, ZN => n1018);
   U1575 : OAI221_X1 port map( B1 => n157, B2 => n2243, C1 => n154, C2 => n2211
                           , A => n1000, ZN => n993);
   U1576 : AOI22_X1 port map( A1 => REGISTERS_29_7_port, A2 => n151, B1 => 
                           REGISTERS_28_7_port, B2 => n148, ZN => n1000);
   U1577 : OAI221_X1 port map( B1 => n157, B2 => n2242, C1 => n154, C2 => n2210
                           , A => n982, ZN => n975);
   U1578 : AOI22_X1 port map( A1 => REGISTERS_29_8_port, A2 => n151, B1 => 
                           REGISTERS_28_8_port, B2 => n148, ZN => n982);
   U1579 : OAI221_X1 port map( B1 => n157, B2 => n2241, C1 => n154, C2 => n2209
                           , A => n964, ZN => n957);
   U1580 : AOI22_X1 port map( A1 => REGISTERS_29_9_port, A2 => n151, B1 => 
                           REGISTERS_28_9_port, B2 => n148, ZN => n964);
   U1581 : OAI221_X1 port map( B1 => n157, B2 => n2240, C1 => n154, C2 => n2208
                           , A => n946, ZN => n939);
   U1582 : AOI22_X1 port map( A1 => REGISTERS_29_10_port, A2 => n151, B1 => 
                           REGISTERS_28_10_port, B2 => n148, ZN => n946);
   U1583 : OAI221_X1 port map( B1 => n157, B2 => n2239, C1 => n155, C2 => n2207
                           , A => n928, ZN => n921);
   U1584 : AOI22_X1 port map( A1 => REGISTERS_29_11_port, A2 => n151, B1 => 
                           REGISTERS_28_11_port, B2 => n148, ZN => n928);
   U1585 : OAI221_X1 port map( B1 => n158, B2 => n2238, C1 => n155, C2 => n2206
                           , A => n910, ZN => n903);
   U1586 : AOI22_X1 port map( A1 => REGISTERS_29_12_port, A2 => n152, B1 => 
                           REGISTERS_28_12_port, B2 => n149, ZN => n910);
   U1587 : OAI221_X1 port map( B1 => n158, B2 => n2237, C1 => n155, C2 => n2205
                           , A => n892, ZN => n885);
   U1588 : AOI22_X1 port map( A1 => REGISTERS_29_13_port, A2 => n152, B1 => 
                           REGISTERS_28_13_port, B2 => n149, ZN => n892);
   U1589 : OAI221_X1 port map( B1 => n158, B2 => n2236, C1 => n155, C2 => n2204
                           , A => n874, ZN => n867);
   U1590 : AOI22_X1 port map( A1 => REGISTERS_29_14_port, A2 => n152, B1 => 
                           REGISTERS_28_14_port, B2 => n149, ZN => n874);
   U1591 : OAI221_X1 port map( B1 => n158, B2 => n2235, C1 => n155, C2 => n2203
                           , A => n856, ZN => n849);
   U1592 : AOI22_X1 port map( A1 => REGISTERS_29_15_port, A2 => n152, B1 => 
                           REGISTERS_28_15_port, B2 => n149, ZN => n856);
   U1593 : OAI221_X1 port map( B1 => n158, B2 => n2234, C1 => n155, C2 => n2202
                           , A => n838, ZN => n831);
   U1594 : AOI22_X1 port map( A1 => REGISTERS_29_16_port, A2 => n152, B1 => 
                           REGISTERS_28_16_port, B2 => n149, ZN => n838);
   U1595 : OAI221_X1 port map( B1 => n158, B2 => n2233, C1 => n155, C2 => n2201
                           , A => n820, ZN => n813);
   U1596 : AOI22_X1 port map( A1 => REGISTERS_29_17_port, A2 => n152, B1 => 
                           REGISTERS_28_17_port, B2 => n149, ZN => n820);
   U1597 : OAI221_X1 port map( B1 => n158, B2 => n2232, C1 => n155, C2 => n2200
                           , A => n802, ZN => n795);
   U1598 : AOI22_X1 port map( A1 => REGISTERS_29_18_port, A2 => n152, B1 => 
                           REGISTERS_28_18_port, B2 => n149, ZN => n802);
   U1599 : OAI221_X1 port map( B1 => n158, B2 => n2231, C1 => n155, C2 => n2199
                           , A => n784, ZN => n777);
   U1600 : AOI22_X1 port map( A1 => REGISTERS_29_19_port, A2 => n152, B1 => 
                           REGISTERS_28_19_port, B2 => n149, ZN => n784);
   U1601 : OAI221_X1 port map( B1 => n158, B2 => n2230, C1 => n155, C2 => n2198
                           , A => n766, ZN => n759);
   U1602 : AOI22_X1 port map( A1 => REGISTERS_29_20_port, A2 => n152, B1 => 
                           REGISTERS_28_20_port, B2 => n149, ZN => n766);
   U1603 : OAI221_X1 port map( B1 => n158, B2 => n2229, C1 => n155, C2 => n2197
                           , A => n748, ZN => n741);
   U1604 : AOI22_X1 port map( A1 => REGISTERS_29_21_port, A2 => n152, B1 => 
                           REGISTERS_28_21_port, B2 => n149, ZN => n748);
   U1605 : OAI221_X1 port map( B1 => n158, B2 => n2228, C1 => n156, C2 => n2196
                           , A => n730, ZN => n723);
   U1606 : AOI22_X1 port map( A1 => REGISTERS_29_22_port, A2 => n152, B1 => 
                           REGISTERS_28_22_port, B2 => n149, ZN => n730);
   U1607 : OAI221_X1 port map( B1 => n158, B2 => n2227, C1 => n156, C2 => n2195
                           , A => n712, ZN => n705);
   U1608 : AOI22_X1 port map( A1 => REGISTERS_29_23_port, A2 => n152, B1 => 
                           REGISTERS_28_23_port, B2 => n149, ZN => n712);
   U1609 : OAI221_X1 port map( B1 => n2239, B2 => n62, C1 => n2207, C2 => n59, 
                           A => n1553, ZN => n1546);
   U1610 : AOI22_X1 port map( A1 => n56, A2 => REGISTERS_29_11_port, B1 => n53,
                           B2 => REGISTERS_28_11_port, ZN => n1553);
   U1611 : OAI221_X1 port map( B1 => n2238, B2 => n62, C1 => n2206, C2 => n59, 
                           A => n1535, ZN => n1528);
   U1612 : AOI22_X1 port map( A1 => n56, A2 => REGISTERS_29_12_port, B1 => n53,
                           B2 => REGISTERS_28_12_port, ZN => n1535);
   U1613 : OAI221_X1 port map( B1 => n2237, B2 => n62, C1 => n2205, C2 => n59, 
                           A => n1517, ZN => n1510);
   U1614 : AOI22_X1 port map( A1 => n56, A2 => REGISTERS_29_13_port, B1 => n53,
                           B2 => REGISTERS_28_13_port, ZN => n1517);
   U1615 : OAI221_X1 port map( B1 => n2236, B2 => n62, C1 => n2204, C2 => n59, 
                           A => n1499, ZN => n1492);
   U1616 : AOI22_X1 port map( A1 => n56, A2 => REGISTERS_29_14_port, B1 => n53,
                           B2 => REGISTERS_28_14_port, ZN => n1499);
   U1617 : OAI221_X1 port map( B1 => n2235, B2 => n62, C1 => n2203, C2 => n59, 
                           A => n1481, ZN => n1474);
   U1618 : AOI22_X1 port map( A1 => n56, A2 => REGISTERS_29_15_port, B1 => n53,
                           B2 => REGISTERS_28_15_port, ZN => n1481);
   U1619 : OAI221_X1 port map( B1 => n2234, B2 => n62, C1 => n2202, C2 => n59, 
                           A => n1463, ZN => n1456);
   U1620 : AOI22_X1 port map( A1 => n56, A2 => REGISTERS_29_16_port, B1 => n53,
                           B2 => REGISTERS_28_16_port, ZN => n1463);
   U1621 : OAI221_X1 port map( B1 => n2233, B2 => n62, C1 => n2201, C2 => n59, 
                           A => n1445, ZN => n1438);
   U1622 : AOI22_X1 port map( A1 => n56, A2 => REGISTERS_29_17_port, B1 => n53,
                           B2 => REGISTERS_28_17_port, ZN => n1445);
   U1623 : OAI221_X1 port map( B1 => n2232, B2 => n62, C1 => n2200, C2 => n59, 
                           A => n1427, ZN => n1420);
   U1624 : AOI22_X1 port map( A1 => n56, A2 => REGISTERS_29_18_port, B1 => n53,
                           B2 => REGISTERS_28_18_port, ZN => n1427);
   U1625 : OAI221_X1 port map( B1 => n2231, B2 => n62, C1 => n2199, C2 => n59, 
                           A => n1409, ZN => n1402);
   U1626 : AOI22_X1 port map( A1 => n56, A2 => REGISTERS_29_19_port, B1 => n53,
                           B2 => REGISTERS_28_19_port, ZN => n1409);
   U1627 : OAI221_X1 port map( B1 => n2230, B2 => n62, C1 => n2198, C2 => n59, 
                           A => n1391, ZN => n1384);
   U1628 : AOI22_X1 port map( A1 => n56, A2 => REGISTERS_29_20_port, B1 => n53,
                           B2 => REGISTERS_28_20_port, ZN => n1391);
   U1629 : OAI221_X1 port map( B1 => n2229, B2 => n62, C1 => n2197, C2 => n59, 
                           A => n1373, ZN => n1366);
   U1630 : AOI22_X1 port map( A1 => n56, A2 => REGISTERS_29_21_port, B1 => n53,
                           B2 => REGISTERS_28_21_port, ZN => n1373);
   U1631 : AOI22_X1 port map( A1 => REGISTERS_15_24_port, A2 => n105, B1 => 
                           REGISTERS_14_24_port, B2 => n102, ZN => n702);
   U1632 : AOI22_X1 port map( A1 => REGISTERS_15_25_port, A2 => n105, B1 => 
                           REGISTERS_14_25_port, B2 => n102, ZN => n684);
   U1633 : AOI22_X1 port map( A1 => REGISTERS_15_26_port, A2 => n105, B1 => 
                           REGISTERS_14_26_port, B2 => n102, ZN => n666);
   U1634 : AOI22_X1 port map( A1 => REGISTERS_15_27_port, A2 => n105, B1 => 
                           REGISTERS_14_27_port, B2 => n102, ZN => n648);
   U1635 : AOI22_X1 port map( A1 => REGISTERS_15_28_port, A2 => n105, B1 => 
                           REGISTERS_14_28_port, B2 => n102, ZN => n630);
   U1636 : AOI22_X1 port map( A1 => REGISTERS_15_29_port, A2 => n105, B1 => 
                           REGISTERS_14_29_port, B2 => n102, ZN => n612);
   U1637 : AOI22_X1 port map( A1 => REGISTERS_15_30_port, A2 => n105, B1 => 
                           REGISTERS_14_30_port, B2 => n102, ZN => n594);
   U1638 : AOI22_X1 port map( A1 => REGISTERS_15_31_port, A2 => n105, B1 => 
                           REGISTERS_14_31_port, B2 => n102, ZN => n574);
   U1639 : AOI22_X1 port map( A1 => REGISTERS_15_0_port, A2 => n103, B1 => 
                           REGISTERS_14_0_port, B2 => n100, ZN => n1149);
   U1640 : AOI22_X1 port map( A1 => REGISTERS_15_1_port, A2 => n103, B1 => 
                           REGISTERS_14_1_port, B2 => n100, ZN => n1116);
   U1641 : AOI22_X1 port map( A1 => REGISTERS_15_2_port, A2 => n103, B1 => 
                           REGISTERS_14_2_port, B2 => n100, ZN => n1098);
   U1642 : AOI22_X1 port map( A1 => REGISTERS_15_3_port, A2 => n103, B1 => 
                           REGISTERS_14_3_port, B2 => n100, ZN => n1080);
   U1643 : AOI22_X1 port map( A1 => REGISTERS_15_4_port, A2 => n103, B1 => 
                           REGISTERS_14_4_port, B2 => n100, ZN => n1062);
   U1644 : AOI22_X1 port map( A1 => REGISTERS_15_5_port, A2 => n103, B1 => 
                           REGISTERS_14_5_port, B2 => n100, ZN => n1044);
   U1645 : AOI22_X1 port map( A1 => REGISTERS_15_6_port, A2 => n103, B1 => 
                           REGISTERS_14_6_port, B2 => n100, ZN => n1026);
   U1646 : AOI22_X1 port map( A1 => REGISTERS_15_7_port, A2 => n103, B1 => 
                           REGISTERS_14_7_port, B2 => n100, ZN => n1008);
   U1647 : AOI22_X1 port map( A1 => REGISTERS_15_8_port, A2 => n103, B1 => 
                           REGISTERS_14_8_port, B2 => n100, ZN => n990);
   U1648 : AOI22_X1 port map( A1 => REGISTERS_15_9_port, A2 => n103, B1 => 
                           REGISTERS_14_9_port, B2 => n100, ZN => n972);
   U1649 : AOI22_X1 port map( A1 => REGISTERS_15_10_port, A2 => n103, B1 => 
                           REGISTERS_14_10_port, B2 => n100, ZN => n954);
   U1650 : AOI22_X1 port map( A1 => REGISTERS_15_11_port, A2 => n103, B1 => 
                           REGISTERS_14_11_port, B2 => n100, ZN => n936);
   U1651 : AOI22_X1 port map( A1 => REGISTERS_15_12_port, A2 => n104, B1 => 
                           REGISTERS_14_12_port, B2 => n101, ZN => n918);
   U1652 : AOI22_X1 port map( A1 => REGISTERS_15_13_port, A2 => n104, B1 => 
                           REGISTERS_14_13_port, B2 => n101, ZN => n900);
   U1653 : AOI22_X1 port map( A1 => REGISTERS_15_14_port, A2 => n104, B1 => 
                           REGISTERS_14_14_port, B2 => n101, ZN => n882);
   U1654 : AOI22_X1 port map( A1 => REGISTERS_15_15_port, A2 => n104, B1 => 
                           REGISTERS_14_15_port, B2 => n101, ZN => n864);
   U1655 : AOI22_X1 port map( A1 => REGISTERS_15_16_port, A2 => n104, B1 => 
                           REGISTERS_14_16_port, B2 => n101, ZN => n846);
   U1656 : AOI22_X1 port map( A1 => REGISTERS_15_17_port, A2 => n104, B1 => 
                           REGISTERS_14_17_port, B2 => n101, ZN => n828);
   U1657 : AOI22_X1 port map( A1 => REGISTERS_15_18_port, A2 => n104, B1 => 
                           REGISTERS_14_18_port, B2 => n101, ZN => n810);
   U1658 : AOI22_X1 port map( A1 => REGISTERS_15_19_port, A2 => n104, B1 => 
                           REGISTERS_14_19_port, B2 => n101, ZN => n792);
   U1659 : AOI22_X1 port map( A1 => REGISTERS_15_20_port, A2 => n104, B1 => 
                           REGISTERS_14_20_port, B2 => n101, ZN => n774);
   U1660 : AOI22_X1 port map( A1 => REGISTERS_15_21_port, A2 => n104, B1 => 
                           REGISTERS_14_21_port, B2 => n101, ZN => n756);
   U1661 : AOI22_X1 port map( A1 => REGISTERS_15_22_port, A2 => n104, B1 => 
                           REGISTERS_14_22_port, B2 => n101, ZN => n738);
   U1662 : AOI22_X1 port map( A1 => REGISTERS_15_23_port, A2 => n104, B1 => 
                           REGISTERS_14_23_port, B2 => n101, ZN => n720);
   U1663 : AOI22_X1 port map( A1 => n7, A2 => REGISTERS_15_0_port, B1 => n4, B2
                           => REGISTERS_14_0_port, ZN => n1774);
   U1664 : AOI22_X1 port map( A1 => n7, A2 => REGISTERS_15_1_port, B1 => n4, B2
                           => REGISTERS_14_1_port, ZN => n1741);
   U1665 : AOI22_X1 port map( A1 => n7, A2 => REGISTERS_15_2_port, B1 => n4, B2
                           => REGISTERS_14_2_port, ZN => n1723);
   U1666 : AOI22_X1 port map( A1 => n7, A2 => REGISTERS_15_3_port, B1 => n4, B2
                           => REGISTERS_14_3_port, ZN => n1705);
   U1667 : AOI22_X1 port map( A1 => n7, A2 => REGISTERS_15_4_port, B1 => n4, B2
                           => REGISTERS_14_4_port, ZN => n1687);
   U1668 : AOI22_X1 port map( A1 => n7, A2 => REGISTERS_15_5_port, B1 => n4, B2
                           => REGISTERS_14_5_port, ZN => n1669);
   U1669 : AOI22_X1 port map( A1 => n7, A2 => REGISTERS_15_6_port, B1 => n4, B2
                           => REGISTERS_14_6_port, ZN => n1651);
   U1670 : AOI22_X1 port map( A1 => n7, A2 => REGISTERS_15_7_port, B1 => n4, B2
                           => REGISTERS_14_7_port, ZN => n1633);
   U1671 : AOI22_X1 port map( A1 => n7, A2 => REGISTERS_15_8_port, B1 => n4, B2
                           => REGISTERS_14_8_port, ZN => n1615);
   U1672 : AOI22_X1 port map( A1 => n7, A2 => REGISTERS_15_9_port, B1 => n4, B2
                           => REGISTERS_14_9_port, ZN => n1597);
   U1673 : AOI22_X1 port map( A1 => n7, A2 => REGISTERS_15_10_port, B1 => n4, 
                           B2 => REGISTERS_14_10_port, ZN => n1579);
   U1674 : AOI22_X1 port map( A1 => n8, A2 => REGISTERS_15_11_port, B1 => n5, 
                           B2 => REGISTERS_14_11_port, ZN => n1561);
   U1675 : AOI22_X1 port map( A1 => n8, A2 => REGISTERS_15_12_port, B1 => n5, 
                           B2 => REGISTERS_14_12_port, ZN => n1543);
   U1676 : AOI22_X1 port map( A1 => n8, A2 => REGISTERS_15_13_port, B1 => n5, 
                           B2 => REGISTERS_14_13_port, ZN => n1525);
   U1677 : AOI22_X1 port map( A1 => n8, A2 => REGISTERS_15_14_port, B1 => n5, 
                           B2 => REGISTERS_14_14_port, ZN => n1507);
   U1678 : AOI22_X1 port map( A1 => n8, A2 => REGISTERS_15_15_port, B1 => n5, 
                           B2 => REGISTERS_14_15_port, ZN => n1489);
   U1679 : AOI22_X1 port map( A1 => n8, A2 => REGISTERS_15_16_port, B1 => n5, 
                           B2 => REGISTERS_14_16_port, ZN => n1471);
   U1680 : AOI22_X1 port map( A1 => n8, A2 => REGISTERS_15_17_port, B1 => n5, 
                           B2 => REGISTERS_14_17_port, ZN => n1453);
   U1681 : AOI22_X1 port map( A1 => n8, A2 => REGISTERS_15_18_port, B1 => n5, 
                           B2 => REGISTERS_14_18_port, ZN => n1435);
   U1682 : AOI22_X1 port map( A1 => n8, A2 => REGISTERS_15_19_port, B1 => n5, 
                           B2 => REGISTERS_14_19_port, ZN => n1417);
   U1683 : AOI22_X1 port map( A1 => n8, A2 => REGISTERS_15_20_port, B1 => n5, 
                           B2 => REGISTERS_14_20_port, ZN => n1399);
   U1684 : AOI22_X1 port map( A1 => n8, A2 => REGISTERS_15_21_port, B1 => n5, 
                           B2 => REGISTERS_14_21_port, ZN => n1381);
   U1685 : AOI22_X1 port map( A1 => n9, A2 => REGISTERS_15_22_port, B1 => n6, 
                           B2 => REGISTERS_14_22_port, ZN => n1363);
   U1686 : AOI22_X1 port map( A1 => n9, A2 => REGISTERS_15_23_port, B1 => n6, 
                           B2 => REGISTERS_14_23_port, ZN => n1345);
   U1687 : AOI22_X1 port map( A1 => n9, A2 => REGISTERS_15_24_port, B1 => n6, 
                           B2 => REGISTERS_14_24_port, ZN => n1327);
   U1688 : AOI22_X1 port map( A1 => n9, A2 => REGISTERS_15_25_port, B1 => n6, 
                           B2 => REGISTERS_14_25_port, ZN => n1309);
   U1689 : AOI22_X1 port map( A1 => n9, A2 => REGISTERS_15_26_port, B1 => n6, 
                           B2 => REGISTERS_14_26_port, ZN => n1291);
   U1690 : AOI22_X1 port map( A1 => n9, A2 => REGISTERS_15_27_port, B1 => n6, 
                           B2 => REGISTERS_14_27_port, ZN => n1273);
   U1691 : AOI22_X1 port map( A1 => n9, A2 => REGISTERS_15_28_port, B1 => n6, 
                           B2 => REGISTERS_14_28_port, ZN => n1255);
   U1692 : AOI22_X1 port map( A1 => n9, A2 => REGISTERS_15_29_port, B1 => n6, 
                           B2 => REGISTERS_14_29_port, ZN => n1237);
   U1693 : AOI22_X1 port map( A1 => n9, A2 => REGISTERS_15_30_port, B1 => n6, 
                           B2 => REGISTERS_14_30_port, ZN => n1219);
   U1694 : AOI22_X1 port map( A1 => n9, A2 => REGISTERS_15_31_port, B1 => n6, 
                           B2 => REGISTERS_14_31_port, ZN => n1199);
   U1695 : INV_X1 port map( A => ADD_WR(0), ZN => n2259);
   U1696 : INV_X1 port map( A => ADD_WR(1), ZN => n2260);
   U1697 : INV_X1 port map( A => ADD_WR(2), ZN => n2261);
   U1698 : INV_X1 port map( A => ADD_WR(3), ZN => n2262);
   U1699 : INV_X1 port map( A => ADD_WR(4), ZN => n2263);
   U1700 : OR3_X1 port map( A1 => ADD_WR(3), A2 => ADD_WR(4), A3 => n1786, ZN 
                           => n1777);
   U1701 : INV_X1 port map( A => REGISTERS_17_0_port, ZN => n2058);
   U1702 : INV_X1 port map( A => REGISTERS_21_0_port, ZN => n2122);
   U1703 : INV_X1 port map( A => REGISTERS_25_0_port, ZN => n2186);
   U1704 : INV_X1 port map( A => REGISTERS_31_0_port, ZN => n2250);
   U1705 : INV_X1 port map( A => REGISTERS_1_0_port, ZN => n1802);
   U1706 : INV_X1 port map( A => REGISTERS_5_0_port, ZN => n1866);
   U1707 : INV_X1 port map( A => REGISTERS_9_0_port, ZN => n1930);
   U1708 : INV_X1 port map( A => REGISTERS_13_0_port, ZN => n1994);
   U1709 : INV_X1 port map( A => REGISTERS_17_1_port, ZN => n2057);
   U1710 : INV_X1 port map( A => REGISTERS_21_1_port, ZN => n2121);
   U1711 : INV_X1 port map( A => REGISTERS_25_1_port, ZN => n2185);
   U1712 : INV_X1 port map( A => REGISTERS_31_1_port, ZN => n2249);
   U1713 : INV_X1 port map( A => REGISTERS_1_1_port, ZN => n1801);
   U1714 : INV_X1 port map( A => REGISTERS_5_1_port, ZN => n1865);
   U1715 : INV_X1 port map( A => REGISTERS_9_1_port, ZN => n1929);
   U1716 : INV_X1 port map( A => REGISTERS_13_1_port, ZN => n1993);
   U1717 : INV_X1 port map( A => REGISTERS_17_2_port, ZN => n2056);
   U1718 : INV_X1 port map( A => REGISTERS_21_2_port, ZN => n2120);
   U1719 : INV_X1 port map( A => REGISTERS_25_2_port, ZN => n2184);
   U1720 : INV_X1 port map( A => REGISTERS_31_2_port, ZN => n2248);
   U1721 : INV_X1 port map( A => REGISTERS_1_2_port, ZN => n1800);
   U1722 : INV_X1 port map( A => REGISTERS_5_2_port, ZN => n1864);
   U1723 : INV_X1 port map( A => REGISTERS_9_2_port, ZN => n1928);
   U1724 : INV_X1 port map( A => REGISTERS_13_2_port, ZN => n1992);
   U1725 : INV_X1 port map( A => REGISTERS_17_3_port, ZN => n2055);
   U1726 : INV_X1 port map( A => REGISTERS_21_3_port, ZN => n2119);
   U1727 : INV_X1 port map( A => REGISTERS_25_3_port, ZN => n2183);
   U1728 : INV_X1 port map( A => REGISTERS_31_3_port, ZN => n2247);
   U1729 : INV_X1 port map( A => REGISTERS_1_3_port, ZN => n1799);
   U1730 : INV_X1 port map( A => REGISTERS_5_3_port, ZN => n1863);
   U1731 : INV_X1 port map( A => REGISTERS_9_3_port, ZN => n1927);
   U1732 : INV_X1 port map( A => REGISTERS_13_3_port, ZN => n1991);
   U1733 : INV_X1 port map( A => REGISTERS_17_4_port, ZN => n2054);
   U1734 : INV_X1 port map( A => REGISTERS_21_4_port, ZN => n2118);
   U1735 : INV_X1 port map( A => REGISTERS_25_4_port, ZN => n2182);
   U1736 : INV_X1 port map( A => REGISTERS_31_4_port, ZN => n2246);
   U1737 : INV_X1 port map( A => REGISTERS_1_4_port, ZN => n1798);
   U1738 : INV_X1 port map( A => REGISTERS_5_4_port, ZN => n1862);
   U1739 : INV_X1 port map( A => REGISTERS_9_4_port, ZN => n1926);
   U1740 : INV_X1 port map( A => REGISTERS_13_4_port, ZN => n1990);
   U1741 : INV_X1 port map( A => REGISTERS_17_5_port, ZN => n2053);
   U1742 : INV_X1 port map( A => REGISTERS_21_5_port, ZN => n2117);
   U1743 : INV_X1 port map( A => REGISTERS_25_5_port, ZN => n2181);
   U1744 : INV_X1 port map( A => REGISTERS_31_5_port, ZN => n2245);
   U1745 : INV_X1 port map( A => REGISTERS_1_5_port, ZN => n1797);
   U1746 : INV_X1 port map( A => REGISTERS_5_5_port, ZN => n1861);
   U1747 : INV_X1 port map( A => REGISTERS_9_5_port, ZN => n1925);
   U1748 : INV_X1 port map( A => REGISTERS_13_5_port, ZN => n1989);
   U1749 : INV_X1 port map( A => REGISTERS_17_6_port, ZN => n2052);
   U1750 : INV_X1 port map( A => REGISTERS_21_6_port, ZN => n2116);
   U1751 : INV_X1 port map( A => REGISTERS_25_6_port, ZN => n2180);
   U1752 : INV_X1 port map( A => REGISTERS_31_6_port, ZN => n2244);
   U1753 : INV_X1 port map( A => REGISTERS_1_6_port, ZN => n1796);
   U1754 : INV_X1 port map( A => REGISTERS_5_6_port, ZN => n1860);
   U1755 : INV_X1 port map( A => REGISTERS_9_6_port, ZN => n1924);
   U1756 : INV_X1 port map( A => REGISTERS_13_6_port, ZN => n1988);
   U1757 : INV_X1 port map( A => REGISTERS_17_7_port, ZN => n2051);
   U1758 : INV_X1 port map( A => REGISTERS_21_7_port, ZN => n2115);
   U1759 : INV_X1 port map( A => REGISTERS_25_7_port, ZN => n2179);
   U1760 : INV_X1 port map( A => REGISTERS_31_7_port, ZN => n2243);
   U1761 : INV_X1 port map( A => REGISTERS_1_7_port, ZN => n1795);
   U1762 : INV_X1 port map( A => REGISTERS_5_7_port, ZN => n1859);
   U1763 : INV_X1 port map( A => REGISTERS_9_7_port, ZN => n1923);
   U1764 : INV_X1 port map( A => REGISTERS_13_7_port, ZN => n1987);
   U1765 : INV_X1 port map( A => REGISTERS_17_8_port, ZN => n2050);
   U1766 : INV_X1 port map( A => REGISTERS_21_8_port, ZN => n2114);
   U1767 : INV_X1 port map( A => REGISTERS_25_8_port, ZN => n2178);
   U1768 : INV_X1 port map( A => REGISTERS_31_8_port, ZN => n2242);
   U1769 : INV_X1 port map( A => REGISTERS_1_8_port, ZN => n1794);
   U1770 : INV_X1 port map( A => REGISTERS_5_8_port, ZN => n1858);
   U1771 : INV_X1 port map( A => REGISTERS_9_8_port, ZN => n1922);
   U1772 : INV_X1 port map( A => REGISTERS_13_8_port, ZN => n1986);
   U1773 : INV_X1 port map( A => REGISTERS_17_9_port, ZN => n2049);
   U1774 : INV_X1 port map( A => REGISTERS_21_9_port, ZN => n2113);
   U1775 : INV_X1 port map( A => REGISTERS_25_9_port, ZN => n2177);
   U1776 : INV_X1 port map( A => REGISTERS_31_9_port, ZN => n2241);
   U1777 : INV_X1 port map( A => REGISTERS_1_9_port, ZN => n1793);
   U1778 : INV_X1 port map( A => REGISTERS_5_9_port, ZN => n1857);
   U1779 : INV_X1 port map( A => REGISTERS_9_9_port, ZN => n1921);
   U1780 : INV_X1 port map( A => REGISTERS_13_9_port, ZN => n1985);
   U1781 : INV_X1 port map( A => REGISTERS_17_10_port, ZN => n2048);
   U1782 : INV_X1 port map( A => REGISTERS_21_10_port, ZN => n2112);
   U1783 : INV_X1 port map( A => REGISTERS_25_10_port, ZN => n2176);
   U1784 : INV_X1 port map( A => REGISTERS_31_10_port, ZN => n2240);
   U1785 : INV_X1 port map( A => REGISTERS_1_10_port, ZN => n1792);
   U1786 : INV_X1 port map( A => REGISTERS_5_10_port, ZN => n1856);
   U1787 : INV_X1 port map( A => REGISTERS_9_10_port, ZN => n1920);
   U1788 : INV_X1 port map( A => REGISTERS_13_10_port, ZN => n1984);
   U1789 : INV_X1 port map( A => REGISTERS_17_11_port, ZN => n2047);
   U1790 : INV_X1 port map( A => REGISTERS_21_11_port, ZN => n2111);
   U1791 : INV_X1 port map( A => REGISTERS_25_11_port, ZN => n2175);
   U1792 : INV_X1 port map( A => REGISTERS_31_11_port, ZN => n2239);
   U1793 : INV_X1 port map( A => REGISTERS_1_11_port, ZN => n1791);
   U1794 : INV_X1 port map( A => REGISTERS_5_11_port, ZN => n1855);
   U1795 : INV_X1 port map( A => REGISTERS_9_11_port, ZN => n1919);
   U1796 : INV_X1 port map( A => REGISTERS_13_11_port, ZN => n1983);
   U1797 : INV_X1 port map( A => REGISTERS_17_12_port, ZN => n2046);
   U1798 : INV_X1 port map( A => REGISTERS_21_12_port, ZN => n2110);
   U1799 : INV_X1 port map( A => REGISTERS_25_12_port, ZN => n2174);
   U1800 : INV_X1 port map( A => REGISTERS_31_12_port, ZN => n2238);
   U1801 : INV_X1 port map( A => REGISTERS_1_12_port, ZN => n526);
   U1802 : INV_X1 port map( A => REGISTERS_5_12_port, ZN => n1854);
   U1803 : INV_X1 port map( A => REGISTERS_9_12_port, ZN => n1918);
   U1804 : INV_X1 port map( A => REGISTERS_13_12_port, ZN => n1982);
   U1805 : INV_X1 port map( A => REGISTERS_17_13_port, ZN => n2045);
   U1806 : INV_X1 port map( A => REGISTERS_21_13_port, ZN => n2109);
   U1807 : INV_X1 port map( A => REGISTERS_25_13_port, ZN => n2173);
   U1808 : INV_X1 port map( A => REGISTERS_31_13_port, ZN => n2237);
   U1809 : INV_X1 port map( A => REGISTERS_1_13_port, ZN => n525);
   U1810 : INV_X1 port map( A => REGISTERS_5_13_port, ZN => n1853);
   U1811 : INV_X1 port map( A => REGISTERS_9_13_port, ZN => n1917);
   U1812 : INV_X1 port map( A => REGISTERS_13_13_port, ZN => n1981);
   U1813 : INV_X1 port map( A => REGISTERS_17_14_port, ZN => n2044);
   U1814 : INV_X1 port map( A => REGISTERS_21_14_port, ZN => n2108);
   U1815 : INV_X1 port map( A => REGISTERS_25_14_port, ZN => n2172);
   U1816 : INV_X1 port map( A => REGISTERS_31_14_port, ZN => n2236);
   U1817 : INV_X1 port map( A => REGISTERS_1_14_port, ZN => n524);
   U1818 : INV_X1 port map( A => REGISTERS_5_14_port, ZN => n1852);
   U1819 : INV_X1 port map( A => REGISTERS_9_14_port, ZN => n1916);
   U1820 : INV_X1 port map( A => REGISTERS_13_14_port, ZN => n1980);
   U1821 : INV_X1 port map( A => REGISTERS_17_15_port, ZN => n2043);
   U1822 : INV_X1 port map( A => REGISTERS_21_15_port, ZN => n2107);
   U1823 : INV_X1 port map( A => REGISTERS_25_15_port, ZN => n2171);
   U1824 : INV_X1 port map( A => REGISTERS_31_15_port, ZN => n2235);
   U1825 : INV_X1 port map( A => REGISTERS_1_15_port, ZN => n523);
   U1826 : INV_X1 port map( A => REGISTERS_5_15_port, ZN => n1851);
   U1827 : INV_X1 port map( A => REGISTERS_9_15_port, ZN => n1915);
   U1828 : INV_X1 port map( A => REGISTERS_13_15_port, ZN => n1979);
   U1829 : INV_X1 port map( A => REGISTERS_17_16_port, ZN => n2042);
   U1830 : INV_X1 port map( A => REGISTERS_21_16_port, ZN => n2106);
   U1831 : INV_X1 port map( A => REGISTERS_25_16_port, ZN => n2170);
   U1832 : INV_X1 port map( A => REGISTERS_31_16_port, ZN => n2234);
   U1833 : INV_X1 port map( A => REGISTERS_1_16_port, ZN => n522);
   U1834 : INV_X1 port map( A => REGISTERS_5_16_port, ZN => n1850);
   U1835 : INV_X1 port map( A => REGISTERS_9_16_port, ZN => n1914);
   U1836 : INV_X1 port map( A => REGISTERS_13_16_port, ZN => n1978);
   U1837 : INV_X1 port map( A => REGISTERS_17_17_port, ZN => n2041);
   U1838 : INV_X1 port map( A => REGISTERS_21_17_port, ZN => n2105);
   U1839 : INV_X1 port map( A => REGISTERS_25_17_port, ZN => n2169);
   U1840 : INV_X1 port map( A => REGISTERS_31_17_port, ZN => n2233);
   U1841 : INV_X1 port map( A => REGISTERS_1_17_port, ZN => n521);
   U1842 : INV_X1 port map( A => REGISTERS_5_17_port, ZN => n1849);
   U1843 : INV_X1 port map( A => REGISTERS_9_17_port, ZN => n1913);
   U1844 : INV_X1 port map( A => REGISTERS_13_17_port, ZN => n1977);
   U1845 : INV_X1 port map( A => REGISTERS_17_18_port, ZN => n2040);
   U1846 : INV_X1 port map( A => REGISTERS_21_18_port, ZN => n2104);
   U1847 : INV_X1 port map( A => REGISTERS_25_18_port, ZN => n2168);
   U1848 : INV_X1 port map( A => REGISTERS_31_18_port, ZN => n2232);
   U1849 : INV_X1 port map( A => REGISTERS_1_18_port, ZN => n520);
   U1850 : INV_X1 port map( A => REGISTERS_5_18_port, ZN => n1848);
   U1851 : INV_X1 port map( A => REGISTERS_9_18_port, ZN => n1912);
   U1852 : INV_X1 port map( A => REGISTERS_13_18_port, ZN => n1976);
   U1853 : INV_X1 port map( A => REGISTERS_17_19_port, ZN => n2039);
   U1854 : INV_X1 port map( A => REGISTERS_21_19_port, ZN => n2103);
   U1855 : INV_X1 port map( A => REGISTERS_25_19_port, ZN => n2167);
   U1856 : INV_X1 port map( A => REGISTERS_31_19_port, ZN => n2231);
   U1857 : INV_X1 port map( A => REGISTERS_1_19_port, ZN => n519);
   U1858 : INV_X1 port map( A => REGISTERS_5_19_port, ZN => n1847);
   U1859 : INV_X1 port map( A => REGISTERS_9_19_port, ZN => n1911);
   U1860 : INV_X1 port map( A => REGISTERS_13_19_port, ZN => n1975);
   U1861 : INV_X1 port map( A => REGISTERS_17_20_port, ZN => n2038);
   U1862 : INV_X1 port map( A => REGISTERS_21_20_port, ZN => n2102);
   U1863 : INV_X1 port map( A => REGISTERS_25_20_port, ZN => n2166);
   U1864 : INV_X1 port map( A => REGISTERS_31_20_port, ZN => n2230);
   U1865 : INV_X1 port map( A => REGISTERS_1_20_port, ZN => n518);
   U1866 : INV_X1 port map( A => REGISTERS_5_20_port, ZN => n1846);
   U1867 : INV_X1 port map( A => REGISTERS_9_20_port, ZN => n1910);
   U1868 : INV_X1 port map( A => REGISTERS_13_20_port, ZN => n1974);
   U1869 : INV_X1 port map( A => REGISTERS_17_21_port, ZN => n2037);
   U1870 : INV_X1 port map( A => REGISTERS_21_21_port, ZN => n2101);
   U1871 : INV_X1 port map( A => REGISTERS_25_21_port, ZN => n2165);
   U1872 : INV_X1 port map( A => REGISTERS_31_21_port, ZN => n2229);
   U1873 : INV_X1 port map( A => REGISTERS_1_21_port, ZN => n517);
   U1874 : INV_X1 port map( A => REGISTERS_5_21_port, ZN => n1845);
   U1875 : INV_X1 port map( A => REGISTERS_9_21_port, ZN => n1909);
   U1876 : INV_X1 port map( A => REGISTERS_13_21_port, ZN => n1973);
   U1877 : INV_X1 port map( A => REGISTERS_17_22_port, ZN => n2036);
   U1878 : INV_X1 port map( A => REGISTERS_21_22_port, ZN => n2100);
   U1879 : INV_X1 port map( A => REGISTERS_25_22_port, ZN => n2164);
   U1880 : INV_X1 port map( A => REGISTERS_31_22_port, ZN => n2228);
   U1881 : INV_X1 port map( A => REGISTERS_1_22_port, ZN => n516);
   U1882 : INV_X1 port map( A => REGISTERS_5_22_port, ZN => n1844);
   U1883 : INV_X1 port map( A => REGISTERS_9_22_port, ZN => n1908);
   U1884 : INV_X1 port map( A => REGISTERS_13_22_port, ZN => n1972);
   U1885 : INV_X1 port map( A => REGISTERS_17_23_port, ZN => n2035);
   U1886 : INV_X1 port map( A => REGISTERS_21_23_port, ZN => n2099);
   U1887 : INV_X1 port map( A => REGISTERS_25_23_port, ZN => n2163);
   U1888 : INV_X1 port map( A => REGISTERS_31_23_port, ZN => n2227);
   U1889 : INV_X1 port map( A => REGISTERS_1_23_port, ZN => n515);
   U1890 : INV_X1 port map( A => REGISTERS_5_23_port, ZN => n1843);
   U1891 : INV_X1 port map( A => REGISTERS_9_23_port, ZN => n1907);
   U1892 : INV_X1 port map( A => REGISTERS_13_23_port, ZN => n1971);
   U1893 : INV_X1 port map( A => REGISTERS_17_24_port, ZN => n2034);
   U1894 : INV_X1 port map( A => REGISTERS_21_24_port, ZN => n2098);
   U1895 : INV_X1 port map( A => REGISTERS_25_24_port, ZN => n2162);
   U1896 : INV_X1 port map( A => REGISTERS_31_24_port, ZN => n2226);
   U1897 : INV_X1 port map( A => REGISTERS_1_24_port, ZN => n514);
   U1898 : INV_X1 port map( A => REGISTERS_5_24_port, ZN => n1842);
   U1899 : INV_X1 port map( A => REGISTERS_9_24_port, ZN => n1906);
   U1900 : INV_X1 port map( A => REGISTERS_13_24_port, ZN => n1970);
   U1901 : INV_X1 port map( A => REGISTERS_17_25_port, ZN => n2033);
   U1902 : INV_X1 port map( A => REGISTERS_21_25_port, ZN => n2097);
   U1903 : INV_X1 port map( A => REGISTERS_25_25_port, ZN => n2161);
   U1904 : INV_X1 port map( A => REGISTERS_31_25_port, ZN => n2225);
   U1905 : INV_X1 port map( A => REGISTERS_1_25_port, ZN => n513);
   U1906 : INV_X1 port map( A => REGISTERS_5_25_port, ZN => n1841);
   U1907 : INV_X1 port map( A => REGISTERS_9_25_port, ZN => n1905);
   U1908 : INV_X1 port map( A => REGISTERS_13_25_port, ZN => n1969);
   U1909 : INV_X1 port map( A => REGISTERS_17_26_port, ZN => n2032);
   U1910 : INV_X1 port map( A => REGISTERS_21_26_port, ZN => n2096);
   U1923 : INV_X1 port map( A => REGISTERS_25_26_port, ZN => n2160);
   U1924 : INV_X1 port map( A => REGISTERS_31_26_port, ZN => n2224);
   U1925 : INV_X1 port map( A => REGISTERS_1_26_port, ZN => n512);
   U1926 : INV_X1 port map( A => REGISTERS_5_26_port, ZN => n1840);
   U1927 : INV_X1 port map( A => REGISTERS_9_26_port, ZN => n1904);
   U1928 : INV_X1 port map( A => REGISTERS_13_26_port, ZN => n1968);
   U1929 : INV_X1 port map( A => REGISTERS_17_27_port, ZN => n2031);
   U1930 : INV_X1 port map( A => REGISTERS_21_27_port, ZN => n2095);
   U1931 : INV_X1 port map( A => REGISTERS_25_27_port, ZN => n2159);
   U1932 : INV_X1 port map( A => REGISTERS_31_27_port, ZN => n2223);
   U1933 : INV_X1 port map( A => REGISTERS_1_27_port, ZN => n511);
   U1934 : INV_X1 port map( A => REGISTERS_5_27_port, ZN => n1839);
   U1935 : INV_X1 port map( A => REGISTERS_9_27_port, ZN => n1903);
   U1936 : INV_X1 port map( A => REGISTERS_13_27_port, ZN => n1967);
   U1937 : INV_X1 port map( A => REGISTERS_17_28_port, ZN => n2030);
   U1938 : INV_X1 port map( A => REGISTERS_21_28_port, ZN => n2094);
   U1939 : INV_X1 port map( A => REGISTERS_25_28_port, ZN => n2158);
   U1940 : INV_X1 port map( A => REGISTERS_31_28_port, ZN => n2222);
   U1941 : INV_X1 port map( A => REGISTERS_1_28_port, ZN => n510);
   U1942 : INV_X1 port map( A => REGISTERS_5_28_port, ZN => n1838);
   U1943 : INV_X1 port map( A => REGISTERS_9_28_port, ZN => n1902);
   U1944 : INV_X1 port map( A => REGISTERS_13_28_port, ZN => n1966);
   U1945 : INV_X1 port map( A => REGISTERS_17_29_port, ZN => n2029);
   U1946 : INV_X1 port map( A => REGISTERS_21_29_port, ZN => n2093);
   U1947 : INV_X1 port map( A => REGISTERS_25_29_port, ZN => n2157);
   U1948 : INV_X1 port map( A => REGISTERS_31_29_port, ZN => n2221);
   U1949 : INV_X1 port map( A => REGISTERS_1_29_port, ZN => n509);
   U1950 : INV_X1 port map( A => REGISTERS_5_29_port, ZN => n1837);
   U1951 : INV_X1 port map( A => REGISTERS_9_29_port, ZN => n1901);
   U1952 : INV_X1 port map( A => REGISTERS_13_29_port, ZN => n1965);
   U1953 : INV_X1 port map( A => REGISTERS_17_30_port, ZN => n2028);
   U1954 : INV_X1 port map( A => REGISTERS_21_30_port, ZN => n2092);
   U1955 : INV_X1 port map( A => REGISTERS_25_30_port, ZN => n2156);
   U1956 : INV_X1 port map( A => REGISTERS_31_30_port, ZN => n2220);
   U1957 : INV_X1 port map( A => REGISTERS_1_30_port, ZN => n508);
   U1958 : INV_X1 port map( A => REGISTERS_5_30_port, ZN => n1836);
   U1959 : INV_X1 port map( A => REGISTERS_9_30_port, ZN => n1900);
   U1960 : INV_X1 port map( A => REGISTERS_13_30_port, ZN => n1964);
   U1961 : INV_X1 port map( A => REGISTERS_17_31_port, ZN => n2027);
   U1962 : INV_X1 port map( A => REGISTERS_21_31_port, ZN => n2091);
   U1963 : INV_X1 port map( A => REGISTERS_25_31_port, ZN => n2155);
   U1964 : INV_X1 port map( A => REGISTERS_31_31_port, ZN => n2219);
   U1965 : INV_X1 port map( A => REGISTERS_1_31_port, ZN => n507);
   U1966 : INV_X1 port map( A => REGISTERS_5_31_port, ZN => n1835);
   U1967 : INV_X1 port map( A => REGISTERS_9_31_port, ZN => n1899);
   U1968 : INV_X1 port map( A => REGISTERS_13_31_port, ZN => n1963);
   U1969 : INV_X1 port map( A => REGISTERS_16_0_port, ZN => n2026);
   U1970 : INV_X1 port map( A => REGISTERS_20_0_port, ZN => n2090);
   U1971 : INV_X1 port map( A => REGISTERS_24_0_port, ZN => n2154);
   U1972 : INV_X1 port map( A => REGISTERS_30_0_port, ZN => n2218);
   U1973 : INV_X1 port map( A => REGISTERS_0_0_port, ZN => n506);
   U1974 : INV_X1 port map( A => REGISTERS_4_0_port, ZN => n1834);
   U1975 : INV_X1 port map( A => REGISTERS_8_0_port, ZN => n1898);
   U1976 : INV_X1 port map( A => REGISTERS_12_0_port, ZN => n1962);
   U1977 : INV_X1 port map( A => REGISTERS_16_1_port, ZN => n2025);
   U1978 : INV_X1 port map( A => REGISTERS_20_1_port, ZN => n2089);
   U1979 : INV_X1 port map( A => REGISTERS_24_1_port, ZN => n2153);
   U1980 : INV_X1 port map( A => REGISTERS_30_1_port, ZN => n2217);
   U1981 : INV_X1 port map( A => REGISTERS_0_1_port, ZN => n505);
   U1982 : INV_X1 port map( A => REGISTERS_4_1_port, ZN => n1833);
   U1983 : INV_X1 port map( A => REGISTERS_8_1_port, ZN => n1897);
   U1984 : INV_X1 port map( A => REGISTERS_12_1_port, ZN => n1961);
   U1985 : INV_X1 port map( A => REGISTERS_16_2_port, ZN => n2024);
   U1986 : INV_X1 port map( A => REGISTERS_20_2_port, ZN => n2088);
   U1987 : INV_X1 port map( A => REGISTERS_24_2_port, ZN => n2152);
   U1988 : INV_X1 port map( A => REGISTERS_30_2_port, ZN => n2216);
   U1989 : INV_X1 port map( A => REGISTERS_0_2_port, ZN => n504);
   U1990 : INV_X1 port map( A => REGISTERS_4_2_port, ZN => n1832);
   U1991 : INV_X1 port map( A => REGISTERS_8_2_port, ZN => n1896);
   U1992 : INV_X1 port map( A => REGISTERS_12_2_port, ZN => n1960);
   U1993 : INV_X1 port map( A => REGISTERS_16_3_port, ZN => n2023);
   U1994 : INV_X1 port map( A => REGISTERS_20_3_port, ZN => n2087);
   U1995 : INV_X1 port map( A => REGISTERS_24_3_port, ZN => n2151);
   U1996 : INV_X1 port map( A => REGISTERS_30_3_port, ZN => n2215);
   U1997 : INV_X1 port map( A => REGISTERS_0_3_port, ZN => n503);
   U1998 : INV_X1 port map( A => REGISTERS_4_3_port, ZN => n1831);
   U1999 : INV_X1 port map( A => REGISTERS_8_3_port, ZN => n1895);
   U2000 : INV_X1 port map( A => REGISTERS_12_3_port, ZN => n1959);
   U2001 : INV_X1 port map( A => REGISTERS_16_4_port, ZN => n2022);
   U2002 : INV_X1 port map( A => REGISTERS_20_4_port, ZN => n2086);
   U2003 : INV_X1 port map( A => REGISTERS_24_4_port, ZN => n2150);
   U2004 : INV_X1 port map( A => REGISTERS_30_4_port, ZN => n2214);
   U2005 : INV_X1 port map( A => REGISTERS_0_4_port, ZN => n502);
   U2006 : INV_X1 port map( A => REGISTERS_4_4_port, ZN => n1830);
   U2007 : INV_X1 port map( A => REGISTERS_8_4_port, ZN => n1894);
   U2008 : INV_X1 port map( A => REGISTERS_12_4_port, ZN => n1958);
   U2009 : INV_X1 port map( A => REGISTERS_16_5_port, ZN => n2021);
   U2010 : INV_X1 port map( A => REGISTERS_20_5_port, ZN => n2085);
   U2011 : INV_X1 port map( A => REGISTERS_24_5_port, ZN => n2149);
   U2012 : INV_X1 port map( A => REGISTERS_30_5_port, ZN => n2213);
   U2013 : INV_X1 port map( A => REGISTERS_0_5_port, ZN => n501);
   U2014 : INV_X1 port map( A => REGISTERS_4_5_port, ZN => n1829);
   U2015 : INV_X1 port map( A => REGISTERS_8_5_port, ZN => n1893);
   U2016 : INV_X1 port map( A => REGISTERS_12_5_port, ZN => n1957);
   U2017 : INV_X1 port map( A => REGISTERS_16_6_port, ZN => n2020);
   U2018 : INV_X1 port map( A => REGISTERS_20_6_port, ZN => n2084);
   U2019 : INV_X1 port map( A => REGISTERS_24_6_port, ZN => n2148);
   U2020 : INV_X1 port map( A => REGISTERS_30_6_port, ZN => n2212);
   U2021 : INV_X1 port map( A => REGISTERS_0_6_port, ZN => n500);
   U2022 : INV_X1 port map( A => REGISTERS_4_6_port, ZN => n1828);
   U2023 : INV_X1 port map( A => REGISTERS_8_6_port, ZN => n1892);
   U2024 : INV_X1 port map( A => REGISTERS_12_6_port, ZN => n1956);
   U2025 : INV_X1 port map( A => REGISTERS_16_7_port, ZN => n2019);
   U2026 : INV_X1 port map( A => REGISTERS_20_7_port, ZN => n2083);
   U2027 : INV_X1 port map( A => REGISTERS_24_7_port, ZN => n2147);
   U2028 : INV_X1 port map( A => REGISTERS_30_7_port, ZN => n2211);
   U2029 : INV_X1 port map( A => REGISTERS_0_7_port, ZN => n499);
   U2030 : INV_X1 port map( A => REGISTERS_4_7_port, ZN => n1827);
   U2031 : INV_X1 port map( A => REGISTERS_8_7_port, ZN => n1891);
   U2032 : INV_X1 port map( A => REGISTERS_12_7_port, ZN => n1955);
   U2033 : INV_X1 port map( A => REGISTERS_16_8_port, ZN => n2018);
   U2034 : INV_X1 port map( A => REGISTERS_20_8_port, ZN => n2082);
   U2035 : INV_X1 port map( A => REGISTERS_24_8_port, ZN => n2146);
   U2036 : INV_X1 port map( A => REGISTERS_30_8_port, ZN => n2210);
   U2037 : INV_X1 port map( A => REGISTERS_0_8_port, ZN => n498);
   U2038 : INV_X1 port map( A => REGISTERS_4_8_port, ZN => n1826);
   U2039 : INV_X1 port map( A => REGISTERS_8_8_port, ZN => n1890);
   U2040 : INV_X1 port map( A => REGISTERS_12_8_port, ZN => n1954);
   U2041 : INV_X1 port map( A => REGISTERS_16_9_port, ZN => n2017);
   U2042 : INV_X1 port map( A => REGISTERS_20_9_port, ZN => n2081);
   U2043 : INV_X1 port map( A => REGISTERS_24_9_port, ZN => n2145);
   U2044 : INV_X1 port map( A => REGISTERS_30_9_port, ZN => n2209);
   U2045 : INV_X1 port map( A => REGISTERS_0_9_port, ZN => n497);
   U2046 : INV_X1 port map( A => REGISTERS_4_9_port, ZN => n1825);
   U2047 : INV_X1 port map( A => REGISTERS_8_9_port, ZN => n1889);
   U2048 : INV_X1 port map( A => REGISTERS_12_9_port, ZN => n1953);
   U2049 : INV_X1 port map( A => REGISTERS_16_10_port, ZN => n2016);
   U2050 : INV_X1 port map( A => REGISTERS_20_10_port, ZN => n2080);
   U2051 : INV_X1 port map( A => REGISTERS_24_10_port, ZN => n2144);
   U2052 : INV_X1 port map( A => REGISTERS_30_10_port, ZN => n2208);
   U2053 : INV_X1 port map( A => REGISTERS_0_10_port, ZN => n496);
   U2054 : INV_X1 port map( A => REGISTERS_4_10_port, ZN => n1824);
   U2055 : INV_X1 port map( A => REGISTERS_8_10_port, ZN => n1888);
   U2056 : INV_X1 port map( A => REGISTERS_12_10_port, ZN => n1952);
   U2057 : INV_X1 port map( A => REGISTERS_16_11_port, ZN => n2015);
   U2058 : INV_X1 port map( A => REGISTERS_20_11_port, ZN => n2079);
   U2059 : INV_X1 port map( A => REGISTERS_24_11_port, ZN => n2143);
   U2060 : INV_X1 port map( A => REGISTERS_30_11_port, ZN => n2207);
   U2061 : INV_X1 port map( A => REGISTERS_0_11_port, ZN => n495);
   U2062 : INV_X1 port map( A => REGISTERS_4_11_port, ZN => n1823);
   U2063 : INV_X1 port map( A => REGISTERS_8_11_port, ZN => n1887);
   U2064 : INV_X1 port map( A => REGISTERS_12_11_port, ZN => n1951);
   U2065 : INV_X1 port map( A => REGISTERS_16_12_port, ZN => n2014);
   U2066 : INV_X1 port map( A => REGISTERS_20_12_port, ZN => n2078);
   U2067 : INV_X1 port map( A => REGISTERS_24_12_port, ZN => n2142);
   U2068 : INV_X1 port map( A => REGISTERS_30_12_port, ZN => n2206);
   U2069 : INV_X1 port map( A => REGISTERS_0_12_port, ZN => n494);
   U2070 : INV_X1 port map( A => REGISTERS_4_12_port, ZN => n1822);
   U2071 : INV_X1 port map( A => REGISTERS_8_12_port, ZN => n1886);
   U2072 : INV_X1 port map( A => REGISTERS_12_12_port, ZN => n1950);
   U2073 : INV_X1 port map( A => REGISTERS_16_13_port, ZN => n2013);
   U2074 : INV_X1 port map( A => REGISTERS_20_13_port, ZN => n2077);
   U2075 : INV_X1 port map( A => REGISTERS_24_13_port, ZN => n2141);
   U2076 : INV_X1 port map( A => REGISTERS_30_13_port, ZN => n2205);
   U2077 : INV_X1 port map( A => REGISTERS_0_13_port, ZN => n493);
   U2078 : INV_X1 port map( A => REGISTERS_4_13_port, ZN => n1821);
   U2079 : INV_X1 port map( A => REGISTERS_8_13_port, ZN => n1885);
   U2080 : INV_X1 port map( A => REGISTERS_12_13_port, ZN => n1949);
   U2081 : INV_X1 port map( A => REGISTERS_16_14_port, ZN => n2012);
   U2082 : INV_X1 port map( A => REGISTERS_20_14_port, ZN => n2076);
   U2083 : INV_X1 port map( A => REGISTERS_24_14_port, ZN => n2140);
   U2084 : INV_X1 port map( A => REGISTERS_30_14_port, ZN => n2204);
   U2085 : INV_X1 port map( A => REGISTERS_0_14_port, ZN => n492);
   U2086 : INV_X1 port map( A => REGISTERS_4_14_port, ZN => n1820);
   U2087 : INV_X1 port map( A => REGISTERS_8_14_port, ZN => n1884);
   U2088 : INV_X1 port map( A => REGISTERS_12_14_port, ZN => n1948);
   U2089 : INV_X1 port map( A => REGISTERS_16_15_port, ZN => n2011);
   U2090 : INV_X1 port map( A => REGISTERS_20_15_port, ZN => n2075);
   U2091 : INV_X1 port map( A => REGISTERS_24_15_port, ZN => n2139);
   U2092 : INV_X1 port map( A => REGISTERS_30_15_port, ZN => n2203);
   U2093 : INV_X1 port map( A => REGISTERS_0_15_port, ZN => n491);
   U2094 : INV_X1 port map( A => REGISTERS_4_15_port, ZN => n1819);
   U2095 : INV_X1 port map( A => REGISTERS_8_15_port, ZN => n1883);
   U2096 : INV_X1 port map( A => REGISTERS_12_15_port, ZN => n1947);
   U2097 : INV_X1 port map( A => REGISTERS_16_16_port, ZN => n2010);
   U2098 : INV_X1 port map( A => REGISTERS_20_16_port, ZN => n2074);
   U2099 : INV_X1 port map( A => REGISTERS_24_16_port, ZN => n2138);
   U2100 : INV_X1 port map( A => REGISTERS_30_16_port, ZN => n2202);
   U2101 : INV_X1 port map( A => REGISTERS_0_16_port, ZN => n490);
   U2102 : INV_X1 port map( A => REGISTERS_4_16_port, ZN => n1818);
   U2103 : INV_X1 port map( A => REGISTERS_8_16_port, ZN => n1882);
   U2104 : INV_X1 port map( A => REGISTERS_12_16_port, ZN => n1946);
   U2105 : INV_X1 port map( A => REGISTERS_16_17_port, ZN => n2009);
   U2106 : INV_X1 port map( A => REGISTERS_20_17_port, ZN => n2073);
   U2107 : INV_X1 port map( A => REGISTERS_24_17_port, ZN => n2137);
   U2108 : INV_X1 port map( A => REGISTERS_30_17_port, ZN => n2201);
   U2109 : INV_X1 port map( A => REGISTERS_0_17_port, ZN => n489);
   U2110 : INV_X1 port map( A => REGISTERS_4_17_port, ZN => n1817);
   U2111 : INV_X1 port map( A => REGISTERS_8_17_port, ZN => n1881);
   U2112 : INV_X1 port map( A => REGISTERS_12_17_port, ZN => n1945);
   U2113 : INV_X1 port map( A => REGISTERS_16_18_port, ZN => n2008);
   U2114 : INV_X1 port map( A => REGISTERS_20_18_port, ZN => n2072);
   U2115 : INV_X1 port map( A => REGISTERS_24_18_port, ZN => n2136);
   U2116 : INV_X1 port map( A => REGISTERS_30_18_port, ZN => n2200);
   U2117 : INV_X1 port map( A => REGISTERS_0_18_port, ZN => n488);
   U2118 : INV_X1 port map( A => REGISTERS_4_18_port, ZN => n1816);
   U2119 : INV_X1 port map( A => REGISTERS_8_18_port, ZN => n1880);
   U2120 : INV_X1 port map( A => REGISTERS_12_18_port, ZN => n1944);
   U2121 : INV_X1 port map( A => REGISTERS_16_19_port, ZN => n2007);
   U2122 : INV_X1 port map( A => REGISTERS_20_19_port, ZN => n2071);
   U2123 : INV_X1 port map( A => REGISTERS_24_19_port, ZN => n2135);
   U2124 : INV_X1 port map( A => REGISTERS_30_19_port, ZN => n2199);
   U2125 : INV_X1 port map( A => REGISTERS_0_19_port, ZN => n487);
   U2126 : INV_X1 port map( A => REGISTERS_4_19_port, ZN => n1815);
   U2127 : INV_X1 port map( A => REGISTERS_8_19_port, ZN => n1879);
   U2128 : INV_X1 port map( A => REGISTERS_12_19_port, ZN => n1943);
   U2129 : INV_X1 port map( A => REGISTERS_16_20_port, ZN => n2006);
   U2130 : INV_X1 port map( A => REGISTERS_20_20_port, ZN => n2070);
   U2131 : INV_X1 port map( A => REGISTERS_24_20_port, ZN => n2134);
   U2132 : INV_X1 port map( A => REGISTERS_30_20_port, ZN => n2198);
   U2133 : INV_X1 port map( A => REGISTERS_0_20_port, ZN => n486);
   U2134 : INV_X1 port map( A => REGISTERS_4_20_port, ZN => n1814);
   U2135 : INV_X1 port map( A => REGISTERS_8_20_port, ZN => n1878);
   U2136 : INV_X1 port map( A => REGISTERS_12_20_port, ZN => n1942);
   U2137 : INV_X1 port map( A => REGISTERS_16_21_port, ZN => n2005);
   U2138 : INV_X1 port map( A => REGISTERS_20_21_port, ZN => n2069);
   U2139 : INV_X1 port map( A => REGISTERS_24_21_port, ZN => n2133);
   U2140 : INV_X1 port map( A => REGISTERS_30_21_port, ZN => n2197);
   U2141 : INV_X1 port map( A => REGISTERS_0_21_port, ZN => n485);
   U2142 : INV_X1 port map( A => REGISTERS_4_21_port, ZN => n1813);
   U2143 : INV_X1 port map( A => REGISTERS_8_21_port, ZN => n1877);
   U2144 : INV_X1 port map( A => REGISTERS_12_21_port, ZN => n1941);
   U2145 : INV_X1 port map( A => REGISTERS_16_22_port, ZN => n2004);
   U2146 : INV_X1 port map( A => REGISTERS_20_22_port, ZN => n2068);
   U2147 : INV_X1 port map( A => REGISTERS_24_22_port, ZN => n2132);
   U2148 : INV_X1 port map( A => REGISTERS_30_22_port, ZN => n2196);
   U2149 : INV_X1 port map( A => REGISTERS_0_22_port, ZN => n484);
   U2150 : INV_X1 port map( A => REGISTERS_4_22_port, ZN => n1812);
   U2151 : INV_X1 port map( A => REGISTERS_8_22_port, ZN => n1876);
   U2152 : INV_X1 port map( A => REGISTERS_12_22_port, ZN => n1940);
   U2153 : INV_X1 port map( A => REGISTERS_16_23_port, ZN => n2003);
   U2154 : INV_X1 port map( A => REGISTERS_20_23_port, ZN => n2067);
   U2155 : INV_X1 port map( A => REGISTERS_24_23_port, ZN => n2131);
   U2156 : INV_X1 port map( A => REGISTERS_30_23_port, ZN => n2195);
   U2157 : INV_X1 port map( A => REGISTERS_0_23_port, ZN => n483);
   U2158 : INV_X1 port map( A => REGISTERS_4_23_port, ZN => n1811);
   U2159 : INV_X1 port map( A => REGISTERS_8_23_port, ZN => n1875);
   U2160 : INV_X1 port map( A => REGISTERS_12_23_port, ZN => n1939);
   U2161 : INV_X1 port map( A => REGISTERS_16_24_port, ZN => n2002);
   U2162 : INV_X1 port map( A => REGISTERS_20_24_port, ZN => n2066);
   U2163 : INV_X1 port map( A => REGISTERS_24_24_port, ZN => n2130);
   U2164 : INV_X1 port map( A => REGISTERS_30_24_port, ZN => n2194);
   U2165 : INV_X1 port map( A => REGISTERS_0_24_port, ZN => n482);
   U2166 : INV_X1 port map( A => REGISTERS_4_24_port, ZN => n1810);
   U2167 : INV_X1 port map( A => REGISTERS_8_24_port, ZN => n1874);
   U2168 : INV_X1 port map( A => REGISTERS_12_24_port, ZN => n1938);
   U2169 : INV_X1 port map( A => REGISTERS_16_25_port, ZN => n2001);
   U2170 : INV_X1 port map( A => REGISTERS_20_25_port, ZN => n2065);
   U2171 : INV_X1 port map( A => REGISTERS_24_25_port, ZN => n2129);
   U2172 : INV_X1 port map( A => REGISTERS_30_25_port, ZN => n2193);
   U2173 : INV_X1 port map( A => REGISTERS_0_25_port, ZN => n481);
   U2174 : INV_X1 port map( A => REGISTERS_4_25_port, ZN => n1809);
   U2175 : INV_X1 port map( A => REGISTERS_8_25_port, ZN => n1873);
   U2176 : INV_X1 port map( A => REGISTERS_12_25_port, ZN => n1937);
   U2177 : INV_X1 port map( A => REGISTERS_16_26_port, ZN => n2000);
   U2178 : INV_X1 port map( A => REGISTERS_20_26_port, ZN => n2064);
   U2179 : INV_X1 port map( A => REGISTERS_24_26_port, ZN => n2128);
   U2180 : INV_X1 port map( A => REGISTERS_30_26_port, ZN => n2192);
   U2181 : INV_X1 port map( A => REGISTERS_0_26_port, ZN => n480);
   U2182 : INV_X1 port map( A => REGISTERS_4_26_port, ZN => n1808);
   U2183 : INV_X1 port map( A => REGISTERS_8_26_port, ZN => n1872);
   U2184 : INV_X1 port map( A => REGISTERS_12_26_port, ZN => n1936);
   U2185 : INV_X1 port map( A => REGISTERS_16_27_port, ZN => n1999);
   U2186 : INV_X1 port map( A => REGISTERS_20_27_port, ZN => n2063);
   U2187 : INV_X1 port map( A => REGISTERS_24_27_port, ZN => n2127);
   U2188 : INV_X1 port map( A => REGISTERS_30_27_port, ZN => n2191);
   U2189 : INV_X1 port map( A => REGISTERS_0_27_port, ZN => n479);
   U2190 : INV_X1 port map( A => REGISTERS_4_27_port, ZN => n1807);
   U2191 : INV_X1 port map( A => REGISTERS_8_27_port, ZN => n1871);
   U2192 : INV_X1 port map( A => REGISTERS_12_27_port, ZN => n1935);
   U2193 : INV_X1 port map( A => REGISTERS_16_28_port, ZN => n1998);
   U2194 : INV_X1 port map( A => REGISTERS_20_28_port, ZN => n2062);
   U2195 : INV_X1 port map( A => REGISTERS_24_28_port, ZN => n2126);
   U2196 : INV_X1 port map( A => REGISTERS_30_28_port, ZN => n2190);
   U2197 : INV_X1 port map( A => REGISTERS_0_28_port, ZN => n478);
   U2198 : INV_X1 port map( A => REGISTERS_4_28_port, ZN => n1806);
   U2199 : INV_X1 port map( A => REGISTERS_8_28_port, ZN => n1870);
   U2200 : INV_X1 port map( A => REGISTERS_12_28_port, ZN => n1934);
   U2201 : INV_X1 port map( A => REGISTERS_16_29_port, ZN => n1997);
   U2202 : INV_X1 port map( A => REGISTERS_20_29_port, ZN => n2061);
   U2203 : INV_X1 port map( A => REGISTERS_24_29_port, ZN => n2125);
   U2204 : INV_X1 port map( A => REGISTERS_30_29_port, ZN => n2189);
   U2205 : INV_X1 port map( A => REGISTERS_0_29_port, ZN => n477);
   U2206 : INV_X1 port map( A => REGISTERS_4_29_port, ZN => n1805);
   U2207 : INV_X1 port map( A => REGISTERS_8_29_port, ZN => n1869);
   U2208 : INV_X1 port map( A => REGISTERS_12_29_port, ZN => n1933);
   U2209 : INV_X1 port map( A => REGISTERS_16_30_port, ZN => n1996);
   U2210 : INV_X1 port map( A => REGISTERS_20_30_port, ZN => n2060);
   U2211 : INV_X1 port map( A => REGISTERS_24_30_port, ZN => n2124);
   U2212 : INV_X1 port map( A => REGISTERS_30_30_port, ZN => n2188);
   U2213 : INV_X1 port map( A => REGISTERS_0_30_port, ZN => n476);
   U2214 : INV_X1 port map( A => REGISTERS_4_30_port, ZN => n1804);
   U2215 : INV_X1 port map( A => REGISTERS_8_30_port, ZN => n1868);
   U2216 : INV_X1 port map( A => REGISTERS_12_30_port, ZN => n1932);
   U2217 : INV_X1 port map( A => REGISTERS_16_31_port, ZN => n1995);
   U2218 : INV_X1 port map( A => REGISTERS_20_31_port, ZN => n2059);
   U2219 : INV_X1 port map( A => REGISTERS_24_31_port, ZN => n2123);
   U2220 : INV_X1 port map( A => REGISTERS_30_31_port, ZN => n2187);
   U2221 : INV_X1 port map( A => REGISTERS_0_31_port, ZN => n475);
   U2222 : INV_X1 port map( A => REGISTERS_4_31_port, ZN => n1803);
   U2223 : INV_X1 port map( A => REGISTERS_8_31_port, ZN => n1867);
   U2224 : INV_X1 port map( A => REGISTERS_12_31_port, ZN => n1931);
   U2225 : INV_X1 port map( A => ADD_RD1(2), ZN => n2257);
   U2226 : NOR2_X1 port map( A1 => n2256, A2 => ADD_RD1(2), ZN => n1750);
   U2227 : NOR2_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(2), ZN => n1752);
   U2228 : CLKBUF_X1 port map( A => N409, Z => n196);
   U2229 : CLKBUF_X1 port map( A => N409, Z => n197);
   U2230 : CLKBUF_X1 port map( A => N409, Z => n198);
   U2231 : CLKBUF_X1 port map( A => N409, Z => n199);
   U2232 : CLKBUF_X1 port map( A => N376, Z => n200);
   U2233 : CLKBUF_X1 port map( A => N376, Z => n201);
   U2234 : CLKBUF_X1 port map( A => N376, Z => n202);
   U2235 : CLKBUF_X1 port map( A => N376, Z => n203);
   U2236 : CLKBUF_X1 port map( A => N375, Z => n204);
   U2237 : CLKBUF_X1 port map( A => N375, Z => n205);
   U2238 : CLKBUF_X1 port map( A => N375, Z => n206);
   U2239 : CLKBUF_X1 port map( A => N375, Z => n207);
   U2240 : CLKBUF_X1 port map( A => N374, Z => n208);
   U2241 : CLKBUF_X1 port map( A => N374, Z => n209);
   U2242 : CLKBUF_X1 port map( A => N374, Z => n210);
   U2243 : CLKBUF_X1 port map( A => N374, Z => n211);
   U2244 : CLKBUF_X1 port map( A => N373, Z => n212);
   U2245 : CLKBUF_X1 port map( A => N373, Z => n213);
   U2246 : CLKBUF_X1 port map( A => N373, Z => n214);
   U2247 : CLKBUF_X1 port map( A => N373, Z => n215);
   U2248 : CLKBUF_X1 port map( A => N372, Z => n216);
   U2249 : CLKBUF_X1 port map( A => N372, Z => n217);
   U2250 : CLKBUF_X1 port map( A => N372, Z => n218);
   U2251 : CLKBUF_X1 port map( A => N372, Z => n219);
   U2252 : CLKBUF_X1 port map( A => N371, Z => n220);
   U2253 : CLKBUF_X1 port map( A => N371, Z => n221);
   U2254 : CLKBUF_X1 port map( A => N371, Z => n222);
   U2255 : CLKBUF_X1 port map( A => N371, Z => n223);
   U2256 : CLKBUF_X1 port map( A => N370, Z => n224);
   U2257 : CLKBUF_X1 port map( A => N370, Z => n225);
   U2258 : CLKBUF_X1 port map( A => N370, Z => n226);
   U2259 : CLKBUF_X1 port map( A => N370, Z => n227);
   U2260 : CLKBUF_X1 port map( A => N369, Z => n228);
   U2261 : CLKBUF_X1 port map( A => N369, Z => n229);
   U2262 : CLKBUF_X1 port map( A => N369, Z => n230);
   U2263 : CLKBUF_X1 port map( A => N369, Z => n231);
   U2264 : CLKBUF_X1 port map( A => N368, Z => n232);
   U2265 : CLKBUF_X1 port map( A => N368, Z => n233);
   U2266 : CLKBUF_X1 port map( A => N368, Z => n234);
   U2267 : CLKBUF_X1 port map( A => N368, Z => n235);
   U2268 : CLKBUF_X1 port map( A => N367, Z => n236);
   U2269 : CLKBUF_X1 port map( A => N367, Z => n237);
   U2270 : CLKBUF_X1 port map( A => N367, Z => n238);
   U2271 : CLKBUF_X1 port map( A => N367, Z => n239);
   U2272 : CLKBUF_X1 port map( A => N366, Z => n240);
   U2273 : CLKBUF_X1 port map( A => N366, Z => n241);
   U2274 : CLKBUF_X1 port map( A => N366, Z => n242);
   U2275 : CLKBUF_X1 port map( A => N366, Z => n243);
   U2276 : CLKBUF_X1 port map( A => N365, Z => n244);
   U2277 : CLKBUF_X1 port map( A => N365, Z => n245);
   U2278 : CLKBUF_X1 port map( A => N365, Z => n246);
   U2279 : CLKBUF_X1 port map( A => N365, Z => n247);
   U2280 : CLKBUF_X1 port map( A => N364, Z => n248);
   U2281 : CLKBUF_X1 port map( A => N364, Z => n249);
   U2282 : CLKBUF_X1 port map( A => N364, Z => n250);
   U2283 : CLKBUF_X1 port map( A => N364, Z => n251);
   U2284 : CLKBUF_X1 port map( A => N363, Z => n252);
   U2285 : CLKBUF_X1 port map( A => N363, Z => n253);
   U2286 : CLKBUF_X1 port map( A => N363, Z => n254);
   U2287 : CLKBUF_X1 port map( A => N363, Z => n255);
   U2288 : CLKBUF_X1 port map( A => N362, Z => n256);
   U2289 : CLKBUF_X1 port map( A => N362, Z => n257);
   U2290 : CLKBUF_X1 port map( A => N362, Z => n258);
   U2291 : CLKBUF_X1 port map( A => N362, Z => n259);
   U2292 : CLKBUF_X1 port map( A => N361, Z => n260);
   U2293 : CLKBUF_X1 port map( A => N361, Z => n261);
   U2294 : CLKBUF_X1 port map( A => N361, Z => n262);
   U2295 : CLKBUF_X1 port map( A => N361, Z => n263);
   U2296 : CLKBUF_X1 port map( A => N360, Z => n264);
   U2297 : CLKBUF_X1 port map( A => N360, Z => n265);
   U2298 : CLKBUF_X1 port map( A => N360, Z => n266);
   U2299 : CLKBUF_X1 port map( A => N360, Z => n267);
   U2300 : CLKBUF_X1 port map( A => N359, Z => n268);
   U2301 : CLKBUF_X1 port map( A => N359, Z => n269);
   U2302 : CLKBUF_X1 port map( A => N359, Z => n270);
   U2303 : CLKBUF_X1 port map( A => N359, Z => n271);
   U2304 : CLKBUF_X1 port map( A => N358, Z => n272);
   U2305 : CLKBUF_X1 port map( A => N358, Z => n273);
   U2306 : CLKBUF_X1 port map( A => N358, Z => n274);
   U2307 : CLKBUF_X1 port map( A => N358, Z => n275);
   U2308 : CLKBUF_X1 port map( A => N357, Z => n276);
   U2309 : CLKBUF_X1 port map( A => N357, Z => n277);
   U2310 : CLKBUF_X1 port map( A => N357, Z => n278);
   U2311 : CLKBUF_X1 port map( A => N357, Z => n279);
   U2312 : CLKBUF_X1 port map( A => N356, Z => n280);
   U2313 : CLKBUF_X1 port map( A => N356, Z => n281);
   U2314 : CLKBUF_X1 port map( A => N356, Z => n282);
   U2315 : CLKBUF_X1 port map( A => N356, Z => n283);
   U2316 : CLKBUF_X1 port map( A => N355, Z => n284);
   U2317 : CLKBUF_X1 port map( A => N355, Z => n285);
   U2318 : CLKBUF_X1 port map( A => N355, Z => n286);
   U2319 : CLKBUF_X1 port map( A => N355, Z => n287);
   U2320 : CLKBUF_X1 port map( A => N354, Z => n288);
   U2321 : CLKBUF_X1 port map( A => N354, Z => n289);
   U2322 : CLKBUF_X1 port map( A => N354, Z => n290);
   U2323 : CLKBUF_X1 port map( A => N354, Z => n291);
   U2324 : CLKBUF_X1 port map( A => N353, Z => n292);
   U2325 : CLKBUF_X1 port map( A => N353, Z => n293);
   U2326 : CLKBUF_X1 port map( A => N353, Z => n294);
   U2327 : CLKBUF_X1 port map( A => N353, Z => n295);
   U2328 : CLKBUF_X1 port map( A => N352, Z => n296);
   U2329 : CLKBUF_X1 port map( A => N352, Z => n297);
   U2330 : CLKBUF_X1 port map( A => N352, Z => n298);
   U2331 : CLKBUF_X1 port map( A => N352, Z => n299);
   U2332 : CLKBUF_X1 port map( A => N351, Z => n300);
   U2333 : CLKBUF_X1 port map( A => N351, Z => n301);
   U2334 : CLKBUF_X1 port map( A => N351, Z => n302);
   U2335 : CLKBUF_X1 port map( A => N351, Z => n303);
   U2336 : CLKBUF_X1 port map( A => N350, Z => n304);
   U2337 : CLKBUF_X1 port map( A => N350, Z => n305);
   U2338 : CLKBUF_X1 port map( A => N350, Z => n306);
   U2339 : CLKBUF_X1 port map( A => N350, Z => n307);
   U2340 : CLKBUF_X1 port map( A => N349, Z => n308);
   U2341 : CLKBUF_X1 port map( A => N349, Z => n309);
   U2342 : CLKBUF_X1 port map( A => N349, Z => n310);
   U2343 : CLKBUF_X1 port map( A => N349, Z => n311);
   U2344 : CLKBUF_X1 port map( A => N348, Z => n312_port);
   U2345 : CLKBUF_X1 port map( A => N348, Z => n313_port);
   U2346 : CLKBUF_X1 port map( A => N348, Z => n314_port);
   U2347 : CLKBUF_X1 port map( A => N348, Z => n315_port);
   U2348 : CLKBUF_X1 port map( A => N347, Z => n316_port);
   U2349 : CLKBUF_X1 port map( A => N347, Z => n317_port);
   U2350 : CLKBUF_X1 port map( A => N347, Z => n318_port);
   U2351 : CLKBUF_X1 port map( A => N347, Z => n319_port);
   U2352 : CLKBUF_X1 port map( A => N346, Z => n320_port);
   U2353 : CLKBUF_X1 port map( A => N346, Z => n321_port);
   U2354 : CLKBUF_X1 port map( A => N346, Z => n322_port);
   U2355 : CLKBUF_X1 port map( A => N346, Z => n323_port);
   U2356 : CLKBUF_X1 port map( A => N345, Z => n324_port);
   U2357 : CLKBUF_X1 port map( A => N345, Z => n325_port);
   U2358 : CLKBUF_X1 port map( A => N345, Z => n326_port);
   U2359 : CLKBUF_X1 port map( A => N345, Z => n327_port);
   U2360 : CLKBUF_X1 port map( A => N344, Z => n331_port);
   U2361 : CLKBUF_X1 port map( A => N343, Z => n335_port);
   U2362 : CLKBUF_X1 port map( A => N342, Z => n339_port);
   U2363 : CLKBUF_X1 port map( A => N341, Z => n343_port);
   U2364 : CLKBUF_X1 port map( A => N340, Z => n347_port);
   U2365 : CLKBUF_X1 port map( A => N339, Z => n351_port);
   U2366 : CLKBUF_X1 port map( A => N338, Z => n355_port);
   U2367 : CLKBUF_X1 port map( A => N337, Z => n359_port);
   U2368 : CLKBUF_X1 port map( A => N336, Z => n363_port);
   U2369 : CLKBUF_X1 port map( A => N335, Z => n367_port);
   U2370 : CLKBUF_X1 port map( A => N334, Z => n371_port);
   U2371 : CLKBUF_X1 port map( A => N333, Z => n375_port);
   U2372 : CLKBUF_X1 port map( A => N332, Z => n379_port);
   U2373 : CLKBUF_X1 port map( A => N331, Z => n383_port);
   U2374 : CLKBUF_X1 port map( A => N330, Z => n387_port);
   U2375 : CLKBUF_X1 port map( A => N329, Z => n391_port);
   U2376 : CLKBUF_X1 port map( A => N328, Z => n395_port);
   U2377 : CLKBUF_X1 port map( A => N327, Z => n399_port);
   U2378 : CLKBUF_X1 port map( A => N326, Z => n403_port);
   U2379 : CLKBUF_X1 port map( A => N325, Z => n407_port);
   U2380 : CLKBUF_X1 port map( A => N324, Z => n411_port);
   U2381 : CLKBUF_X1 port map( A => N323, Z => n415_port);
   U2382 : CLKBUF_X1 port map( A => N322, Z => n419_port);
   U2383 : CLKBUF_X1 port map( A => N321, Z => n423_port);
   U2384 : CLKBUF_X1 port map( A => N320, Z => n427_port);
   U2385 : CLKBUF_X1 port map( A => N319, Z => n431_port);
   U2386 : CLKBUF_X1 port map( A => N318, Z => n435_port);
   U2387 : CLKBUF_X1 port map( A => N317, Z => n439_port);
   U2388 : CLKBUF_X1 port map( A => N316, Z => n443);
   U2389 : CLKBUF_X1 port map( A => N315, Z => n447);
   U2390 : CLKBUF_X1 port map( A => N314, Z => n451);
   U2391 : CLKBUF_X1 port map( A => N313, Z => n455);
   U2392 : CLKBUF_X1 port map( A => N312, Z => n456);
   U2393 : CLKBUF_X1 port map( A => N312, Z => n457);
   U2394 : CLKBUF_X1 port map( A => N312, Z => n458);
   U2395 : CLKBUF_X1 port map( A => N312, Z => n459);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity 
   stall_detection_unit_op_code_size6_func_size11_PC_reg_size32_reg_file_size32
   is

   port( opcode : in std_logic_vector (5 downto 0);  RSA, RSB, RD : in 
         std_logic_vector (4 downto 0);  FUNC : in std_logic_vector (10 downto 
         0);  EXE_RD : in std_logic_vector (4 downto 0);  NPC_in : in 
         std_logic_vector (31 downto 0);  Ld : in std_logic;  RD_inmul : in 
         std_logic_vector (4 downto 0);  flag_structHzd, flag_ismul : in 
         std_logic;  opcode_out : out std_logic_vector (5 downto 0);  RD_out : 
         out std_logic_vector (4 downto 0);  FUNC_out : out std_logic_vector 
         (10 downto 0);  NPC_out : out std_logic_vector (31 downto 0);  PC_sel 
         : out std_logic);

end 
   stall_detection_unit_op_code_size6_func_size11_PC_reg_size32_reg_file_size32
   ;

architecture SYN_Behavioral of 
   stall_detection_unit_op_code_size6_func_size11_PC_reg_size32_reg_file_size32
   is

   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component 
      stall_detection_unit_op_code_size6_func_size11_PC_reg_size32_reg_file_size32_DW01_sub_3
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  DIFF
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   component 
      stall_detection_unit_op_code_size6_func_size11_PC_reg_size32_reg_file_size32_DW01_sub_2
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  DIFF
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   component 
      stall_detection_unit_op_code_size6_func_size11_PC_reg_size32_reg_file_size32_DW01_sub_1
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  DIFF
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   component 
      stall_detection_unit_op_code_size6_func_size11_PC_reg_size32_reg_file_size32_DW01_sub_0
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  DIFF
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   signal n172, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46
      , N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, 
      N61, N62, N63, N64, N65, N104, N105, N106, N107, N108, N109, N110, N111, 
      N112, N113, N114, N115, N116, N117, N118, N119, N120, N121, N122, N123, 
      N124, N125, N126, N127, N128, N129, N130, N131, N132, N133, N134, N135, 
      N141, N142, N143, N144, N145, N146, N147, N148, N149, N150, N151, N152, 
      N153, N154, N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, 
      N165, N166, N167, N168, N169, N170, N171, N172_port, N265, N266, N267, 
      N268, N269, N270, N271, N272, N273, N274, N275, N276, N277, N278, N279, 
      N280, N281, N282, N283, N284, N285, N286, N287, N288, N289, N290, N291, 
      N292, N293, N294, N295, N296, n26, n27, n28, n30, n31, n32, PC_sel_port, 
      n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, 
      n18, n19, n20, n21, n22, n23, n24, n25, n29, n33, n34_port, n35_port, 
      n36_port, n37_port, n38_port, n39_port, n40_port, n41_port, n42_port, 
      n43_port, n44_port, n45_port, n46_port, n47_port, n48_port, n49_port, 
      n50_port, n51_port, n52_port, n53_port, n54_port, n55_port, n56_port, 
      n57_port, n58_port, n59_port, n60_port, n61_port, n62_port, n63_port, 
      n64_port, n65_port, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76
      , n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, 
      n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, 
      n104_port, n105_port, n106_port, n107_port, n108_port, n109_port, 
      n110_port, n111_port, n112_port, n113_port, n114_port, n115_port, 
      n116_port, n117_port, n118_port, n119_port, n120_port, n121_port, 
      n122_port, n123_port, n124_port, n125_port, n126_port, n127_port, 
      n128_port, n129_port, n130_port, n131_port, n132_port, n133_port, 
      n134_port, n135_port, n136, n137, n138, n139, n140, n141_port, n142_port,
      n143_port, n144_port, n145_port, n146_port, n147_port, n148_port, 
      n149_port, n150_port, n151_port, n152_port, n153_port, n154_port, 
      n155_port, n156_port, n157_port, n158_port, n159_port, n160_port, 
      n161_port, n162_port, n163_port, n164_port, n165_port, n166_port, 
      n167_port, n168_port, n169_port, n170_port, n171_port, n_1939, n_1940, 
      n_1941, n_1942 : std_logic;

begin
   FUNC_out <= ( FUNC(10), FUNC(9), FUNC(8), FUNC(7), FUNC(6), FUNC(5), FUNC(4)
      , FUNC(3), FUNC(2), FUNC(1), FUNC(0) );
   PC_sel <= PC_sel_port;
   
   n26 <= '0';
   n27 <= '1';
   n28 <= '0';
   n30 <= '0';
   n31 <= '0';
   n32 <= '0';
   sub_100_aco : 
                           stall_detection_unit_op_code_size6_func_size11_PC_reg_size32_reg_file_size32_DW01_sub_0 
                           port map( A(31) => NPC_in(31), A(30) => NPC_in(30), 
                           A(29) => NPC_in(29), A(28) => NPC_in(28), A(27) => 
                           NPC_in(27), A(26) => NPC_in(26), A(25) => NPC_in(25)
                           , A(24) => NPC_in(24), A(23) => NPC_in(23), A(22) =>
                           NPC_in(22), A(21) => NPC_in(21), A(20) => NPC_in(20)
                           , A(19) => NPC_in(19), A(18) => NPC_in(18), A(17) =>
                           NPC_in(17), A(16) => NPC_in(16), A(15) => NPC_in(15)
                           , A(14) => NPC_in(14), A(13) => NPC_in(13), A(12) =>
                           NPC_in(12), A(11) => NPC_in(11), A(10) => NPC_in(10)
                           , A(9) => NPC_in(9), A(8) => NPC_in(8), A(7) => 
                           NPC_in(7), A(6) => NPC_in(6), A(5) => NPC_in(5), 
                           A(4) => NPC_in(4), A(3) => NPC_in(3), A(2) => 
                           NPC_in(2), A(1) => NPC_in(1), A(0) => NPC_in(0), 
                           B(31) => n28, B(30) => n28, B(29) => n28, B(28) => 
                           n28, B(27) => n28, B(26) => n28, B(25) => n28, B(24)
                           => n28, B(23) => n28, B(22) => n28, B(21) => n28, 
                           B(20) => n28, B(19) => n28, B(18) => n28, B(17) => 
                           n28, B(16) => n28, B(15) => n28, B(14) => n28, B(13)
                           => n28, B(12) => n28, B(11) => n28, B(10) => n28, 
                           B(9) => n28, B(8) => n28, B(7) => n28, B(6) => n28, 
                           B(5) => n28, B(4) => n28, B(3) => n28, B(2) => 
                           flag_structHzd, B(1) => n26, B(0) => n26, CI => n28,
                           DIFF(31) => N296, DIFF(30) => N295, DIFF(29) => N294
                           , DIFF(28) => N293, DIFF(27) => N292, DIFF(26) => 
                           N291, DIFF(25) => N290, DIFF(24) => N289, DIFF(23) 
                           => N288, DIFF(22) => N287, DIFF(21) => N286, 
                           DIFF(20) => N285, DIFF(19) => N284, DIFF(18) => N283
                           , DIFF(17) => N282, DIFF(16) => N281, DIFF(15) => 
                           N280, DIFF(14) => N279, DIFF(13) => N278, DIFF(12) 
                           => N277, DIFF(11) => N276, DIFF(10) => N275, DIFF(9)
                           => N274, DIFF(8) => N273, DIFF(7) => N272, DIFF(6) 
                           => N271, DIFF(5) => N270, DIFF(4) => N269, DIFF(3) 
                           => N268, DIFF(2) => N267, DIFF(1) => N266, DIFF(0) 
                           => N265, CO => n_1939);
   sub_73_aco : 
                           stall_detection_unit_op_code_size6_func_size11_PC_reg_size32_reg_file_size32_DW01_sub_1 
                           port map( A(31) => NPC_in(31), A(30) => NPC_in(30), 
                           A(29) => NPC_in(29), A(28) => NPC_in(28), A(27) => 
                           NPC_in(27), A(26) => NPC_in(26), A(25) => NPC_in(25)
                           , A(24) => NPC_in(24), A(23) => NPC_in(23), A(22) =>
                           NPC_in(22), A(21) => NPC_in(21), A(20) => NPC_in(20)
                           , A(19) => NPC_in(19), A(18) => NPC_in(18), A(17) =>
                           NPC_in(17), A(16) => NPC_in(16), A(15) => NPC_in(15)
                           , A(14) => NPC_in(14), A(13) => NPC_in(13), A(12) =>
                           NPC_in(12), A(11) => NPC_in(11), A(10) => NPC_in(10)
                           , A(9) => NPC_in(9), A(8) => NPC_in(8), A(7) => 
                           NPC_in(7), A(6) => NPC_in(6), A(5) => NPC_in(5), 
                           A(4) => NPC_in(4), A(3) => NPC_in(3), A(2) => 
                           NPC_in(2), A(1) => NPC_in(1), A(0) => NPC_in(0), 
                           B(31) => n30, B(30) => n30, B(29) => n30, B(28) => 
                           n30, B(27) => n30, B(26) => n30, B(25) => n30, B(24)
                           => n30, B(23) => n30, B(22) => n30, B(21) => n30, 
                           B(20) => n30, B(19) => n30, B(18) => n30, B(17) => 
                           n30, B(16) => n30, B(15) => n30, B(14) => n30, B(13)
                           => n30, B(12) => n30, B(11) => n30, B(10) => n30, 
                           B(9) => n30, B(8) => n30, B(7) => n30, B(6) => n30, 
                           B(5) => n30, B(4) => n30, B(3) => n30, B(2) => 
                           n171_port, B(1) => n26, B(0) => n26, CI => n30, 
                           DIFF(31) => N135, DIFF(30) => N134, DIFF(29) => N133
                           , DIFF(28) => N132, DIFF(27) => N131, DIFF(26) => 
                           N130, DIFF(25) => N129, DIFF(24) => N128, DIFF(23) 
                           => N127, DIFF(22) => N126, DIFF(21) => N125, 
                           DIFF(20) => N124, DIFF(19) => N123, DIFF(18) => N122
                           , DIFF(17) => N121, DIFF(16) => N120, DIFF(15) => 
                           N119, DIFF(14) => N118, DIFF(13) => N117, DIFF(12) 
                           => N116, DIFF(11) => N115, DIFF(10) => N114, DIFF(9)
                           => N113, DIFF(8) => N112, DIFF(7) => N111, DIFF(6) 
                           => N110, DIFF(5) => N109, DIFF(4) => N108, DIFF(3) 
                           => N107, DIFF(2) => N106, DIFF(1) => N105, DIFF(0) 
                           => N104, CO => n_1940);
   sub_60_aco : 
                           stall_detection_unit_op_code_size6_func_size11_PC_reg_size32_reg_file_size32_DW01_sub_2 
                           port map( A(31) => NPC_in(31), A(30) => NPC_in(30), 
                           A(29) => NPC_in(29), A(28) => NPC_in(28), A(27) => 
                           NPC_in(27), A(26) => NPC_in(26), A(25) => NPC_in(25)
                           , A(24) => NPC_in(24), A(23) => NPC_in(23), A(22) =>
                           NPC_in(22), A(21) => NPC_in(21), A(20) => NPC_in(20)
                           , A(19) => NPC_in(19), A(18) => NPC_in(18), A(17) =>
                           NPC_in(17), A(16) => NPC_in(16), A(15) => NPC_in(15)
                           , A(14) => NPC_in(14), A(13) => NPC_in(13), A(12) =>
                           NPC_in(12), A(11) => NPC_in(11), A(10) => NPC_in(10)
                           , A(9) => NPC_in(9), A(8) => NPC_in(8), A(7) => 
                           NPC_in(7), A(6) => NPC_in(6), A(5) => NPC_in(5), 
                           A(4) => NPC_in(4), A(3) => NPC_in(3), A(2) => 
                           NPC_in(2), A(1) => NPC_in(1), A(0) => NPC_in(0), 
                           B(31) => n31, B(30) => n31, B(29) => n31, B(28) => 
                           n31, B(27) => n31, B(26) => n31, B(25) => n31, B(24)
                           => n31, B(23) => n31, B(22) => n31, B(21) => n31, 
                           B(20) => n31, B(19) => n31, B(18) => n31, B(17) => 
                           n31, B(16) => n31, B(15) => n31, B(14) => n31, B(13)
                           => n31, B(12) => n31, B(11) => n31, B(10) => n31, 
                           B(9) => n31, B(8) => n31, B(7) => n31, B(6) => n31, 
                           B(5) => n31, B(4) => n31, B(3) => n31, B(2) => 
                           n170_port, B(1) => n26, B(0) => n26, CI => n31, 
                           DIFF(31) => N65, DIFF(30) => N64, DIFF(29) => N63, 
                           DIFF(28) => N62, DIFF(27) => N61, DIFF(26) => N60, 
                           DIFF(25) => N59, DIFF(24) => N58, DIFF(23) => N57, 
                           DIFF(22) => N56, DIFF(21) => N55, DIFF(20) => N54, 
                           DIFF(19) => N53, DIFF(18) => N52, DIFF(17) => N51, 
                           DIFF(16) => N50, DIFF(15) => N49, DIFF(14) => N48, 
                           DIFF(13) => N47, DIFF(12) => N46, DIFF(11) => N45, 
                           DIFF(10) => N44, DIFF(9) => N43, DIFF(8) => N42, 
                           DIFF(7) => N41, DIFF(6) => N40, DIFF(5) => N39, 
                           DIFF(4) => N38, DIFF(3) => N37, DIFF(2) => N36, 
                           DIFF(1) => N35, DIFF(0) => N34, CO => n_1941);
   r107 : 
                           stall_detection_unit_op_code_size6_func_size11_PC_reg_size32_reg_file_size32_DW01_sub_3 
                           port map( A(31) => NPC_in(31), A(30) => NPC_in(30), 
                           A(29) => NPC_in(29), A(28) => NPC_in(28), A(27) => 
                           NPC_in(27), A(26) => NPC_in(26), A(25) => NPC_in(25)
                           , A(24) => NPC_in(24), A(23) => NPC_in(23), A(22) =>
                           NPC_in(22), A(21) => NPC_in(21), A(20) => NPC_in(20)
                           , A(19) => NPC_in(19), A(18) => NPC_in(18), A(17) =>
                           NPC_in(17), A(16) => NPC_in(16), A(15) => NPC_in(15)
                           , A(14) => NPC_in(14), A(13) => NPC_in(13), A(12) =>
                           NPC_in(12), A(11) => NPC_in(11), A(10) => NPC_in(10)
                           , A(9) => NPC_in(9), A(8) => NPC_in(8), A(7) => 
                           NPC_in(7), A(6) => NPC_in(6), A(5) => NPC_in(5), 
                           A(4) => NPC_in(4), A(3) => NPC_in(3), A(2) => 
                           NPC_in(2), A(1) => NPC_in(1), A(0) => NPC_in(0), 
                           B(31) => n32, B(30) => n32, B(29) => n32, B(28) => 
                           n32, B(27) => n32, B(26) => n32, B(25) => n32, B(24)
                           => n32, B(23) => n32, B(22) => n32, B(21) => n32, 
                           B(20) => n32, B(19) => n32, B(18) => n32, B(17) => 
                           n32, B(16) => n32, B(15) => n32, B(14) => n32, B(13)
                           => n32, B(12) => n32, B(11) => n32, B(10) => n32, 
                           B(9) => n32, B(8) => n32, B(7) => n32, B(6) => n32, 
                           B(5) => n32, B(4) => n32, B(3) => n32, B(2) => n27, 
                           B(1) => n26, B(0) => n26, CI => n32, DIFF(31) => 
                           N172_port, DIFF(30) => N171, DIFF(29) => N170, 
                           DIFF(28) => N169, DIFF(27) => N168, DIFF(26) => N167
                           , DIFF(25) => N166, DIFF(24) => N165, DIFF(23) => 
                           N164, DIFF(22) => N163, DIFF(21) => N162, DIFF(20) 
                           => N161, DIFF(19) => N160, DIFF(18) => N159, 
                           DIFF(17) => N158, DIFF(16) => N157, DIFF(15) => N156
                           , DIFF(14) => N155, DIFF(13) => N154, DIFF(12) => 
                           N153, DIFF(11) => N152, DIFF(10) => N151, DIFF(9) =>
                           N150, DIFF(8) => N149, DIFF(7) => N148, DIFF(6) => 
                           N147, DIFF(5) => N146, DIFF(4) => N145, DIFF(3) => 
                           N144, DIFF(2) => N143, DIFF(1) => N142, DIFF(0) => 
                           N141, CO => n_1942);
   U6 : NOR2_X2 port map( A1 => PC_sel_port, A2 => n25, ZN => opcode_out(3));
   U9 : NOR2_X2 port map( A1 => PC_sel_port, A2 => n22, ZN => opcode_out(5));
   U10 : BUF_X1 port map( A => n172, Z => PC_sel_port);
   U11 : BUF_X1 port map( A => n16, Z => n18);
   U12 : BUF_X1 port map( A => n19, Z => n21);
   U13 : BUF_X1 port map( A => n57_port, Z => n15);
   U14 : BUF_X1 port map( A => n4, Z => n6);
   U15 : BUF_X1 port map( A => n4, Z => n7);
   U16 : BUF_X1 port map( A => n5, Z => n9);
   U17 : BUF_X1 port map( A => n57_port, Z => n13);
   U18 : BUF_X1 port map( A => n5, Z => n8);
   U20 : BUF_X1 port map( A => n57_port, Z => n14);
   U21 : BUF_X1 port map( A => n42_port, Z => n10);
   U22 : BUF_X1 port map( A => n42_port, Z => n11);
   U23 : BUF_X1 port map( A => n41_port, Z => n4);
   U24 : BUF_X1 port map( A => n41_port, Z => n5);
   U25 : BUF_X1 port map( A => n42_port, Z => n12);
   U26 : NOR2_X1 port map( A1 => n23, A2 => n9, ZN => n172);
   U27 : BUF_X1 port map( A => n58_port, Z => n16);
   U28 : CLKBUF_X1 port map( A => n16, Z => n17);
   U29 : BUF_X1 port map( A => n59_port, Z => n19);
   U30 : CLKBUF_X1 port map( A => n19, Z => n20);
   U31 : OAI33_X1 port map( A1 => n155_port, A2 => n156_port, A3 => n157_port, 
                           B1 => n158_port, B2 => n159_port, B3 => n160_port, 
                           ZN => n2);
   U32 : CLKBUF_X1 port map( A => n23, Z => n3);
   U33 : NAND2_X1 port map( A1 => n3, A2 => n24, ZN => opcode_out(4));
   U34 : INV_X1 port map( A => opcode(4), ZN => n24);
   U35 : NAND2_X1 port map( A1 => n3, A2 => n29, ZN => opcode_out(2));
   U36 : INV_X1 port map( A => opcode(2), ZN => n29);
   U37 : NOR2_X1 port map( A1 => PC_sel_port, A2 => n33, ZN => opcode_out(1));
   U38 : NAND2_X1 port map( A1 => n3, A2 => n34_port, ZN => opcode_out(0));
   U39 : INV_X1 port map( A => opcode(0), ZN => n34_port);
   U40 : NOR2_X1 port map( A1 => n35_port, A2 => n36_port, ZN => RD_out(4));
   U41 : INV_X1 port map( A => RD(4), ZN => n36_port);
   U42 : NOR2_X1 port map( A1 => n35_port, A2 => n37_port, ZN => RD_out(3));
   U43 : NOR2_X1 port map( A1 => n35_port, A2 => n38_port, ZN => RD_out(2));
   U44 : INV_X1 port map( A => RD(2), ZN => n38_port);
   U45 : NOR2_X1 port map( A1 => n35_port, A2 => n39_port, ZN => RD_out(1));
   U46 : NOR2_X1 port map( A1 => n35_port, A2 => n40_port, ZN => RD_out(0));
   U47 : NOR3_X1 port map( A1 => n6, A2 => n10, A3 => n43_port, ZN => n35_port)
                           ;
   U48 : INV_X1 port map( A => n44_port, ZN => n43_port);
   U49 : MUX2_X1 port map( A => n45_port, B => n170_port, S => Ld, Z => 
                           n44_port);
   U50 : AOI222_X1 port map( A1 => n171_port, A2 => n10, B1 => n45_port, B2 => 
                           n46_port, C1 => n170_port, C2 => Ld, ZN => n23);
   U51 : INV_X1 port map( A => n47_port, ZN => n46_port);
   U52 : OR2_X1 port map( A1 => flag_structHzd, A2 => n48_port, ZN => n45_port)
                           ;
   U53 : NOR2_X1 port map( A1 => n49_port, A2 => n50_port, ZN => n171_port);
   U54 : AND4_X1 port map( A1 => n51_port, A2 => n52_port, A3 => n53_port, A4 
                           => n54_port, ZN => n50_port);
   U55 : NOR2_X1 port map( A1 => RSA(1), A2 => RSA(0), ZN => n54_port);
   U56 : INV_X1 port map( A => RSA(2), ZN => n53_port);
   U57 : INV_X1 port map( A => RSA(4), ZN => n52_port);
   U58 : NAND2_X1 port map( A1 => n55_port, A2 => n56_port, ZN => NPC_out(9));
   U59 : AOI222_X1 port map( A1 => N43, A2 => n15, B1 => N150, B2 => n18, C1 =>
                           N274, C2 => n21, ZN => n56_port);
   U60 : AOI22_X1 port map( A1 => NPC_in(9), A2 => n6, B1 => N113, B2 => n10, 
                           ZN => n55_port);
   U61 : NAND2_X1 port map( A1 => n60_port, A2 => n61_port, ZN => NPC_out(8));
   U62 : AOI222_X1 port map( A1 => N42, A2 => n15, B1 => N149, B2 => n18, C1 =>
                           N273, C2 => n21, ZN => n61_port);
   U63 : AOI22_X1 port map( A1 => NPC_in(8), A2 => n6, B1 => N112, B2 => n10, 
                           ZN => n60_port);
   U64 : NAND2_X1 port map( A1 => n62_port, A2 => n63_port, ZN => NPC_out(7));
   U65 : AOI222_X1 port map( A1 => N41, A2 => n15, B1 => N148, B2 => n18, C1 =>
                           N272, C2 => n21, ZN => n63_port);
   U66 : AOI22_X1 port map( A1 => NPC_in(7), A2 => n6, B1 => N111, B2 => n10, 
                           ZN => n62_port);
   U67 : NAND2_X1 port map( A1 => n64_port, A2 => n65_port, ZN => NPC_out(6));
   U68 : AOI222_X1 port map( A1 => N40, A2 => n15, B1 => N147, B2 => n18, C1 =>
                           N271, C2 => n21, ZN => n65_port);
   U69 : AOI22_X1 port map( A1 => NPC_in(6), A2 => n6, B1 => N110, B2 => n10, 
                           ZN => n64_port);
   U70 : NAND2_X1 port map( A1 => n66, A2 => n67, ZN => NPC_out(5));
   U71 : AOI222_X1 port map( A1 => N39, A2 => n15, B1 => N146, B2 => n17, C1 =>
                           N270, C2 => n20, ZN => n67);
   U72 : AOI22_X1 port map( A1 => NPC_in(5), A2 => n6, B1 => N109, B2 => n10, 
                           ZN => n66);
   U73 : NAND2_X1 port map( A1 => n68, A2 => n69, ZN => NPC_out(4));
   U74 : AOI222_X1 port map( A1 => N38, A2 => n15, B1 => N145, B2 => n16, C1 =>
                           N269, C2 => n19, ZN => n69);
   U75 : AOI22_X1 port map( A1 => NPC_in(4), A2 => n6, B1 => N108, B2 => n10, 
                           ZN => n68);
   U76 : NAND2_X1 port map( A1 => n70, A2 => n71, ZN => NPC_out(3));
   U77 : AOI222_X1 port map( A1 => N37, A2 => n15, B1 => N144, B2 => n58_port, 
                           C1 => N268, C2 => n59_port, ZN => n71);
   U78 : AOI22_X1 port map( A1 => NPC_in(3), A2 => n7, B1 => N107, B2 => n11, 
                           ZN => n70);
   U79 : NAND2_X1 port map( A1 => n72, A2 => n73, ZN => NPC_out(31));
   U80 : AOI222_X1 port map( A1 => N65, A2 => n15, B1 => N172_port, B2 => n18, 
                           C1 => N296, C2 => n21, ZN => n73);
   U81 : AOI22_X1 port map( A1 => NPC_in(31), A2 => n6, B1 => N135, B2 => n10, 
                           ZN => n72);
   U82 : NAND2_X1 port map( A1 => n74, A2 => n75, ZN => NPC_out(30));
   U83 : AOI222_X1 port map( A1 => N64, A2 => n15, B1 => N171, B2 => n18, C1 =>
                           N295, C2 => n21, ZN => n75);
   U84 : AOI22_X1 port map( A1 => NPC_in(30), A2 => n6, B1 => N134, B2 => n10, 
                           ZN => n74);
   U85 : NAND2_X1 port map( A1 => n76, A2 => n77, ZN => NPC_out(2));
   U86 : AOI222_X1 port map( A1 => N36, A2 => n15, B1 => N143, B2 => n58_port, 
                           C1 => N267, C2 => n59_port, ZN => n77);
   U87 : AOI22_X1 port map( A1 => NPC_in(2), A2 => n6, B1 => N106, B2 => n11, 
                           ZN => n76);
   U88 : NAND2_X1 port map( A1 => n78, A2 => n79, ZN => NPC_out(29));
   U89 : AOI222_X1 port map( A1 => N63, A2 => n14, B1 => N170, B2 => n18, C1 =>
                           N294, C2 => n21, ZN => n79);
   U90 : AOI22_X1 port map( A1 => NPC_in(29), A2 => n7, B1 => N133, B2 => n11, 
                           ZN => n78);
   U91 : NAND2_X1 port map( A1 => n80, A2 => n81, ZN => NPC_out(28));
   U92 : AOI222_X1 port map( A1 => N62, A2 => n14, B1 => N169, B2 => n18, C1 =>
                           N293, C2 => n21, ZN => n81);
   U93 : AOI22_X1 port map( A1 => NPC_in(28), A2 => n7, B1 => N132, B2 => n11, 
                           ZN => n80);
   U94 : NAND2_X1 port map( A1 => n82, A2 => n83, ZN => NPC_out(27));
   U95 : AOI222_X1 port map( A1 => N61, A2 => n14, B1 => N168, B2 => n18, C1 =>
                           N292, C2 => n21, ZN => n83);
   U96 : AOI22_X1 port map( A1 => NPC_in(27), A2 => n7, B1 => N131, B2 => n11, 
                           ZN => n82);
   U97 : NAND2_X1 port map( A1 => n84, A2 => n85, ZN => NPC_out(26));
   U98 : AOI222_X1 port map( A1 => N60, A2 => n14, B1 => N167, B2 => n18, C1 =>
                           N291, C2 => n21, ZN => n85);
   U99 : AOI22_X1 port map( A1 => NPC_in(26), A2 => n7, B1 => N130, B2 => n11, 
                           ZN => n84);
   U100 : NAND2_X1 port map( A1 => n86, A2 => n87, ZN => NPC_out(25));
   U101 : AOI222_X1 port map( A1 => N59, A2 => n14, B1 => N166, B2 => n18, C1 
                           => N290, C2 => n21, ZN => n87);
   U102 : AOI22_X1 port map( A1 => NPC_in(25), A2 => n7, B1 => N129, B2 => n11,
                           ZN => n86);
   U103 : NAND2_X1 port map( A1 => n88, A2 => n89, ZN => NPC_out(24));
   U104 : AOI222_X1 port map( A1 => N58, A2 => n14, B1 => N165, B2 => n18, C1 
                           => N289, C2 => n21, ZN => n89);
   U105 : AOI22_X1 port map( A1 => NPC_in(24), A2 => n7, B1 => N128, B2 => n11,
                           ZN => n88);
   U106 : NAND2_X1 port map( A1 => n90, A2 => n91, ZN => NPC_out(23));
   U107 : AOI222_X1 port map( A1 => N57, A2 => n14, B1 => N164, B2 => n18, C1 
                           => N288, C2 => n21, ZN => n91);
   U108 : AOI22_X1 port map( A1 => NPC_in(23), A2 => n7, B1 => N127, B2 => n11,
                           ZN => n90);
   U109 : NAND2_X1 port map( A1 => n92, A2 => n93, ZN => NPC_out(22));
   U110 : AOI222_X1 port map( A1 => N56, A2 => n14, B1 => N163, B2 => n18, C1 
                           => N287, C2 => n21, ZN => n93);
   U111 : AOI22_X1 port map( A1 => NPC_in(22), A2 => n7, B1 => N126, B2 => n11,
                           ZN => n92);
   U112 : NAND2_X1 port map( A1 => n94, A2 => n95, ZN => NPC_out(21));
   U113 : AOI222_X1 port map( A1 => N55, A2 => n14, B1 => N162, B2 => n18, C1 
                           => N286, C2 => n21, ZN => n95);
   U114 : AOI22_X1 port map( A1 => NPC_in(21), A2 => n7, B1 => N125, B2 => n11,
                           ZN => n94);
   U115 : NAND2_X1 port map( A1 => n96, A2 => n97, ZN => NPC_out(20));
   U116 : AOI222_X1 port map( A1 => N54, A2 => n14, B1 => N161, B2 => n18, C1 
                           => N285, C2 => n21, ZN => n97);
   U117 : AOI22_X1 port map( A1 => NPC_in(20), A2 => n7, B1 => N124, B2 => n12,
                           ZN => n96);
   U118 : NAND2_X1 port map( A1 => n98, A2 => n99, ZN => NPC_out(1));
   U119 : AOI222_X1 port map( A1 => N35, A2 => n14, B1 => N142, B2 => n18, C1 
                           => N266, C2 => n21, ZN => n99);
   U120 : AOI22_X1 port map( A1 => NPC_in(1), A2 => n8, B1 => N105, B2 => n12, 
                           ZN => n98);
   U121 : NAND2_X1 port map( A1 => n100, A2 => n101, ZN => NPC_out(19));
   U122 : AOI222_X1 port map( A1 => N53, A2 => n13, B1 => N160, B2 => n17, C1 
                           => N284, C2 => n20, ZN => n101);
   U123 : AOI22_X1 port map( A1 => NPC_in(19), A2 => n8, B1 => N123, B2 => n12,
                           ZN => n100);
   U124 : NAND2_X1 port map( A1 => n102, A2 => n103, ZN => NPC_out(18));
   U125 : AOI222_X1 port map( A1 => N52, A2 => n13, B1 => N159, B2 => n17, C1 
                           => N283, C2 => n20, ZN => n103);
   U126 : AOI22_X1 port map( A1 => NPC_in(18), A2 => n8, B1 => N122, B2 => n12,
                           ZN => n102);
   U127 : NAND2_X1 port map( A1 => n104_port, A2 => n105_port, ZN => 
                           NPC_out(17));
   U128 : AOI222_X1 port map( A1 => N51, A2 => n13, B1 => N158, B2 => n17, C1 
                           => N282, C2 => n20, ZN => n105_port);
   U129 : AOI22_X1 port map( A1 => NPC_in(17), A2 => n8, B1 => N121, B2 => n12,
                           ZN => n104_port);
   U130 : NAND2_X1 port map( A1 => n106_port, A2 => n107_port, ZN => 
                           NPC_out(16));
   U131 : AOI222_X1 port map( A1 => N50, A2 => n13, B1 => N157, B2 => n17, C1 
                           => N281, C2 => n20, ZN => n107_port);
   U132 : AOI22_X1 port map( A1 => NPC_in(16), A2 => n8, B1 => N120, B2 => n12,
                           ZN => n106_port);
   U133 : NAND2_X1 port map( A1 => n108_port, A2 => n109_port, ZN => 
                           NPC_out(15));
   U134 : AOI222_X1 port map( A1 => N49, A2 => n13, B1 => N156, B2 => n17, C1 
                           => N280, C2 => n20, ZN => n109_port);
   U135 : AOI22_X1 port map( A1 => NPC_in(15), A2 => n8, B1 => N119, B2 => n12,
                           ZN => n108_port);
   U136 : NAND2_X1 port map( A1 => n110_port, A2 => n111_port, ZN => 
                           NPC_out(14));
   U137 : AOI222_X1 port map( A1 => N48, A2 => n13, B1 => N155, B2 => n17, C1 
                           => N279, C2 => n20, ZN => n111_port);
   U138 : AOI22_X1 port map( A1 => NPC_in(14), A2 => n8, B1 => N118, B2 => n12,
                           ZN => n110_port);
   U139 : NAND2_X1 port map( A1 => n112_port, A2 => n113_port, ZN => 
                           NPC_out(13));
   U140 : AOI222_X1 port map( A1 => N47, A2 => n13, B1 => N154, B2 => n17, C1 
                           => N278, C2 => n20, ZN => n113_port);
   U141 : AOI22_X1 port map( A1 => NPC_in(13), A2 => n8, B1 => N117, B2 => n12,
                           ZN => n112_port);
   U142 : NAND2_X1 port map( A1 => n114_port, A2 => n115_port, ZN => 
                           NPC_out(12));
   U143 : AOI222_X1 port map( A1 => N46, A2 => n13, B1 => N153, B2 => n17, C1 
                           => N277, C2 => n20, ZN => n115_port);
   U144 : AOI22_X1 port map( A1 => NPC_in(12), A2 => n8, B1 => N116, B2 => n12,
                           ZN => n114_port);
   U145 : NAND2_X1 port map( A1 => n116_port, A2 => n117_port, ZN => 
                           NPC_out(11));
   U146 : AOI222_X1 port map( A1 => N45, A2 => n13, B1 => N152, B2 => n17, C1 
                           => N276, C2 => n20, ZN => n117_port);
   U147 : AOI22_X1 port map( A1 => NPC_in(11), A2 => n8, B1 => N115, B2 => n12,
                           ZN => n116_port);
   U148 : NAND2_X1 port map( A1 => n118_port, A2 => n119_port, ZN => 
                           NPC_out(10));
   U149 : AOI222_X1 port map( A1 => N44, A2 => n13, B1 => N151, B2 => n17, C1 
                           => N275, C2 => n20, ZN => n119_port);
   U150 : AOI22_X1 port map( A1 => NPC_in(10), A2 => n8, B1 => N114, B2 => n12,
                           ZN => n118_port);
   U151 : NAND2_X1 port map( A1 => n120_port, A2 => n121_port, ZN => NPC_out(0)
                           );
   U152 : AOI222_X1 port map( A1 => N34, A2 => n13, B1 => N141, B2 => n17, C1 
                           => N265, C2 => n20, ZN => n121_port);
   U153 : NOR3_X1 port map( A1 => n48_port, A2 => n9, A3 => n47_port, ZN => 
                           n59_port);
   U154 : NOR3_X1 port map( A1 => n122_port, A2 => n9, A3 => n47_port, ZN => 
                           n58_port);
   U155 : NAND2_X1 port map( A1 => n123_port, A2 => n124_port, ZN => n47_port);
   U156 : INV_X1 port map( A => n48_port, ZN => n122_port);
   U157 : NAND2_X1 port map( A1 => n125_port, A2 => n126_port, ZN => n48_port);
   U158 : OAI21_X1 port map( B1 => n170_port, B2 => n2, A => flag_ismul, ZN => 
                           n126_port);
   U159 : NAND2_X1 port map( A1 => n49_port, A2 => n127_port, ZN => n170_port);
   U160 : NAND4_X1 port map( A1 => n131_port, A2 => n129_port, A3 => n130_port,
                           A4 => n128_port, ZN => n49_port);
   U161 : NOR2_X1 port map( A1 => n133_port, A2 => n132_port, ZN => n131_port);
   U162 : XOR2_X1 port map( A => RSA(4), B => EXE_RD(4), Z => n133_port);
   U163 : XOR2_X1 port map( A => RSA(2), B => EXE_RD(2), Z => n132_port);
   U164 : XNOR2_X1 port map( A => EXE_RD(0), B => RSA(0), ZN => n130_port);
   U165 : XNOR2_X1 port map( A => EXE_RD(1), B => RSA(1), ZN => n129_port);
   U166 : XOR2_X1 port map( A => EXE_RD(3), B => n51_port, Z => n128_port);
   U167 : NAND4_X1 port map( A1 => n134_port, A2 => n135_port, A3 => n136, A4 
                           => n137, ZN => n127_port);
   U168 : NOR2_X1 port map( A1 => n138, A2 => n139, ZN => n137);
   U169 : XOR2_X1 port map( A => RSB(4), B => EXE_RD(4), Z => n139);
   U170 : XOR2_X1 port map( A => RSB(3), B => EXE_RD(3), Z => n138);
   U171 : XNOR2_X1 port map( A => EXE_RD(1), B => RSB(1), ZN => n136);
   U172 : XNOR2_X1 port map( A => EXE_RD(2), B => RSB(2), ZN => n135_port);
   U173 : XNOR2_X1 port map( A => EXE_RD(0), B => RSB(0), ZN => n134_port);
   U174 : OAI21_X1 port map( B1 => n2, B2 => n140, A => n141_port, ZN => 
                           n125_port);
   U175 : OR4_X1 port map( A1 => RD_inmul(3), A2 => RD_inmul(4), A3 => 
                           RD_inmul(2), A4 => n142_port, ZN => n141_port);
   U176 : OR2_X1 port map( A1 => RD_inmul(1), A2 => RD_inmul(0), ZN => 
                           n142_port);
   U177 : OAI33_X1 port map( A1 => n143_port, A2 => n144_port, A3 => n145_port,
                           B1 => n146_port, B2 => n147_port, B3 => n148_port, 
                           ZN => n140);
   U178 : XOR2_X1 port map( A => RSA(4), B => RD_inmul(4), Z => n148_port);
   U179 : XOR2_X1 port map( A => RSA(2), B => RD_inmul(2), Z => n147_port);
   U180 : NAND3_X1 port map( A1 => n149_port, A2 => n150_port, A3 => n151_port,
                           ZN => n146_port);
   U181 : XNOR2_X1 port map( A => RSA(0), B => RD_inmul(0), ZN => n151_port);
   U182 : XNOR2_X1 port map( A => RSA(1), B => RD_inmul(1), ZN => n150_port);
   U183 : XOR2_X1 port map( A => n51_port, B => RD_inmul(3), Z => n149_port);
   U184 : INV_X1 port map( A => RSA(3), ZN => n51_port);
   U185 : XOR2_X1 port map( A => RSB(4), B => RD_inmul(4), Z => n145_port);
   U186 : XOR2_X1 port map( A => RSB(3), B => RD_inmul(3), Z => n144_port);
   U187 : NAND3_X1 port map( A1 => n152_port, A2 => n153_port, A3 => n154_port,
                           ZN => n143_port);
   U188 : XNOR2_X1 port map( A => RSB(1), B => RD_inmul(1), ZN => n154_port);
   U189 : XNOR2_X1 port map( A => RSB(2), B => RD_inmul(2), ZN => n153_port);
   U190 : XNOR2_X1 port map( A => RSB(0), B => RD_inmul(0), ZN => n152_port);
   U191 : XOR2_X1 port map( A => RD_inmul(4), B => RD(4), Z => n160_port);
   U192 : XOR2_X1 port map( A => RD_inmul(2), B => RD(2), Z => n159_port);
   U193 : NAND3_X1 port map( A1 => n161_port, A2 => n162_port, A3 => n163_port,
                           ZN => n158_port);
   U194 : XOR2_X1 port map( A => n40_port, B => RD_inmul(0), Z => n163_port);
   U195 : XOR2_X1 port map( A => n39_port, B => RD_inmul(1), Z => n162_port);
   U196 : XOR2_X1 port map( A => n37_port, B => RD_inmul(3), Z => n161_port);
   U197 : XOR2_X1 port map( A => RD(4), B => EXE_RD(4), Z => n157_port);
   U198 : XOR2_X1 port map( A => RD(2), B => EXE_RD(2), Z => n156_port);
   U199 : NAND3_X1 port map( A1 => n164_port, A2 => n165_port, A3 => n166_port,
                           ZN => n155_port);
   U200 : XOR2_X1 port map( A => n40_port, B => EXE_RD(0), Z => n166_port);
   U201 : INV_X1 port map( A => RD(0), ZN => n40_port);
   U202 : XOR2_X1 port map( A => n39_port, B => EXE_RD(1), Z => n165_port);
   U203 : INV_X1 port map( A => RD(1), ZN => n39_port);
   U204 : XOR2_X1 port map( A => EXE_RD(3), B => n37_port, Z => n164_port);
   U205 : INV_X1 port map( A => RD(3), ZN => n37_port);
   U206 : NOR2_X1 port map( A1 => n124_port, A2 => n9, ZN => n57_port);
   U207 : INV_X1 port map( A => Ld, ZN => n124_port);
   U208 : AOI22_X1 port map( A1 => NPC_in(0), A2 => n6, B1 => N104, B2 => n10, 
                           ZN => n120_port);
   U209 : NOR2_X1 port map( A1 => n123_port, A2 => Ld, ZN => n42_port);
   U210 : NAND4_X1 port map( A1 => n167_port, A2 => n168_port, A3 => n25, A4 =>
                           n22, ZN => n123_port);
   U211 : INV_X1 port map( A => opcode(5), ZN => n22);
   U212 : INV_X1 port map( A => opcode(3), ZN => n25);
   U213 : NAND2_X1 port map( A1 => opcode(4), A2 => n33, ZN => n168_port);
   U214 : MUX2_X1 port map( A => opcode(4), B => n33, S => opcode(2), Z => 
                           n167_port);
   U215 : INV_X1 port map( A => opcode(1), ZN => n33);
   U216 : AND4_X1 port map( A1 => opcode(2), A2 => opcode(0), A3 => opcode(4), 
                           A4 => n169_port, ZN => n41_port);
   U217 : NOR3_X1 port map( A1 => opcode(1), A2 => opcode(5), A3 => opcode(3), 
                           ZN => n169_port);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity jump_logic_WORD_size32_NREG32_reg_file_size32 is

   port( opcode : in std_logic_vector (5 downto 0);  RSA, WB_RD, MEM_RD : in 
         std_logic_vector (4 downto 0);  Rega, ALU_out, MEM_out : in 
         std_logic_vector (31 downto 0);  Rega_new : out std_logic_vector (31 
         downto 0);  mux_s, flag : out std_logic);

end jump_logic_WORD_size32_NREG32_reg_file_size32;

architecture SYN_Behavioral of jump_logic_WORD_size32_NREG32_reg_file_size32 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, Rega_new_31_port, Rega_new_30_port, Rega_new_29_port, 
      Rega_new_28_port, Rega_new_27_port, Rega_new_26_port, Rega_new_25_port, 
      Rega_new_24_port, Rega_new_23_port, Rega_new_22_port, Rega_new_21_port, 
      Rega_new_20_port, Rega_new_19_port, Rega_new_18_port, Rega_new_17_port, 
      Rega_new_16_port, Rega_new_15_port, Rega_new_14_port, Rega_new_13_port, 
      Rega_new_12_port, Rega_new_11_port, Rega_new_10_port, Rega_new_9_port, 
      Rega_new_8_port, Rega_new_7_port, Rega_new_6_port, Rega_new_5_port, 
      Rega_new_4_port, Rega_new_3_port, Rega_new_2_port, Rega_new_1_port, 
      Rega_new_0_port : std_logic;

begin
   Rega_new <= ( Rega_new_31_port, Rega_new_30_port, Rega_new_29_port, 
      Rega_new_28_port, Rega_new_27_port, Rega_new_26_port, Rega_new_25_port, 
      Rega_new_24_port, Rega_new_23_port, Rega_new_22_port, Rega_new_21_port, 
      Rega_new_20_port, Rega_new_19_port, Rega_new_18_port, Rega_new_17_port, 
      Rega_new_16_port, Rega_new_15_port, Rega_new_14_port, Rega_new_13_port, 
      Rega_new_12_port, Rega_new_11_port, Rega_new_10_port, Rega_new_9_port, 
      Rega_new_8_port, Rega_new_7_port, Rega_new_6_port, Rega_new_5_port, 
      Rega_new_4_port, Rega_new_3_port, Rega_new_2_port, Rega_new_1_port, 
      Rega_new_0_port );
   
   U3 : BUF_X1 port map( A => n11, Z => n1);
   U4 : BUF_X1 port map( A => n11, Z => n2);
   U5 : BUF_X1 port map( A => n11, Z => n3);
   U6 : BUF_X1 port map( A => n12, Z => n5);
   U7 : BUF_X1 port map( A => n12, Z => n4);
   U8 : BUF_X1 port map( A => n13, Z => n8);
   U9 : BUF_X1 port map( A => n13, Z => n7);
   U10 : BUF_X1 port map( A => n12, Z => n6);
   U11 : BUF_X1 port map( A => n13, Z => n9);
   U12 : INV_X1 port map( A => n10, ZN => Rega_new_31_port);
   U13 : AOI222_X1 port map( A1 => ALU_out(31), A2 => n1, B1 => MEM_out(31), B2
                           => n6, C1 => Rega(31), C2 => n9, ZN => n10);
   U14 : INV_X1 port map( A => n14, ZN => Rega_new_30_port);
   U15 : INV_X1 port map( A => n15, ZN => Rega_new_29_port);
   U16 : INV_X1 port map( A => n16, ZN => Rega_new_28_port);
   U17 : INV_X1 port map( A => n17, ZN => Rega_new_27_port);
   U18 : INV_X1 port map( A => n18, ZN => Rega_new_26_port);
   U19 : INV_X1 port map( A => n19, ZN => Rega_new_25_port);
   U20 : INV_X1 port map( A => n20, ZN => Rega_new_24_port);
   U21 : INV_X1 port map( A => n21, ZN => Rega_new_23_port);
   U22 : INV_X1 port map( A => n22, ZN => Rega_new_22_port);
   U23 : INV_X1 port map( A => n23, ZN => Rega_new_21_port);
   U24 : INV_X1 port map( A => n24, ZN => Rega_new_20_port);
   U25 : INV_X1 port map( A => n25, ZN => Rega_new_19_port);
   U26 : INV_X1 port map( A => n26, ZN => Rega_new_18_port);
   U27 : INV_X1 port map( A => n27, ZN => Rega_new_17_port);
   U28 : INV_X1 port map( A => n28, ZN => Rega_new_16_port);
   U29 : INV_X1 port map( A => n29, ZN => Rega_new_15_port);
   U30 : INV_X1 port map( A => n30, ZN => Rega_new_6_port);
   U31 : INV_X1 port map( A => n31, ZN => Rega_new_5_port);
   U32 : INV_X1 port map( A => n32, ZN => Rega_new_4_port);
   U33 : INV_X1 port map( A => n33, ZN => Rega_new_3_port);
   U34 : AND4_X1 port map( A1 => n34, A2 => n35, A3 => opcode(1), A4 => 
                           opcode(4), ZN => mux_s);
   U35 : OAI22_X1 port map( A1 => n36, A2 => n37, B1 => n38, B2 => n39, ZN => 
                           flag);
   U36 : INV_X1 port map( A => n35, ZN => n39);
   U37 : AOI22_X1 port map( A1 => n40, A2 => n41, B1 => opcode(1), B2 => n34, 
                           ZN => n38);
   U38 : AND2_X1 port map( A1 => n37, A2 => n36, ZN => n40);
   U39 : NAND3_X1 port map( A1 => n42, A2 => n35, A3 => n41, ZN => n37);
   U40 : NOR3_X1 port map( A1 => opcode(1), A2 => opcode(4), A3 => n34, ZN => 
                           n41);
   U41 : INV_X1 port map( A => opcode(2), ZN => n34);
   U42 : NOR2_X1 port map( A1 => opcode(5), A2 => opcode(3), ZN => n35);
   U43 : INV_X1 port map( A => opcode(0), ZN => n42);
   U44 : NAND4_X1 port map( A1 => n43, A2 => n44, A3 => n45, A4 => n46, ZN => 
                           n36);
   U45 : NOR4_X1 port map( A1 => n47, A2 => n48, A3 => n49, A4 => n50, ZN => 
                           n46);
   U46 : NAND4_X1 port map( A1 => n29, A2 => n28, A3 => n27, A4 => n26, ZN => 
                           n50);
   U47 : AOI222_X1 port map( A1 => ALU_out(18), A2 => n1, B1 => MEM_out(18), B2
                           => n6, C1 => Rega(18), C2 => n9, ZN => n26);
   U48 : AOI222_X1 port map( A1 => ALU_out(17), A2 => n1, B1 => MEM_out(17), B2
                           => n6, C1 => Rega(17), C2 => n9, ZN => n27);
   U49 : AOI222_X1 port map( A1 => ALU_out(16), A2 => n1, B1 => MEM_out(16), B2
                           => n6, C1 => Rega(16), C2 => n9, ZN => n28);
   U50 : AOI222_X1 port map( A1 => ALU_out(15), A2 => n1, B1 => MEM_out(15), B2
                           => n6, C1 => Rega(15), C2 => n9, ZN => n29);
   U51 : NAND4_X1 port map( A1 => n25, A2 => n24, A3 => n23, A4 => n22, ZN => 
                           n49);
   U52 : AOI222_X1 port map( A1 => ALU_out(22), A2 => n1, B1 => MEM_out(22), B2
                           => n6, C1 => Rega(22), C2 => n9, ZN => n22);
   U53 : AOI222_X1 port map( A1 => ALU_out(21), A2 => n1, B1 => MEM_out(21), B2
                           => n6, C1 => Rega(21), C2 => n9, ZN => n23);
   U54 : AOI222_X1 port map( A1 => ALU_out(20), A2 => n1, B1 => MEM_out(20), B2
                           => n6, C1 => Rega(20), C2 => n9, ZN => n24);
   U55 : AOI222_X1 port map( A1 => ALU_out(19), A2 => n1, B1 => MEM_out(19), B2
                           => n6, C1 => Rega(19), C2 => n9, ZN => n25);
   U56 : NAND4_X1 port map( A1 => n21, A2 => n20, A3 => n19, A4 => n18, ZN => 
                           n48);
   U57 : AOI222_X1 port map( A1 => ALU_out(26), A2 => n1, B1 => MEM_out(26), B2
                           => n6, C1 => Rega(26), C2 => n9, ZN => n18);
   U58 : AOI222_X1 port map( A1 => ALU_out(25), A2 => n1, B1 => MEM_out(25), B2
                           => n5, C1 => Rega(25), C2 => n8, ZN => n19);
   U59 : AOI222_X1 port map( A1 => ALU_out(24), A2 => n2, B1 => MEM_out(24), B2
                           => n5, C1 => Rega(24), C2 => n8, ZN => n20);
   U60 : AOI222_X1 port map( A1 => ALU_out(23), A2 => n2, B1 => MEM_out(23), B2
                           => n5, C1 => Rega(23), C2 => n8, ZN => n21);
   U61 : NAND4_X1 port map( A1 => n17, A2 => n16, A3 => n15, A4 => n14, ZN => 
                           n47);
   U62 : AOI222_X1 port map( A1 => ALU_out(30), A2 => n2, B1 => MEM_out(30), B2
                           => n5, C1 => Rega(30), C2 => n8, ZN => n14);
   U63 : AOI222_X1 port map( A1 => ALU_out(29), A2 => n2, B1 => MEM_out(29), B2
                           => n5, C1 => Rega(29), C2 => n8, ZN => n15);
   U64 : AOI222_X1 port map( A1 => ALU_out(28), A2 => n2, B1 => MEM_out(28), B2
                           => n5, C1 => Rega(28), C2 => n8, ZN => n16);
   U65 : AOI222_X1 port map( A1 => ALU_out(27), A2 => n2, B1 => MEM_out(27), B2
                           => n5, C1 => Rega(27), C2 => n8, ZN => n17);
   U66 : NOR4_X1 port map( A1 => n51, A2 => Rega_new_0_port, A3 => 
                           Rega_new_2_port, A4 => Rega_new_1_port, ZN => n45);
   U67 : INV_X1 port map( A => n52, ZN => Rega_new_1_port);
   U68 : AOI222_X1 port map( A1 => ALU_out(1), A2 => n2, B1 => MEM_out(1), B2 
                           => n5, C1 => Rega(1), C2 => n8, ZN => n52);
   U69 : INV_X1 port map( A => n53, ZN => Rega_new_2_port);
   U70 : AOI222_X1 port map( A1 => ALU_out(2), A2 => n2, B1 => MEM_out(2), B2 
                           => n5, C1 => Rega(2), C2 => n8, ZN => n53);
   U71 : INV_X1 port map( A => n54, ZN => Rega_new_0_port);
   U72 : AOI222_X1 port map( A1 => ALU_out(0), A2 => n2, B1 => MEM_out(0), B2 
                           => n5, C1 => Rega(0), C2 => n8, ZN => n54);
   U73 : NAND4_X1 port map( A1 => n33, A2 => n32, A3 => n31, A4 => n30, ZN => 
                           n51);
   U74 : AOI222_X1 port map( A1 => ALU_out(6), A2 => n2, B1 => MEM_out(6), B2 
                           => n5, C1 => Rega(6), C2 => n8, ZN => n30);
   U75 : AOI222_X1 port map( A1 => ALU_out(5), A2 => n2, B1 => MEM_out(5), B2 
                           => n4, C1 => Rega(5), C2 => n7, ZN => n31);
   U76 : AOI222_X1 port map( A1 => ALU_out(4), A2 => n3, B1 => MEM_out(4), B2 
                           => n4, C1 => Rega(4), C2 => n7, ZN => n32);
   U77 : AOI222_X1 port map( A1 => ALU_out(3), A2 => n3, B1 => MEM_out(3), B2 
                           => n4, C1 => Rega(3), C2 => n7, ZN => n33);
   U78 : NOR4_X1 port map( A1 => Rega_new_14_port, A2 => Rega_new_13_port, A3 
                           => Rega_new_12_port, A4 => Rega_new_11_port, ZN => 
                           n44);
   U79 : INV_X1 port map( A => n55, ZN => Rega_new_11_port);
   U80 : AOI222_X1 port map( A1 => ALU_out(11), A2 => n3, B1 => MEM_out(11), B2
                           => n4, C1 => Rega(11), C2 => n7, ZN => n55);
   U81 : INV_X1 port map( A => n56, ZN => Rega_new_12_port);
   U82 : AOI222_X1 port map( A1 => ALU_out(12), A2 => n3, B1 => MEM_out(12), B2
                           => n4, C1 => Rega(12), C2 => n7, ZN => n56);
   U83 : INV_X1 port map( A => n57, ZN => Rega_new_13_port);
   U84 : AOI222_X1 port map( A1 => ALU_out(13), A2 => n3, B1 => MEM_out(13), B2
                           => n4, C1 => Rega(13), C2 => n7, ZN => n57);
   U85 : INV_X1 port map( A => n58, ZN => Rega_new_14_port);
   U86 : AOI222_X1 port map( A1 => ALU_out(14), A2 => n3, B1 => MEM_out(14), B2
                           => n4, C1 => Rega(14), C2 => n7, ZN => n58);
   U87 : NOR4_X1 port map( A1 => Rega_new_10_port, A2 => Rega_new_9_port, A3 =>
                           Rega_new_8_port, A4 => Rega_new_7_port, ZN => n43);
   U88 : INV_X1 port map( A => n59, ZN => Rega_new_7_port);
   U89 : AOI222_X1 port map( A1 => ALU_out(7), A2 => n3, B1 => MEM_out(7), B2 
                           => n4, C1 => Rega(7), C2 => n7, ZN => n59);
   U90 : INV_X1 port map( A => n60, ZN => Rega_new_8_port);
   U91 : AOI222_X1 port map( A1 => ALU_out(8), A2 => n3, B1 => MEM_out(8), B2 
                           => n4, C1 => Rega(8), C2 => n7, ZN => n60);
   U92 : INV_X1 port map( A => n61, ZN => Rega_new_9_port);
   U93 : AOI222_X1 port map( A1 => ALU_out(9), A2 => n3, B1 => MEM_out(9), B2 
                           => n4, C1 => Rega(9), C2 => n7, ZN => n61);
   U94 : INV_X1 port map( A => n62, ZN => Rega_new_10_port);
   U95 : AOI222_X1 port map( A1 => ALU_out(10), A2 => n3, B1 => MEM_out(10), B2
                           => n4, C1 => Rega(10), C2 => n7, ZN => n62);
   U96 : AND2_X1 port map( A1 => n63, A2 => n64, ZN => n13);
   U97 : NOR2_X1 port map( A1 => n63, A2 => n3, ZN => n12);
   U98 : NAND4_X1 port map( A1 => n65, A2 => n66, A3 => n67, A4 => n68, ZN => 
                           n63);
   U99 : NOR2_X1 port map( A1 => n69, A2 => n70, ZN => n68);
   U100 : XOR2_X1 port map( A => WB_RD(4), B => RSA(4), Z => n70);
   U101 : XOR2_X1 port map( A => WB_RD(2), B => RSA(2), Z => n69);
   U102 : XNOR2_X1 port map( A => RSA(0), B => WB_RD(0), ZN => n67);
   U103 : XNOR2_X1 port map( A => RSA(1), B => WB_RD(1), ZN => n66);
   U104 : XNOR2_X1 port map( A => RSA(3), B => WB_RD(3), ZN => n65);
   U105 : INV_X1 port map( A => n64, ZN => n11);
   U106 : NAND3_X1 port map( A1 => n71, A2 => n72, A3 => n73, ZN => n64);
   U107 : NOR3_X1 port map( A1 => n74, A2 => n75, A3 => n76, ZN => n73);
   U108 : XOR2_X1 port map( A => RSA(3), B => MEM_RD(3), Z => n76);
   U109 : XOR2_X1 port map( A => RSA(1), B => MEM_RD(1), Z => n75);
   U110 : XOR2_X1 port map( A => RSA(0), B => MEM_RD(0), Z => n74);
   U111 : XNOR2_X1 port map( A => RSA(2), B => MEM_RD(2), ZN => n72);
   U112 : XNOR2_X1 port map( A => RSA(4), B => MEM_RD(4), ZN => n71);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity P4_ADDER_NBIT32_0 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  S : 
         out std_logic_vector (31 downto 0);  Cout, ovf : out std_logic);

end P4_ADDER_NBIT32_0;

architecture SYN_STRUCTURAL of P4_ADDER_NBIT32_0 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component sum_generator_n_bit32_n_CSB8_0
      port( A, B : in std_logic_vector (31 downto 0);  C_in : in 
            std_logic_vector (7 downto 0);  S : out std_logic_vector (31 downto
            0));
   end component;
   
   component CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_0
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  Co 
            : out std_logic_vector (7 downto 0));
   end component;
   
   component my_xor_225
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_226
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_227
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_228
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_229
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_230
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_231
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_232
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_233
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_234
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_235
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_236
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_237
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_238
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_239
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_240
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_241
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_242
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_243
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_244
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_245
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_246
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_247
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_248
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_249
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_250
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_251
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_252
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_253
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_254
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_255
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component my_xor_0
      port( A, B : in std_logic;  xor_out : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal S_31_port, S_30_port, S_29_port, S_28_port, S_27_port, S_26_port, 
      S_25_port, S_24_port, S_23_port, S_22_port, S_21_port, S_20_port, 
      S_19_port, S_18_port, S_17_port, S_16_port, S_15_port, S_14_port, 
      S_13_port, S_12_port, S_11_port, S_10_port, S_9_port, S_8_port, S_7_port,
      S_6_port, S_5_port, S_4_port, S_3_port, S_2_port, S_1_port, S_0_port, 
      xor_b_31_port, xor_b_30_port, xor_b_29_port, xor_b_28_port, xor_b_27_port
      , xor_b_26_port, xor_b_25_port, xor_b_24_port, xor_b_23_port, 
      xor_b_22_port, xor_b_21_port, xor_b_20_port, xor_b_19_port, xor_b_18_port
      , xor_b_17_port, xor_b_16_port, xor_b_15_port, xor_b_14_port, 
      xor_b_13_port, xor_b_12_port, xor_b_11_port, xor_b_10_port, xor_b_9_port,
      xor_b_8_port, xor_b_7_port, xor_b_6_port, xor_b_5_port, xor_b_4_port, 
      xor_b_3_port, xor_b_2_port, xor_b_1_port, xor_b_0_port, carry_6_port, 
      carry_5_port, carry_4_port, carry_3_port, carry_2_port, carry_1_port, 
      carry_0_port, n1, n2 : std_logic;

begin
   S <= ( S_31_port, S_30_port, S_29_port, S_28_port, S_27_port, S_26_port, 
      S_25_port, S_24_port, S_23_port, S_22_port, S_21_port, S_20_port, 
      S_19_port, S_18_port, S_17_port, S_16_port, S_15_port, S_14_port, 
      S_13_port, S_12_port, S_11_port, S_10_port, S_9_port, S_8_port, S_7_port,
      S_6_port, S_5_port, S_4_port, S_3_port, S_2_port, S_1_port, S_0_port );
   
   U3 : XOR2_X1 port map( A => xor_b_31_port, B => A(31), Z => n2);
   bc_xor_31 : my_xor_0 port map( A => B(31), B => Cin, xor_out => 
                           xor_b_31_port);
   bc_xor_30 : my_xor_255 port map( A => B(30), B => Cin, xor_out => 
                           xor_b_30_port);
   bc_xor_29 : my_xor_254 port map( A => B(29), B => Cin, xor_out => 
                           xor_b_29_port);
   bc_xor_28 : my_xor_253 port map( A => B(28), B => Cin, xor_out => 
                           xor_b_28_port);
   bc_xor_27 : my_xor_252 port map( A => B(27), B => Cin, xor_out => 
                           xor_b_27_port);
   bc_xor_26 : my_xor_251 port map( A => B(26), B => Cin, xor_out => 
                           xor_b_26_port);
   bc_xor_25 : my_xor_250 port map( A => B(25), B => Cin, xor_out => 
                           xor_b_25_port);
   bc_xor_24 : my_xor_249 port map( A => B(24), B => Cin, xor_out => 
                           xor_b_24_port);
   bc_xor_23 : my_xor_248 port map( A => B(23), B => Cin, xor_out => 
                           xor_b_23_port);
   bc_xor_22 : my_xor_247 port map( A => B(22), B => Cin, xor_out => 
                           xor_b_22_port);
   bc_xor_21 : my_xor_246 port map( A => B(21), B => Cin, xor_out => 
                           xor_b_21_port);
   bc_xor_20 : my_xor_245 port map( A => B(20), B => Cin, xor_out => 
                           xor_b_20_port);
   bc_xor_19 : my_xor_244 port map( A => B(19), B => Cin, xor_out => 
                           xor_b_19_port);
   bc_xor_18 : my_xor_243 port map( A => B(18), B => Cin, xor_out => 
                           xor_b_18_port);
   bc_xor_17 : my_xor_242 port map( A => B(17), B => Cin, xor_out => 
                           xor_b_17_port);
   bc_xor_16 : my_xor_241 port map( A => B(16), B => Cin, xor_out => 
                           xor_b_16_port);
   bc_xor_15 : my_xor_240 port map( A => B(15), B => Cin, xor_out => 
                           xor_b_15_port);
   bc_xor_14 : my_xor_239 port map( A => B(14), B => Cin, xor_out => 
                           xor_b_14_port);
   bc_xor_13 : my_xor_238 port map( A => B(13), B => Cin, xor_out => 
                           xor_b_13_port);
   bc_xor_12 : my_xor_237 port map( A => B(12), B => Cin, xor_out => 
                           xor_b_12_port);
   bc_xor_11 : my_xor_236 port map( A => B(11), B => Cin, xor_out => 
                           xor_b_11_port);
   bc_xor_10 : my_xor_235 port map( A => B(10), B => Cin, xor_out => 
                           xor_b_10_port);
   bc_xor_9 : my_xor_234 port map( A => B(9), B => Cin, xor_out => xor_b_9_port
                           );
   bc_xor_8 : my_xor_233 port map( A => B(8), B => Cin, xor_out => xor_b_8_port
                           );
   bc_xor_7 : my_xor_232 port map( A => B(7), B => Cin, xor_out => xor_b_7_port
                           );
   bc_xor_6 : my_xor_231 port map( A => B(6), B => Cin, xor_out => xor_b_6_port
                           );
   bc_xor_5 : my_xor_230 port map( A => B(5), B => Cin, xor_out => xor_b_5_port
                           );
   bc_xor_4 : my_xor_229 port map( A => B(4), B => Cin, xor_out => xor_b_4_port
                           );
   bc_xor_3 : my_xor_228 port map( A => B(3), B => Cin, xor_out => xor_b_3_port
                           );
   bc_xor_2 : my_xor_227 port map( A => B(2), B => Cin, xor_out => xor_b_2_port
                           );
   bc_xor_1 : my_xor_226 port map( A => B(1), B => Cin, xor_out => xor_b_1_port
                           );
   bc_xor_0 : my_xor_225 port map( A => B(0), B => Cin, xor_out => xor_b_0_port
                           );
   CG : CARRY_GENERATOR_NBIT32_NBIT_PER_BLOCK4_0 port map( A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(31) => 
                           xor_b_31_port, B(30) => xor_b_30_port, B(29) => 
                           xor_b_29_port, B(28) => xor_b_28_port, B(27) => 
                           xor_b_27_port, B(26) => xor_b_26_port, B(25) => 
                           xor_b_25_port, B(24) => xor_b_24_port, B(23) => 
                           xor_b_23_port, B(22) => xor_b_22_port, B(21) => 
                           xor_b_21_port, B(20) => xor_b_20_port, B(19) => 
                           xor_b_19_port, B(18) => xor_b_18_port, B(17) => 
                           xor_b_17_port, B(16) => xor_b_16_port, B(15) => 
                           xor_b_15_port, B(14) => xor_b_14_port, B(13) => 
                           xor_b_13_port, B(12) => xor_b_12_port, B(11) => 
                           xor_b_11_port, B(10) => xor_b_10_port, B(9) => 
                           xor_b_9_port, B(8) => xor_b_8_port, B(7) => 
                           xor_b_7_port, B(6) => xor_b_6_port, B(5) => 
                           xor_b_5_port, B(4) => xor_b_4_port, B(3) => 
                           xor_b_3_port, B(2) => xor_b_2_port, B(1) => 
                           xor_b_1_port, B(0) => xor_b_0_port, Cin => Cin, 
                           Co(7) => Cout, Co(6) => carry_6_port, Co(5) => 
                           carry_5_port, Co(4) => carry_4_port, Co(3) => 
                           carry_3_port, Co(2) => carry_2_port, Co(1) => 
                           carry_1_port, Co(0) => carry_0_port);
   SG : sum_generator_n_bit32_n_CSB8_0 port map( A(31) => A(31), A(30) => A(30)
                           , A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(31) => xor_b_31_port, B(30) =>
                           xor_b_30_port, B(29) => xor_b_29_port, B(28) => 
                           xor_b_28_port, B(27) => xor_b_27_port, B(26) => 
                           xor_b_26_port, B(25) => xor_b_25_port, B(24) => 
                           xor_b_24_port, B(23) => xor_b_23_port, B(22) => 
                           xor_b_22_port, B(21) => xor_b_21_port, B(20) => 
                           xor_b_20_port, B(19) => xor_b_19_port, B(18) => 
                           xor_b_18_port, B(17) => xor_b_17_port, B(16) => 
                           xor_b_16_port, B(15) => xor_b_15_port, B(14) => 
                           xor_b_14_port, B(13) => xor_b_13_port, B(12) => 
                           xor_b_12_port, B(11) => xor_b_11_port, B(10) => 
                           xor_b_10_port, B(9) => xor_b_9_port, B(8) => 
                           xor_b_8_port, B(7) => xor_b_7_port, B(6) => 
                           xor_b_6_port, B(5) => xor_b_5_port, B(4) => 
                           xor_b_4_port, B(3) => xor_b_3_port, B(2) => 
                           xor_b_2_port, B(1) => xor_b_1_port, B(0) => 
                           xor_b_0_port, C_in(7) => carry_6_port, C_in(6) => 
                           carry_5_port, C_in(5) => carry_4_port, C_in(4) => 
                           carry_3_port, C_in(3) => carry_2_port, C_in(2) => 
                           carry_1_port, C_in(1) => carry_0_port, C_in(0) => 
                           Cin, S(31) => S_31_port, S(30) => S_30_port, S(29) 
                           => S_29_port, S(28) => S_28_port, S(27) => S_27_port
                           , S(26) => S_26_port, S(25) => S_25_port, S(24) => 
                           S_24_port, S(23) => S_23_port, S(22) => S_22_port, 
                           S(21) => S_21_port, S(20) => S_20_port, S(19) => 
                           S_19_port, S(18) => S_18_port, S(17) => S_17_port, 
                           S(16) => S_16_port, S(15) => S_15_port, S(14) => 
                           S_14_port, S(13) => S_13_port, S(12) => S_12_port, 
                           S(11) => S_11_port, S(10) => S_10_port, S(9) => 
                           S_9_port, S(8) => S_8_port, S(7) => S_7_port, S(6) 
                           => S_6_port, S(5) => S_5_port, S(4) => S_4_port, 
                           S(3) => S_3_port, S(2) => S_2_port, S(1) => S_1_port
                           , S(0) => S_0_port);
   U1 : NOR2_X1 port map( A1 => n1, A2 => n2, ZN => ovf);
   U2 : XNOR2_X1 port map( A => A(31), B => S_31_port, ZN => n1);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity dec_logic_WORD_size32_NREG32 is

   port( instr, NPC_in : in std_logic_vector (31 downto 0);  opcode : out 
         std_logic_vector (5 downto 0);  RS1, RS2, RD : out std_logic_vector (4
         downto 0);  FUNC : out std_logic_vector (10 downto 0);  IMM : out 
         std_logic_vector (15 downto 0);  IMM26 : out std_logic_vector (25 
         downto 0));

end dec_logic_WORD_size32_NREG32;

architecture SYN_Behavioral of dec_logic_WORD_size32_NREG32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   signal N246, N247, N248, N249, N250, N251, N252, N253, N254, N255, N256, 
      N257, N258, N259, N260, N261, N262, N263, N264, N265, N266, N267, N268, 
      N269, N270, N271, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, 
      n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58
      , n59, n60, n61, n62, n63, n64, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, 
      n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25
      , n26, n27, n28, n29, n30, n31, n32, n65, n66, n67, n68, n69, n70 : 
      std_logic;

begin
   opcode <= ( instr(31), instr(30), instr(29), instr(28), instr(27), instr(26)
      );
   
   IMM26_reg_25_inst : DLL_X1 port map( D => N271, GN => n4, Q => IMM26(25));
   IMM26_reg_24_inst : DLL_X1 port map( D => N270, GN => n4, Q => IMM26(24));
   IMM26_reg_23_inst : DLL_X1 port map( D => N269, GN => n4, Q => IMM26(23));
   IMM26_reg_22_inst : DLL_X1 port map( D => N268, GN => n4, Q => IMM26(22));
   IMM26_reg_21_inst : DLL_X1 port map( D => N267, GN => n4, Q => IMM26(21));
   IMM26_reg_20_inst : DLL_X1 port map( D => N266, GN => n4, Q => IMM26(20));
   IMM26_reg_19_inst : DLL_X1 port map( D => N265, GN => n4, Q => IMM26(19));
   IMM26_reg_18_inst : DLL_X1 port map( D => N264, GN => n4, Q => IMM26(18));
   IMM26_reg_17_inst : DLL_X1 port map( D => N263, GN => n4, Q => IMM26(17));
   IMM26_reg_16_inst : DLL_X1 port map( D => N262, GN => n4, Q => IMM26(16));
   IMM26_reg_15_inst : DLL_X1 port map( D => N261, GN => n5, Q => IMM26(15));
   IMM26_reg_14_inst : DLL_X1 port map( D => N260, GN => n5, Q => IMM26(14));
   IMM26_reg_13_inst : DLL_X1 port map( D => N259, GN => n5, Q => IMM26(13));
   IMM26_reg_12_inst : DLL_X1 port map( D => N258, GN => n5, Q => IMM26(12));
   IMM26_reg_11_inst : DLL_X1 port map( D => N257, GN => n5, Q => IMM26(11));
   IMM26_reg_10_inst : DLL_X1 port map( D => N256, GN => n5, Q => IMM26(10));
   IMM26_reg_9_inst : DLL_X1 port map( D => N255, GN => n5, Q => IMM26(9));
   IMM26_reg_8_inst : DLL_X1 port map( D => N254, GN => n5, Q => IMM26(8));
   IMM26_reg_7_inst : DLL_X1 port map( D => N253, GN => n5, Q => IMM26(7));
   IMM26_reg_6_inst : DLL_X1 port map( D => N252, GN => n5, Q => IMM26(6));
   IMM26_reg_5_inst : DLL_X1 port map( D => N251, GN => n6, Q => IMM26(5));
   IMM26_reg_4_inst : DLL_X1 port map( D => N250, GN => n6, Q => IMM26(4));
   IMM26_reg_3_inst : DLL_X1 port map( D => N249, GN => n6, Q => IMM26(3));
   IMM26_reg_2_inst : DLL_X1 port map( D => N248, GN => n6, Q => IMM26(2));
   IMM26_reg_1_inst : DLL_X1 port map( D => N247, GN => n6, Q => IMM26(1));
   IMM26_reg_0_inst : DLL_X1 port map( D => N246, GN => n6, Q => IMM26(0));
   U134 : NAND3_X1 port map( A1 => n39, A2 => n1, A3 => instr(15), ZN => n46);
   U3 : AND2_X1 port map( A1 => n36, A2 => n41, ZN => n33);
   U4 : NOR2_X1 port map( A1 => n68, A2 => n32, ZN => RS1(4));
   U5 : NOR2_X1 port map( A1 => n68, A2 => n28, ZN => RS1(0));
   U6 : BUF_X1 port map( A => n36, Z => n2);
   U7 : INV_X1 port map( A => n34, ZN => n68);
   U8 : OR2_X1 port map( A1 => n45, A2 => n65, ZN => n47);
   U9 : NOR2_X1 port map( A1 => n68, A2 => n29, ZN => RS1(1));
   U10 : NOR2_X1 port map( A1 => n68, A2 => n30, ZN => RS1(2));
   U11 : NOR2_X1 port map( A1 => n68, A2 => n31, ZN => RS1(3));
   U12 : INV_X1 port map( A => n37, ZN => n66);
   U13 : NAND2_X1 port map( A1 => n39, A2 => n1, ZN => n45);
   U14 : INV_X1 port map( A => n39, ZN => n67);
   U15 : OAI21_X1 port map( B1 => n1, B2 => n22, A => n46, ZN => N261);
   U16 : OAI21_X1 port map( B1 => n1, B2 => n23, A => n46, ZN => N262);
   U17 : OAI21_X1 port map( B1 => n1, B2 => n24, A => n46, ZN => N263);
   U18 : OAI21_X1 port map( B1 => n1, B2 => n25, A => n46, ZN => N264);
   U19 : OAI21_X1 port map( B1 => n1, B2 => n26, A => n46, ZN => N265);
   U20 : OAI21_X1 port map( B1 => n1, B2 => n27, A => n46, ZN => N266);
   U21 : OAI21_X1 port map( B1 => n1, B2 => n28, A => n46, ZN => N267);
   U22 : OAI21_X1 port map( B1 => n1, B2 => n29, A => n46, ZN => N268);
   U23 : OAI21_X1 port map( B1 => n1, B2 => n30, A => n46, ZN => N269);
   U24 : OAI21_X1 port map( B1 => n1, B2 => n31, A => n46, ZN => N270);
   U25 : OAI21_X1 port map( B1 => n1, B2 => n32, A => n46, ZN => N271);
   U26 : BUF_X1 port map( A => n44, Z => n5);
   U27 : BUF_X1 port map( A => n44, Z => n4);
   U28 : NOR2_X1 port map( A1 => n67, A2 => n7, ZN => N246);
   U29 : NOR2_X1 port map( A1 => n67, A2 => n8, ZN => N247);
   U30 : NOR2_X1 port map( A1 => n67, A2 => n9, ZN => N248);
   U31 : NOR2_X1 port map( A1 => n67, A2 => n10, ZN => N249);
   U32 : NOR2_X1 port map( A1 => n67, A2 => n11, ZN => N250);
   U33 : NOR2_X1 port map( A1 => n67, A2 => n12, ZN => N251);
   U34 : NOR2_X1 port map( A1 => n67, A2 => n13, ZN => N252);
   U35 : NOR2_X1 port map( A1 => n67, A2 => n14, ZN => N253);
   U36 : NOR2_X1 port map( A1 => n67, A2 => n15, ZN => N254);
   U37 : NOR2_X1 port map( A1 => n67, A2 => n16, ZN => N255);
   U38 : NOR2_X1 port map( A1 => n67, A2 => n17, ZN => N256);
   U39 : NOR2_X1 port map( A1 => n67, A2 => n18, ZN => N257);
   U40 : NOR2_X1 port map( A1 => n67, A2 => n19, ZN => N258);
   U41 : NOR2_X1 port map( A1 => n67, A2 => n20, ZN => N259);
   U42 : NOR2_X1 port map( A1 => n67, A2 => n21, ZN => N260);
   U43 : BUF_X1 port map( A => n44, Z => n6);
   U44 : NOR4_X1 port map( A1 => n69, A2 => instr(28), A3 => instr(29), A4 => 
                           instr(31), ZN => n64);
   U45 : INV_X1 port map( A => instr(11), ZN => n18);
   U46 : INV_X1 port map( A => instr(12), ZN => n19);
   U47 : INV_X1 port map( A => instr(14), ZN => n21);
   U48 : INV_X1 port map( A => instr(13), ZN => n20);
   U49 : INV_X1 port map( A => instr(16), ZN => n23);
   U50 : INV_X1 port map( A => instr(17), ZN => n24);
   U51 : INV_X1 port map( A => instr(18), ZN => n25);
   U52 : INV_X1 port map( A => instr(19), ZN => n26);
   U53 : INV_X1 port map( A => instr(20), ZN => n27);
   U54 : INV_X1 port map( A => instr(25), ZN => n32);
   U55 : INV_X1 port map( A => instr(24), ZN => n31);
   U56 : INV_X1 port map( A => instr(23), ZN => n30);
   U57 : INV_X1 port map( A => instr(22), ZN => n29);
   U58 : INV_X1 port map( A => instr(21), ZN => n28);
   U59 : INV_X1 port map( A => instr(15), ZN => n22);
   U60 : OAI21_X1 port map( B1 => n65, B2 => n46, A => n57, ZN => IMM(15));
   U61 : NAND2_X1 port map( A1 => NPC_in(15), A2 => n66, ZN => n57);
   U62 : OAI21_X1 port map( B1 => n21, B2 => n47, A => n58, ZN => IMM(14));
   U63 : NAND2_X1 port map( A1 => NPC_in(14), A2 => n66, ZN => n58);
   U64 : OAI21_X1 port map( B1 => n20, B2 => n47, A => n59, ZN => IMM(13));
   U65 : NAND2_X1 port map( A1 => NPC_in(13), A2 => n66, ZN => n59);
   U66 : OAI21_X1 port map( B1 => n19, B2 => n47, A => n60, ZN => IMM(12));
   U67 : NAND2_X1 port map( A1 => NPC_in(12), A2 => n66, ZN => n60);
   U68 : OAI21_X1 port map( B1 => n18, B2 => n47, A => n61, ZN => IMM(11));
   U69 : NAND2_X1 port map( A1 => NPC_in(11), A2 => n66, ZN => n61);
   U70 : OAI21_X1 port map( B1 => n17, B2 => n47, A => n62, ZN => IMM(10));
   U71 : NAND2_X1 port map( A1 => NPC_in(10), A2 => n66, ZN => n62);
   U72 : OAI21_X1 port map( B1 => n16, B2 => n47, A => n48, ZN => IMM(9));
   U73 : NAND2_X1 port map( A1 => NPC_in(9), A2 => n66, ZN => n48);
   U74 : OAI21_X1 port map( B1 => n15, B2 => n47, A => n49, ZN => IMM(8));
   U75 : NAND2_X1 port map( A1 => NPC_in(8), A2 => n66, ZN => n49);
   U76 : OAI21_X1 port map( B1 => n14, B2 => n47, A => n50, ZN => IMM(7));
   U77 : NAND2_X1 port map( A1 => NPC_in(7), A2 => n66, ZN => n50);
   U78 : OAI21_X1 port map( B1 => n13, B2 => n47, A => n51, ZN => IMM(6));
   U79 : NAND2_X1 port map( A1 => NPC_in(6), A2 => n66, ZN => n51);
   U80 : OAI21_X1 port map( B1 => n12, B2 => n47, A => n52, ZN => IMM(5));
   U81 : NAND2_X1 port map( A1 => NPC_in(5), A2 => n66, ZN => n52);
   U82 : OAI21_X1 port map( B1 => n11, B2 => n47, A => n53, ZN => IMM(4));
   U83 : NAND2_X1 port map( A1 => NPC_in(4), A2 => n66, ZN => n53);
   U84 : OAI21_X1 port map( B1 => n10, B2 => n47, A => n54, ZN => IMM(3));
   U85 : NAND2_X1 port map( A1 => NPC_in(3), A2 => n66, ZN => n54);
   U86 : OAI21_X1 port map( B1 => n9, B2 => n47, A => n55, ZN => IMM(2));
   U87 : NAND2_X1 port map( A1 => NPC_in(2), A2 => n66, ZN => n55);
   U88 : OAI21_X1 port map( B1 => n8, B2 => n47, A => n56, ZN => IMM(1));
   U89 : NAND2_X1 port map( A1 => NPC_in(1), A2 => n66, ZN => n56);
   U90 : OAI21_X1 port map( B1 => n7, B2 => n47, A => n63, ZN => IMM(0));
   U91 : NAND2_X1 port map( A1 => NPC_in(0), A2 => n66, ZN => n63);
   U92 : INV_X1 port map( A => instr(8), ZN => n15);
   U93 : INV_X1 port map( A => instr(9), ZN => n16);
   U94 : INV_X1 port map( A => instr(10), ZN => n17);
   U95 : INV_X1 port map( A => instr(7), ZN => n14);
   U96 : INV_X1 port map( A => instr(3), ZN => n10);
   U97 : INV_X1 port map( A => instr(4), ZN => n11);
   U98 : INV_X1 port map( A => instr(6), ZN => n13);
   U99 : INV_X1 port map( A => instr(5), ZN => n12);
   U100 : INV_X1 port map( A => instr(1), ZN => n8);
   U101 : INV_X1 port map( A => instr(2), ZN => n9);
   U102 : INV_X1 port map( A => instr(0), ZN => n7);
   U103 : NAND2_X1 port map( A1 => instr(26), A2 => n64, ZN => n37);
   U104 : NOR2_X1 port map( A1 => n33, A2 => n27, ZN => RS2(4));
   U105 : NOR2_X1 port map( A1 => n33, A2 => n25, ZN => RS2(2));
   U106 : NOR2_X1 port map( A1 => n33, A2 => n23, ZN => RS2(0));
   U107 : NOR2_X1 port map( A1 => n33, A2 => n24, ZN => RS2(1));
   U108 : NOR2_X1 port map( A1 => n33, A2 => n26, ZN => RS2(3));
   U109 : NAND4_X1 port map( A1 => instr(31), A2 => instr(29), A3 => n42, A4 =>
                           n70, ZN => n41);
   U110 : CLKBUF_X1 port map( A => n34, Z => n1);
   U111 : NAND2_X1 port map( A1 => n64, A2 => n70, ZN => n34);
   U112 : NAND2_X1 port map( A1 => n3, A2 => n43, ZN => n36);
   U113 : BUF_X1 port map( A => n40, Z => n3);
   U114 : NOR4_X1 port map( A1 => instr(27), A2 => instr(29), A3 => instr(30), 
                           A4 => instr(31), ZN => n40);
   U115 : NOR2_X1 port map( A1 => instr(28), A2 => instr(26), ZN => n43);
   U116 : OAI221_X1 port map( B1 => n26, B2 => n35, C1 => n2, C2 => n21, A => 
                           n37, ZN => RD(3));
   U117 : OAI221_X1 port map( B1 => n27, B2 => n35, C1 => n2, C2 => n22, A => 
                           n37, ZN => RD(4));
   U118 : OAI221_X1 port map( B1 => n25, B2 => n35, C1 => n2, C2 => n20, A => 
                           n37, ZN => RD(2));
   U119 : INV_X1 port map( A => instr(27), ZN => n69);
   U120 : OAI22_X1 port map( A1 => instr(28), A2 => instr(27), B1 => n43, B2 =>
                           n69, ZN => n42);
   U121 : OAI221_X1 port map( B1 => n23, B2 => n35, C1 => n2, C2 => n18, A => 
                           n37, ZN => RD(0));
   U122 : OAI221_X1 port map( B1 => n24, B2 => n35, C1 => n2, C2 => n19, A => 
                           n37, ZN => RD(1));
   U123 : NAND4_X1 port map( A1 => n33, A2 => n38, A3 => n39, A4 => n34, ZN => 
                           n35);
   U124 : AOI21_X1 port map( B1 => n3, B2 => instr(28), A => n45, ZN => n44);
   U125 : INV_X1 port map( A => n2, ZN => n65);
   U126 : NOR2_X1 port map( A1 => n2, A2 => n11, ZN => FUNC(4));
   U127 : NOR2_X1 port map( A1 => n2, A2 => n13, ZN => FUNC(6));
   U128 : NOR2_X1 port map( A1 => n2, A2 => n12, ZN => FUNC(5));
   U129 : NOR2_X1 port map( A1 => n2, A2 => n8, ZN => FUNC(1));
   U130 : NOR2_X1 port map( A1 => n2, A2 => n7, ZN => FUNC(0));
   U131 : NOR2_X1 port map( A1 => n2, A2 => n10, ZN => FUNC(3));
   U132 : NOR2_X1 port map( A1 => n2, A2 => n9, ZN => FUNC(2));
   U133 : NOR2_X1 port map( A1 => n2, A2 => n14, ZN => FUNC(7));
   U135 : NOR2_X1 port map( A1 => n2, A2 => n17, ZN => FUNC(10));
   U136 : NOR2_X1 port map( A1 => n2, A2 => n16, ZN => FUNC(9));
   U137 : NOR2_X1 port map( A1 => n2, A2 => n15, ZN => FUNC(8));
   U138 : NAND2_X1 port map( A1 => instr(28), A2 => n3, ZN => n38);
   U139 : NAND2_X1 port map( A1 => instr(30), A2 => n64, ZN => n39);
   U140 : INV_X1 port map( A => instr(30), ZN => n70);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_0 is

   port( A, B, S : in std_logic;  Y : out std_logic);

end MUX21_0;

architecture SYN_BEHAVIORAL_1 of MUX21_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n1 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => Y);
   U2 : AOI22_X1 port map( A1 => A, A2 => n1, B1 => S, B2 => B, ZN => n3);
   U3 : INV_X1 port map( A => S, ZN => n1);

end SYN_BEHAVIORAL_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity WB is

   port( mem_out, alu_out : in std_logic_vector (31 downto 0);  S3 : in 
         std_logic;  output : out std_logic_vector (31 downto 0));

end WB;

architecture SYN_Behavioral of WB is

   component MUX21_GENERIC_NBIT32_2
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;

begin
   
   MUX : MUX21_GENERIC_NBIT32_2 port map( A(31) => mem_out(31), A(30) => 
                           mem_out(30), A(29) => mem_out(29), A(28) => 
                           mem_out(28), A(27) => mem_out(27), A(26) => 
                           mem_out(26), A(25) => mem_out(25), A(24) => 
                           mem_out(24), A(23) => mem_out(23), A(22) => 
                           mem_out(22), A(21) => mem_out(21), A(20) => 
                           mem_out(20), A(19) => mem_out(19), A(18) => 
                           mem_out(18), A(17) => mem_out(17), A(16) => 
                           mem_out(16), A(15) => mem_out(15), A(14) => 
                           mem_out(14), A(13) => mem_out(13), A(12) => 
                           mem_out(12), A(11) => mem_out(11), A(10) => 
                           mem_out(10), A(9) => mem_out(9), A(8) => mem_out(8),
                           A(7) => mem_out(7), A(6) => mem_out(6), A(5) => 
                           mem_out(5), A(4) => mem_out(4), A(3) => mem_out(3), 
                           A(2) => mem_out(2), A(1) => mem_out(1), A(0) => 
                           mem_out(0), B(31) => alu_out(31), B(30) => 
                           alu_out(30), B(29) => alu_out(29), B(28) => 
                           alu_out(28), B(27) => alu_out(27), B(26) => 
                           alu_out(26), B(25) => alu_out(25), B(24) => 
                           alu_out(24), B(23) => alu_out(23), B(22) => 
                           alu_out(22), B(21) => alu_out(21), B(20) => 
                           alu_out(20), B(19) => alu_out(19), B(18) => 
                           alu_out(18), B(17) => alu_out(17), B(16) => 
                           alu_out(16), B(15) => alu_out(15), B(14) => 
                           alu_out(14), B(13) => alu_out(13), B(12) => 
                           alu_out(12), B(11) => alu_out(11), B(10) => 
                           alu_out(10), B(9) => alu_out(9), B(8) => alu_out(8),
                           B(7) => alu_out(7), B(6) => alu_out(6), B(5) => 
                           alu_out(5), B(4) => alu_out(4), B(3) => alu_out(3), 
                           B(2) => alu_out(2), B(1) => alu_out(1), B(0) => 
                           alu_out(0), SEL => S3, Y(31) => output(31), Y(30) =>
                           output(30), Y(29) => output(29), Y(28) => output(28)
                           , Y(27) => output(27), Y(26) => output(26), Y(25) =>
                           output(25), Y(24) => output(24), Y(23) => output(23)
                           , Y(22) => output(22), Y(21) => output(21), Y(20) =>
                           output(20), Y(19) => output(19), Y(18) => output(18)
                           , Y(17) => output(17), Y(16) => output(16), Y(15) =>
                           output(15), Y(14) => output(14), Y(13) => output(13)
                           , Y(12) => output(12), Y(11) => output(11), Y(10) =>
                           output(10), Y(9) => output(9), Y(8) => output(8), 
                           Y(7) => output(7), Y(6) => output(6), Y(5) => 
                           output(5), Y(4) => output(4), Y(3) => output(3), 
                           Y(2) => output(2), Y(1) => output(1), Y(0) => 
                           output(0));

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MEM_MEMORY_SIZE128 is

   port( CLK, RST : in std_logic;  ALUout, MEout : in std_logic_vector (31 
         downto 0);  RDin : in std_logic_vector (4 downto 0);  DRAM_data_out : 
         in std_logic_vector (31 downto 0);  LnS, Wrd, BHU1, BHU0, EN3 : in 
         std_logic;  DRAM_addr : out std_logic_vector (8 downto 0);  
         DRAM_data_in : out std_logic_vector (31 downto 0);  MMU_out : out 
         std_logic_vector (1 downto 0);  output, alu_out : out std_logic_vector
         (31 downto 0);  RDout : out std_logic_vector (4 downto 0));

end MEM_MEMORY_SIZE128;

architecture SYN_Structural of MEM_MEMORY_SIZE128 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX51_GENERIC_NBIT32
      port( A, B, C, D, E : in std_logic_vector (31 downto 0);  SEL : in 
            std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component MMU_WORD_size32
      port( Wrd, BHU0 : in std_logic;  wdata_size : out std_logic_vector (1 
            downto 0));
   end component;
   
   signal X_Logic0_port, n1, n2, n3, n4, n5, n6 : std_logic;

begin
   DRAM_addr <= ( ALUout(8), ALUout(7), ALUout(6), ALUout(5), ALUout(4), 
      ALUout(3), ALUout(2), ALUout(1), ALUout(0) );
   DRAM_data_in <= ( MEout(31), MEout(30), MEout(29), MEout(28), MEout(27), 
      MEout(26), MEout(25), MEout(24), MEout(23), MEout(22), MEout(21), 
      MEout(20), MEout(19), MEout(18), MEout(17), MEout(16), MEout(15), 
      MEout(14), MEout(13), MEout(12), MEout(11), MEout(10), MEout(9), MEout(8)
      , MEout(7), MEout(6), MEout(5), MEout(4), MEout(3), MEout(2), MEout(1), 
      MEout(0) );
   alu_out <= ( ALUout(31), ALUout(30), ALUout(29), ALUout(28), ALUout(27), 
      ALUout(26), ALUout(25), ALUout(24), ALUout(23), ALUout(22), ALUout(21), 
      ALUout(20), ALUout(19), ALUout(18), ALUout(17), ALUout(16), ALUout(15), 
      ALUout(14), ALUout(13), ALUout(12), ALUout(11), ALUout(10), ALUout(9), 
      ALUout(8), ALUout(7), ALUout(6), ALUout(5), ALUout(4), ALUout(3), 
      ALUout(2), ALUout(1), ALUout(0) );
   RDout <= ( RDin(4), RDin(3), RDin(2), RDin(1), RDin(0) );
   
   X_Logic0_port <= '0';
   mem_MU : MMU_WORD_size32 port map( Wrd => Wrd, BHU0 => BHU0, wdata_size(1) 
                           => MMU_out(1), wdata_size(0) => MMU_out(0));
   mux : MUX51_GENERIC_NBIT32 port map( A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => n4, A(6) => DRAM_data_out(30)
                           , A(5) => DRAM_data_out(29), A(4) => 
                           DRAM_data_out(28), A(3) => DRAM_data_out(27), A(2) 
                           => DRAM_data_out(26), A(1) => DRAM_data_out(25), 
                           A(0) => DRAM_data_out(24), B(31) => X_Logic0_port, 
                           B(30) => X_Logic0_port, B(29) => X_Logic0_port, 
                           B(28) => X_Logic0_port, B(27) => X_Logic0_port, 
                           B(26) => X_Logic0_port, B(25) => X_Logic0_port, 
                           B(24) => X_Logic0_port, B(23) => X_Logic0_port, 
                           B(22) => X_Logic0_port, B(21) => X_Logic0_port, 
                           B(20) => X_Logic0_port, B(19) => X_Logic0_port, 
                           B(18) => X_Logic0_port, B(17) => X_Logic0_port, 
                           B(16) => X_Logic0_port, B(15) => n3, B(14) => 
                           DRAM_data_out(30), B(13) => DRAM_data_out(29), B(12)
                           => DRAM_data_out(28), B(11) => DRAM_data_out(27), 
                           B(10) => DRAM_data_out(26), B(9) => 
                           DRAM_data_out(25), B(8) => DRAM_data_out(24), B(7) 
                           => DRAM_data_out(23), B(6) => DRAM_data_out(22), 
                           B(5) => DRAM_data_out(21), B(4) => DRAM_data_out(20)
                           , B(3) => DRAM_data_out(19), B(2) => 
                           DRAM_data_out(18), B(1) => DRAM_data_out(17), B(0) 
                           => DRAM_data_out(16), C(31) => n3, C(30) => n3, 
                           C(29) => n3, C(28) => n3, C(27) => n3, C(26) => n3, 
                           C(25) => n3, C(24) => n3, C(23) => n3, C(22) => n3, 
                           C(21) => n4, C(20) => n4, C(19) => n4, C(18) => n4, 
                           C(17) => n4, C(16) => n4, C(15) => n4, C(14) => n4, 
                           C(13) => n4, C(12) => n4, C(11) => n4, C(10) => n5, 
                           C(9) => n5, C(8) => n5, C(7) => n5, C(6) => 
                           DRAM_data_out(30), C(5) => DRAM_data_out(29), C(4) 
                           => DRAM_data_out(28), C(3) => DRAM_data_out(27), 
                           C(2) => DRAM_data_out(26), C(1) => DRAM_data_out(25)
                           , C(0) => DRAM_data_out(24), D(31) => n5, D(30) => 
                           n5, D(29) => n5, D(28) => n5, D(27) => n5, D(26) => 
                           n5, D(25) => n5, D(24) => n5, D(23) => n5, D(22) => 
                           n6, D(21) => n6, D(20) => n6, D(19) => n6, D(18) => 
                           n6, D(17) => n6, D(16) => n6, D(15) => n6, D(14) => 
                           DRAM_data_out(30), D(13) => DRAM_data_out(29), D(12)
                           => DRAM_data_out(28), D(11) => DRAM_data_out(27), 
                           D(10) => DRAM_data_out(26), D(9) => 
                           DRAM_data_out(25), D(8) => DRAM_data_out(24), D(7) 
                           => DRAM_data_out(23), D(6) => DRAM_data_out(22), 
                           D(5) => DRAM_data_out(21), D(4) => DRAM_data_out(20)
                           , D(3) => DRAM_data_out(19), D(2) => 
                           DRAM_data_out(18), D(1) => DRAM_data_out(17), D(0) 
                           => DRAM_data_out(16), E(31) => n3, E(30) => 
                           DRAM_data_out(30), E(29) => DRAM_data_out(29), E(28)
                           => DRAM_data_out(28), E(27) => DRAM_data_out(27), 
                           E(26) => DRAM_data_out(26), E(25) => 
                           DRAM_data_out(25), E(24) => DRAM_data_out(24), E(23)
                           => DRAM_data_out(23), E(22) => DRAM_data_out(22), 
                           E(21) => DRAM_data_out(21), E(20) => 
                           DRAM_data_out(20), E(19) => DRAM_data_out(19), E(18)
                           => DRAM_data_out(18), E(17) => DRAM_data_out(17), 
                           E(16) => DRAM_data_out(16), E(15) => 
                           DRAM_data_out(15), E(14) => DRAM_data_out(14), E(13)
                           => DRAM_data_out(13), E(12) => DRAM_data_out(12), 
                           E(11) => DRAM_data_out(11), E(10) => 
                           DRAM_data_out(10), E(9) => DRAM_data_out(9), E(8) =>
                           DRAM_data_out(8), E(7) => DRAM_data_out(7), E(6) => 
                           DRAM_data_out(6), E(5) => DRAM_data_out(5), E(4) => 
                           DRAM_data_out(4), E(3) => DRAM_data_out(3), E(2) => 
                           DRAM_data_out(2), E(1) => DRAM_data_out(1), E(0) => 
                           DRAM_data_out(0), SEL(2) => Wrd, SEL(1) => BHU1, 
                           SEL(0) => BHU0, Y(31) => output(31), Y(30) => 
                           output(30), Y(29) => output(29), Y(28) => output(28)
                           , Y(27) => output(27), Y(26) => output(26), Y(25) =>
                           output(25), Y(24) => output(24), Y(23) => output(23)
                           , Y(22) => output(22), Y(21) => output(21), Y(20) =>
                           output(20), Y(19) => output(19), Y(18) => output(18)
                           , Y(17) => output(17), Y(16) => output(16), Y(15) =>
                           output(15), Y(14) => output(14), Y(13) => output(13)
                           , Y(12) => output(12), Y(11) => output(11), Y(10) =>
                           output(10), Y(9) => output(9), Y(8) => output(8), 
                           Y(7) => output(7), Y(6) => output(6), Y(5) => 
                           output(5), Y(4) => output(4), Y(3) => output(3), 
                           Y(2) => output(2), Y(1) => output(1), Y(0) => 
                           output(0));
   U2 : BUF_X1 port map( A => n2, Z => n5);
   U3 : BUF_X1 port map( A => n1, Z => n3);
   U4 : BUF_X1 port map( A => n1, Z => n4);
   U5 : BUF_X1 port map( A => n2, Z => n6);
   U6 : BUF_X1 port map( A => DRAM_data_out(31), Z => n1);
   U7 : BUF_X1 port map( A => DRAM_data_out(31), Z => n2);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity EXE is

   port( CLK, RST : in std_logic;  IMM, RA, RB : in std_logic_vector (31 downto
         0);  WA, RSA, RSB : in std_logic_vector (4 downto 0);  ALU_outmem, 
         WB_out : in std_logic_vector (31 downto 0);  MEM_RD, WB_RD : in 
         std_logic_vector (4 downto 0);  LD_EN, WB_EN, S1, S2, ALU3, ALU2, ALU1
         , ALU0, SN : in std_logic;  RD_inmul : out std_logic_vector (4 downto 
         0);  flag_structHzd, flag_ismul, OVF : out std_logic;  output, ME : 
         out std_logic_vector (31 downto 0);  WAout : out std_logic_vector (4 
         downto 0));

end EXE;

architecture SYN_Structural of EXE is

   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX21_GENERIC_NBIT5_1
      port( A, B : in std_logic_vector (4 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (4 downto 0));
   end component;
   
   component EXU_N32
      port( DATA1, DATA2 : in std_logic_vector (31 downto 0);  FUNC : in 
            std_logic_vector (3 downto 0);  RD_in : in std_logic_vector (4 
            downto 0);  SN, CLK, RST : in std_logic;  OVF, stall_flag, 
            RD_sel_flag : out std_logic;  OUTPUT : out std_logic_vector (31 
            downto 0);  RD_stall, RD_out : out std_logic_vector (4 downto 0);  
            H_MULOUT : out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT5_0
      port( A, B : in std_logic_vector (4 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (4 downto 0));
   end component;
   
   component MUX41_GENERIC_NBIT32_1
      port( A, B, C, D : in std_logic_vector (31 downto 0);  SEL : in 
            std_logic_vector (1 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component MUX41_GENERIC_NBIT32_2
      port( A, B, C, D : in std_logic_vector (31 downto 0);  SEL : in 
            std_logic_vector (1 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component MUX41_GENERIC_NBIT32_0
      port( A, B, C, D : in std_logic_vector (31 downto 0);  SEL : in 
            std_logic_vector (1 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component forwarding_unit_WORD_size32_NREG32
      port( RSA, RSB : in std_logic_vector (4 downto 0);  ALU_outmem, WB_out : 
            in std_logic_vector (31 downto 0);  MEM_RD, WB_RD : in 
            std_logic_vector (4 downto 0);  LD_EN, WB_EN, S1, S2 : in std_logic
            ;  SEL1, SEL2, SEL3 : out std_logic_vector (1 downto 0));
   end component;
   
   signal X_Logic0_port, N4, s_S1_1_port, s_S1_0_port, s_S2_1_port, s_S2_0_port
      , s_S3_1_port, s_S3_0_port, MUX1out_31_port, MUX1out_30_port, 
      MUX1out_29_port, MUX1out_28_port, MUX1out_27_port, MUX1out_26_port, 
      MUX1out_25_port, MUX1out_24_port, MUX1out_23_port, MUX1out_22_port, 
      MUX1out_21_port, MUX1out_20_port, MUX1out_19_port, MUX1out_18_port, 
      MUX1out_17_port, MUX1out_16_port, MUX1out_15_port, MUX1out_14_port, 
      MUX1out_13_port, MUX1out_12_port, MUX1out_11_port, MUX1out_10_port, 
      MUX1out_9_port, MUX1out_8_port, MUX1out_7_port, MUX1out_6_port, 
      MUX1out_5_port, MUX1out_4_port, MUX1out_3_port, MUX1out_2_port, 
      MUX1out_1_port, MUX1out_0_port, MUX2out_31_port, MUX2out_30_port, 
      MUX2out_29_port, MUX2out_28_port, MUX2out_27_port, MUX2out_26_port, 
      MUX2out_25_port, MUX2out_24_port, MUX2out_23_port, MUX2out_22_port, 
      MUX2out_21_port, MUX2out_20_port, MUX2out_19_port, MUX2out_18_port, 
      MUX2out_17_port, MUX2out_16_port, MUX2out_15_port, MUX2out_14_port, 
      MUX2out_13_port, MUX2out_12_port, MUX2out_11_port, MUX2out_10_port, 
      MUX2out_9_port, MUX2out_8_port, MUX2out_7_port, MUX2out_6_port, 
      MUX2out_5_port, MUX2out_4_port, MUX2out_3_port, MUX2out_2_port, 
      MUX2out_1_port, MUX2out_0_port, s_ALU_RD_4_port, s_ALU_RD_3_port, 
      s_ALU_RD_2_port, s_ALU_RD_1_port, s_ALU_RD_0_port, s_ovf, s_RD_sel2, 
      s_mul_RD_out_4_port, s_mul_RD_out_3_port, s_mul_RD_out_2_port, 
      s_mul_RD_out_1_port, s_mul_RD_out_0_port, n_1943, n_1944, n_1945, n_1946,
      n_1947, n_1948, n_1949, n_1950, n_1951, n_1952, n_1953, n_1954, n_1955, 
      n_1956, n_1957, n_1958, n_1959, n_1960, n_1961, n_1962, n_1963, n_1964, 
      n_1965, n_1966, n_1967, n_1968, n_1969, n_1970, n_1971, n_1972, n_1973, 
      n_1974 : std_logic;

begin
   flag_ismul <= N4;
   
   X_Logic0_port <= '0';
   FWU : forwarding_unit_WORD_size32_NREG32 port map( RSA(4) => RSA(4), RSA(3) 
                           => RSA(3), RSA(2) => RSA(2), RSA(1) => RSA(1), 
                           RSA(0) => RSA(0), RSB(4) => RSB(4), RSB(3) => RSB(3)
                           , RSB(2) => RSB(2), RSB(1) => RSB(1), RSB(0) => 
                           RSB(0), ALU_outmem(31) => ALU_outmem(31), 
                           ALU_outmem(30) => ALU_outmem(30), ALU_outmem(29) => 
                           ALU_outmem(29), ALU_outmem(28) => ALU_outmem(28), 
                           ALU_outmem(27) => ALU_outmem(27), ALU_outmem(26) => 
                           ALU_outmem(26), ALU_outmem(25) => ALU_outmem(25), 
                           ALU_outmem(24) => ALU_outmem(24), ALU_outmem(23) => 
                           ALU_outmem(23), ALU_outmem(22) => ALU_outmem(22), 
                           ALU_outmem(21) => ALU_outmem(21), ALU_outmem(20) => 
                           ALU_outmem(20), ALU_outmem(19) => ALU_outmem(19), 
                           ALU_outmem(18) => ALU_outmem(18), ALU_outmem(17) => 
                           ALU_outmem(17), ALU_outmem(16) => ALU_outmem(16), 
                           ALU_outmem(15) => ALU_outmem(15), ALU_outmem(14) => 
                           ALU_outmem(14), ALU_outmem(13) => ALU_outmem(13), 
                           ALU_outmem(12) => ALU_outmem(12), ALU_outmem(11) => 
                           ALU_outmem(11), ALU_outmem(10) => ALU_outmem(10), 
                           ALU_outmem(9) => ALU_outmem(9), ALU_outmem(8) => 
                           ALU_outmem(8), ALU_outmem(7) => ALU_outmem(7), 
                           ALU_outmem(6) => ALU_outmem(6), ALU_outmem(5) => 
                           ALU_outmem(5), ALU_outmem(4) => ALU_outmem(4), 
                           ALU_outmem(3) => ALU_outmem(3), ALU_outmem(2) => 
                           ALU_outmem(2), ALU_outmem(1) => ALU_outmem(1), 
                           ALU_outmem(0) => ALU_outmem(0), WB_out(31) => 
                           WB_out(31), WB_out(30) => WB_out(30), WB_out(29) => 
                           WB_out(29), WB_out(28) => WB_out(28), WB_out(27) => 
                           WB_out(27), WB_out(26) => WB_out(26), WB_out(25) => 
                           WB_out(25), WB_out(24) => WB_out(24), WB_out(23) => 
                           WB_out(23), WB_out(22) => WB_out(22), WB_out(21) => 
                           WB_out(21), WB_out(20) => WB_out(20), WB_out(19) => 
                           WB_out(19), WB_out(18) => WB_out(18), WB_out(17) => 
                           WB_out(17), WB_out(16) => WB_out(16), WB_out(15) => 
                           WB_out(15), WB_out(14) => WB_out(14), WB_out(13) => 
                           WB_out(13), WB_out(12) => WB_out(12), WB_out(11) => 
                           WB_out(11), WB_out(10) => WB_out(10), WB_out(9) => 
                           WB_out(9), WB_out(8) => WB_out(8), WB_out(7) => 
                           WB_out(7), WB_out(6) => WB_out(6), WB_out(5) => 
                           WB_out(5), WB_out(4) => WB_out(4), WB_out(3) => 
                           WB_out(3), WB_out(2) => WB_out(2), WB_out(1) => 
                           WB_out(1), WB_out(0) => WB_out(0), MEM_RD(4) => 
                           MEM_RD(4), MEM_RD(3) => MEM_RD(3), MEM_RD(2) => 
                           MEM_RD(2), MEM_RD(1) => MEM_RD(1), MEM_RD(0) => 
                           MEM_RD(0), WB_RD(4) => WB_RD(4), WB_RD(3) => 
                           WB_RD(3), WB_RD(2) => WB_RD(2), WB_RD(1) => WB_RD(1)
                           , WB_RD(0) => WB_RD(0), LD_EN => LD_EN, WB_EN => 
                           WB_EN, S1 => S1, S2 => S2, SEL1(1) => s_S1_1_port, 
                           SEL1(0) => s_S1_0_port, SEL2(1) => s_S2_1_port, 
                           SEL2(0) => s_S2_0_port, SEL3(1) => s_S3_1_port, 
                           SEL3(0) => s_S3_0_port);
   FW_MUX1 : MUX41_GENERIC_NBIT32_0 port map( A(31) => IMM(31), A(30) => 
                           IMM(30), A(29) => IMM(29), A(28) => IMM(28), A(27) 
                           => IMM(27), A(26) => IMM(26), A(25) => IMM(25), 
                           A(24) => IMM(24), A(23) => IMM(23), A(22) => IMM(22)
                           , A(21) => IMM(21), A(20) => IMM(20), A(19) => 
                           IMM(19), A(18) => IMM(18), A(17) => IMM(17), A(16) 
                           => IMM(16), A(15) => IMM(15), A(14) => IMM(14), 
                           A(13) => IMM(13), A(12) => IMM(12), A(11) => IMM(11)
                           , A(10) => IMM(10), A(9) => IMM(9), A(8) => IMM(8), 
                           A(7) => IMM(7), A(6) => IMM(6), A(5) => IMM(5), A(4)
                           => IMM(4), A(3) => IMM(3), A(2) => IMM(2), A(1) => 
                           IMM(1), A(0) => IMM(0), B(31) => RA(31), B(30) => 
                           RA(30), B(29) => RA(29), B(28) => RA(28), B(27) => 
                           RA(27), B(26) => RA(26), B(25) => RA(25), B(24) => 
                           RA(24), B(23) => RA(23), B(22) => RA(22), B(21) => 
                           RA(21), B(20) => RA(20), B(19) => RA(19), B(18) => 
                           RA(18), B(17) => RA(17), B(16) => RA(16), B(15) => 
                           RA(15), B(14) => RA(14), B(13) => RA(13), B(12) => 
                           RA(12), B(11) => RA(11), B(10) => RA(10), B(9) => 
                           RA(9), B(8) => RA(8), B(7) => RA(7), B(6) => RA(6), 
                           B(5) => RA(5), B(4) => RA(4), B(3) => RA(3), B(2) =>
                           RA(2), B(1) => RA(1), B(0) => RA(0), C(31) => 
                           ALU_outmem(31), C(30) => ALU_outmem(30), C(29) => 
                           ALU_outmem(29), C(28) => ALU_outmem(28), C(27) => 
                           ALU_outmem(27), C(26) => ALU_outmem(26), C(25) => 
                           ALU_outmem(25), C(24) => ALU_outmem(24), C(23) => 
                           ALU_outmem(23), C(22) => ALU_outmem(22), C(21) => 
                           ALU_outmem(21), C(20) => ALU_outmem(20), C(19) => 
                           ALU_outmem(19), C(18) => ALU_outmem(18), C(17) => 
                           ALU_outmem(17), C(16) => ALU_outmem(16), C(15) => 
                           ALU_outmem(15), C(14) => ALU_outmem(14), C(13) => 
                           ALU_outmem(13), C(12) => ALU_outmem(12), C(11) => 
                           ALU_outmem(11), C(10) => ALU_outmem(10), C(9) => 
                           ALU_outmem(9), C(8) => ALU_outmem(8), C(7) => 
                           ALU_outmem(7), C(6) => ALU_outmem(6), C(5) => 
                           ALU_outmem(5), C(4) => ALU_outmem(4), C(3) => 
                           ALU_outmem(3), C(2) => ALU_outmem(2), C(1) => 
                           ALU_outmem(1), C(0) => ALU_outmem(0), D(31) => 
                           WB_out(31), D(30) => WB_out(30), D(29) => WB_out(29)
                           , D(28) => WB_out(28), D(27) => WB_out(27), D(26) =>
                           WB_out(26), D(25) => WB_out(25), D(24) => WB_out(24)
                           , D(23) => WB_out(23), D(22) => WB_out(22), D(21) =>
                           WB_out(21), D(20) => WB_out(20), D(19) => WB_out(19)
                           , D(18) => WB_out(18), D(17) => WB_out(17), D(16) =>
                           WB_out(16), D(15) => WB_out(15), D(14) => WB_out(14)
                           , D(13) => WB_out(13), D(12) => WB_out(12), D(11) =>
                           WB_out(11), D(10) => WB_out(10), D(9) => WB_out(9), 
                           D(8) => WB_out(8), D(7) => WB_out(7), D(6) => 
                           WB_out(6), D(5) => WB_out(5), D(4) => WB_out(4), 
                           D(3) => WB_out(3), D(2) => WB_out(2), D(1) => 
                           WB_out(1), D(0) => WB_out(0), SEL(1) => s_S1_1_port,
                           SEL(0) => s_S1_0_port, Y(31) => MUX1out_31_port, 
                           Y(30) => MUX1out_30_port, Y(29) => MUX1out_29_port, 
                           Y(28) => MUX1out_28_port, Y(27) => MUX1out_27_port, 
                           Y(26) => MUX1out_26_port, Y(25) => MUX1out_25_port, 
                           Y(24) => MUX1out_24_port, Y(23) => MUX1out_23_port, 
                           Y(22) => MUX1out_22_port, Y(21) => MUX1out_21_port, 
                           Y(20) => MUX1out_20_port, Y(19) => MUX1out_19_port, 
                           Y(18) => MUX1out_18_port, Y(17) => MUX1out_17_port, 
                           Y(16) => MUX1out_16_port, Y(15) => MUX1out_15_port, 
                           Y(14) => MUX1out_14_port, Y(13) => MUX1out_13_port, 
                           Y(12) => MUX1out_12_port, Y(11) => MUX1out_11_port, 
                           Y(10) => MUX1out_10_port, Y(9) => MUX1out_9_port, 
                           Y(8) => MUX1out_8_port, Y(7) => MUX1out_7_port, Y(6)
                           => MUX1out_6_port, Y(5) => MUX1out_5_port, Y(4) => 
                           MUX1out_4_port, Y(3) => MUX1out_3_port, Y(2) => 
                           MUX1out_2_port, Y(1) => MUX1out_1_port, Y(0) => 
                           MUX1out_0_port);
   FW_MUX2 : MUX41_GENERIC_NBIT32_2 port map( A(31) => RB(31), A(30) => RB(30),
                           A(29) => RB(29), A(28) => RB(28), A(27) => RB(27), 
                           A(26) => RB(26), A(25) => RB(25), A(24) => RB(24), 
                           A(23) => RB(23), A(22) => RB(22), A(21) => RB(21), 
                           A(20) => RB(20), A(19) => RB(19), A(18) => RB(18), 
                           A(17) => RB(17), A(16) => RB(16), A(15) => RB(15), 
                           A(14) => RB(14), A(13) => RB(13), A(12) => RB(12), 
                           A(11) => RB(11), A(10) => RB(10), A(9) => RB(9), 
                           A(8) => RB(8), A(7) => RB(7), A(6) => RB(6), A(5) =>
                           RB(5), A(4) => RB(4), A(3) => RB(3), A(2) => RB(2), 
                           A(1) => RB(1), A(0) => RB(0), B(31) => IMM(31), 
                           B(30) => IMM(30), B(29) => IMM(29), B(28) => IMM(28)
                           , B(27) => IMM(27), B(26) => IMM(26), B(25) => 
                           IMM(25), B(24) => IMM(24), B(23) => IMM(23), B(22) 
                           => IMM(22), B(21) => IMM(21), B(20) => IMM(20), 
                           B(19) => IMM(19), B(18) => IMM(18), B(17) => IMM(17)
                           , B(16) => IMM(16), B(15) => IMM(15), B(14) => 
                           IMM(14), B(13) => IMM(13), B(12) => IMM(12), B(11) 
                           => IMM(11), B(10) => IMM(10), B(9) => IMM(9), B(8) 
                           => IMM(8), B(7) => IMM(7), B(6) => IMM(6), B(5) => 
                           IMM(5), B(4) => IMM(4), B(3) => IMM(3), B(2) => 
                           IMM(2), B(1) => IMM(1), B(0) => IMM(0), C(31) => 
                           ALU_outmem(31), C(30) => ALU_outmem(30), C(29) => 
                           ALU_outmem(29), C(28) => ALU_outmem(28), C(27) => 
                           ALU_outmem(27), C(26) => ALU_outmem(26), C(25) => 
                           ALU_outmem(25), C(24) => ALU_outmem(24), C(23) => 
                           ALU_outmem(23), C(22) => ALU_outmem(22), C(21) => 
                           ALU_outmem(21), C(20) => ALU_outmem(20), C(19) => 
                           ALU_outmem(19), C(18) => ALU_outmem(18), C(17) => 
                           ALU_outmem(17), C(16) => ALU_outmem(16), C(15) => 
                           ALU_outmem(15), C(14) => ALU_outmem(14), C(13) => 
                           ALU_outmem(13), C(12) => ALU_outmem(12), C(11) => 
                           ALU_outmem(11), C(10) => ALU_outmem(10), C(9) => 
                           ALU_outmem(9), C(8) => ALU_outmem(8), C(7) => 
                           ALU_outmem(7), C(6) => ALU_outmem(6), C(5) => 
                           ALU_outmem(5), C(4) => ALU_outmem(4), C(3) => 
                           ALU_outmem(3), C(2) => ALU_outmem(2), C(1) => 
                           ALU_outmem(1), C(0) => ALU_outmem(0), D(31) => 
                           WB_out(31), D(30) => WB_out(30), D(29) => WB_out(29)
                           , D(28) => WB_out(28), D(27) => WB_out(27), D(26) =>
                           WB_out(26), D(25) => WB_out(25), D(24) => WB_out(24)
                           , D(23) => WB_out(23), D(22) => WB_out(22), D(21) =>
                           WB_out(21), D(20) => WB_out(20), D(19) => WB_out(19)
                           , D(18) => WB_out(18), D(17) => WB_out(17), D(16) =>
                           WB_out(16), D(15) => WB_out(15), D(14) => WB_out(14)
                           , D(13) => WB_out(13), D(12) => WB_out(12), D(11) =>
                           WB_out(11), D(10) => WB_out(10), D(9) => WB_out(9), 
                           D(8) => WB_out(8), D(7) => WB_out(7), D(6) => 
                           WB_out(6), D(5) => WB_out(5), D(4) => WB_out(4), 
                           D(3) => WB_out(3), D(2) => WB_out(2), D(1) => 
                           WB_out(1), D(0) => WB_out(0), SEL(1) => s_S2_1_port,
                           SEL(0) => s_S2_0_port, Y(31) => MUX2out_31_port, 
                           Y(30) => MUX2out_30_port, Y(29) => MUX2out_29_port, 
                           Y(28) => MUX2out_28_port, Y(27) => MUX2out_27_port, 
                           Y(26) => MUX2out_26_port, Y(25) => MUX2out_25_port, 
                           Y(24) => MUX2out_24_port, Y(23) => MUX2out_23_port, 
                           Y(22) => MUX2out_22_port, Y(21) => MUX2out_21_port, 
                           Y(20) => MUX2out_20_port, Y(19) => MUX2out_19_port, 
                           Y(18) => MUX2out_18_port, Y(17) => MUX2out_17_port, 
                           Y(16) => MUX2out_16_port, Y(15) => MUX2out_15_port, 
                           Y(14) => MUX2out_14_port, Y(13) => MUX2out_13_port, 
                           Y(12) => MUX2out_12_port, Y(11) => MUX2out_11_port, 
                           Y(10) => MUX2out_10_port, Y(9) => MUX2out_9_port, 
                           Y(8) => MUX2out_8_port, Y(7) => MUX2out_7_port, Y(6)
                           => MUX2out_6_port, Y(5) => MUX2out_5_port, Y(4) => 
                           MUX2out_4_port, Y(3) => MUX2out_3_port, Y(2) => 
                           MUX2out_2_port, Y(1) => MUX2out_1_port, Y(0) => 
                           MUX2out_0_port);
   FW_MUX3 : MUX41_GENERIC_NBIT32_1 port map( A(31) => IMM(31), A(30) => 
                           IMM(30), A(29) => IMM(29), A(28) => IMM(28), A(27) 
                           => IMM(27), A(26) => IMM(26), A(25) => IMM(25), 
                           A(24) => IMM(24), A(23) => IMM(23), A(22) => IMM(22)
                           , A(21) => IMM(21), A(20) => IMM(20), A(19) => 
                           IMM(19), A(18) => IMM(18), A(17) => IMM(17), A(16) 
                           => IMM(16), A(15) => IMM(15), A(14) => IMM(14), 
                           A(13) => IMM(13), A(12) => IMM(12), A(11) => IMM(11)
                           , A(10) => IMM(10), A(9) => IMM(9), A(8) => IMM(8), 
                           A(7) => IMM(7), A(6) => IMM(6), A(5) => IMM(5), A(4)
                           => IMM(4), A(3) => IMM(3), A(2) => IMM(2), A(1) => 
                           IMM(1), A(0) => IMM(0), B(31) => RB(31), B(30) => 
                           RB(30), B(29) => RB(29), B(28) => RB(28), B(27) => 
                           RB(27), B(26) => RB(26), B(25) => RB(25), B(24) => 
                           RB(24), B(23) => RB(23), B(22) => RB(22), B(21) => 
                           RB(21), B(20) => RB(20), B(19) => RB(19), B(18) => 
                           RB(18), B(17) => RB(17), B(16) => RB(16), B(15) => 
                           RB(15), B(14) => RB(14), B(13) => RB(13), B(12) => 
                           RB(12), B(11) => RB(11), B(10) => RB(10), B(9) => 
                           RB(9), B(8) => RB(8), B(7) => RB(7), B(6) => RB(6), 
                           B(5) => RB(5), B(4) => RB(4), B(3) => RB(3), B(2) =>
                           RB(2), B(1) => RB(1), B(0) => RB(0), C(31) => 
                           ALU_outmem(31), C(30) => ALU_outmem(30), C(29) => 
                           ALU_outmem(29), C(28) => ALU_outmem(28), C(27) => 
                           ALU_outmem(27), C(26) => ALU_outmem(26), C(25) => 
                           ALU_outmem(25), C(24) => ALU_outmem(24), C(23) => 
                           ALU_outmem(23), C(22) => ALU_outmem(22), C(21) => 
                           ALU_outmem(21), C(20) => ALU_outmem(20), C(19) => 
                           ALU_outmem(19), C(18) => ALU_outmem(18), C(17) => 
                           ALU_outmem(17), C(16) => ALU_outmem(16), C(15) => 
                           ALU_outmem(15), C(14) => ALU_outmem(14), C(13) => 
                           ALU_outmem(13), C(12) => ALU_outmem(12), C(11) => 
                           ALU_outmem(11), C(10) => ALU_outmem(10), C(9) => 
                           ALU_outmem(9), C(8) => ALU_outmem(8), C(7) => 
                           ALU_outmem(7), C(6) => ALU_outmem(6), C(5) => 
                           ALU_outmem(5), C(4) => ALU_outmem(4), C(3) => 
                           ALU_outmem(3), C(2) => ALU_outmem(2), C(1) => 
                           ALU_outmem(1), C(0) => ALU_outmem(0), D(31) => 
                           WB_out(31), D(30) => WB_out(30), D(29) => WB_out(29)
                           , D(28) => WB_out(28), D(27) => WB_out(27), D(26) =>
                           WB_out(26), D(25) => WB_out(25), D(24) => WB_out(24)
                           , D(23) => WB_out(23), D(22) => WB_out(22), D(21) =>
                           WB_out(21), D(20) => WB_out(20), D(19) => WB_out(19)
                           , D(18) => WB_out(18), D(17) => WB_out(17), D(16) =>
                           WB_out(16), D(15) => WB_out(15), D(14) => WB_out(14)
                           , D(13) => WB_out(13), D(12) => WB_out(12), D(11) =>
                           WB_out(11), D(10) => WB_out(10), D(9) => WB_out(9), 
                           D(8) => WB_out(8), D(7) => WB_out(7), D(6) => 
                           WB_out(6), D(5) => WB_out(5), D(4) => WB_out(4), 
                           D(3) => WB_out(3), D(2) => WB_out(2), D(1) => 
                           WB_out(1), D(0) => WB_out(0), SEL(1) => s_S3_1_port,
                           SEL(0) => s_S3_0_port, Y(31) => ME(31), Y(30) => 
                           ME(30), Y(29) => ME(29), Y(28) => ME(28), Y(27) => 
                           ME(27), Y(26) => ME(26), Y(25) => ME(25), Y(24) => 
                           ME(24), Y(23) => ME(23), Y(22) => ME(22), Y(21) => 
                           ME(21), Y(20) => ME(20), Y(19) => ME(19), Y(18) => 
                           ME(18), Y(17) => ME(17), Y(16) => ME(16), Y(15) => 
                           ME(15), Y(14) => ME(14), Y(13) => ME(13), Y(12) => 
                           ME(12), Y(11) => ME(11), Y(10) => ME(10), Y(9) => 
                           ME(9), Y(8) => ME(8), Y(7) => ME(7), Y(6) => ME(6), 
                           Y(5) => ME(5), Y(4) => ME(4), Y(3) => ME(3), Y(2) =>
                           ME(2), Y(1) => ME(1), Y(0) => ME(0));
   RD_MUX1 : MUX21_GENERIC_NBIT5_0 port map( A(4) => WA(4), A(3) => WA(3), A(2)
                           => WA(2), A(1) => WA(1), A(0) => WA(0), B(4) => 
                           X_Logic0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           X_Logic0_port, SEL => N4, Y(4) => s_ALU_RD_4_port, 
                           Y(3) => s_ALU_RD_3_port, Y(2) => s_ALU_RD_2_port, 
                           Y(1) => s_ALU_RD_1_port, Y(0) => s_ALU_RD_0_port);
   EXUx : EXU_N32 port map( DATA1(31) => MUX1out_31_port, DATA1(30) => 
                           MUX1out_30_port, DATA1(29) => MUX1out_29_port, 
                           DATA1(28) => MUX1out_28_port, DATA1(27) => 
                           MUX1out_27_port, DATA1(26) => MUX1out_26_port, 
                           DATA1(25) => MUX1out_25_port, DATA1(24) => 
                           MUX1out_24_port, DATA1(23) => MUX1out_23_port, 
                           DATA1(22) => MUX1out_22_port, DATA1(21) => 
                           MUX1out_21_port, DATA1(20) => MUX1out_20_port, 
                           DATA1(19) => MUX1out_19_port, DATA1(18) => 
                           MUX1out_18_port, DATA1(17) => MUX1out_17_port, 
                           DATA1(16) => MUX1out_16_port, DATA1(15) => 
                           MUX1out_15_port, DATA1(14) => MUX1out_14_port, 
                           DATA1(13) => MUX1out_13_port, DATA1(12) => 
                           MUX1out_12_port, DATA1(11) => MUX1out_11_port, 
                           DATA1(10) => MUX1out_10_port, DATA1(9) => 
                           MUX1out_9_port, DATA1(8) => MUX1out_8_port, DATA1(7)
                           => MUX1out_7_port, DATA1(6) => MUX1out_6_port, 
                           DATA1(5) => MUX1out_5_port, DATA1(4) => 
                           MUX1out_4_port, DATA1(3) => MUX1out_3_port, DATA1(2)
                           => MUX1out_2_port, DATA1(1) => MUX1out_1_port, 
                           DATA1(0) => MUX1out_0_port, DATA2(31) => 
                           MUX2out_31_port, DATA2(30) => MUX2out_30_port, 
                           DATA2(29) => MUX2out_29_port, DATA2(28) => 
                           MUX2out_28_port, DATA2(27) => MUX2out_27_port, 
                           DATA2(26) => MUX2out_26_port, DATA2(25) => 
                           MUX2out_25_port, DATA2(24) => MUX2out_24_port, 
                           DATA2(23) => MUX2out_23_port, DATA2(22) => 
                           MUX2out_22_port, DATA2(21) => MUX2out_21_port, 
                           DATA2(20) => MUX2out_20_port, DATA2(19) => 
                           MUX2out_19_port, DATA2(18) => MUX2out_18_port, 
                           DATA2(17) => MUX2out_17_port, DATA2(16) => 
                           MUX2out_16_port, DATA2(15) => MUX2out_15_port, 
                           DATA2(14) => MUX2out_14_port, DATA2(13) => 
                           MUX2out_13_port, DATA2(12) => MUX2out_12_port, 
                           DATA2(11) => MUX2out_11_port, DATA2(10) => 
                           MUX2out_10_port, DATA2(9) => MUX2out_9_port, 
                           DATA2(8) => MUX2out_8_port, DATA2(7) => 
                           MUX2out_7_port, DATA2(6) => MUX2out_6_port, DATA2(5)
                           => MUX2out_5_port, DATA2(4) => MUX2out_4_port, 
                           DATA2(3) => MUX2out_3_port, DATA2(2) => 
                           MUX2out_2_port, DATA2(1) => MUX2out_1_port, DATA2(0)
                           => MUX2out_0_port, FUNC(3) => ALU3, FUNC(2) => ALU2,
                           FUNC(1) => ALU1, FUNC(0) => ALU0, RD_in(4) => WA(4),
                           RD_in(3) => WA(3), RD_in(2) => WA(2), RD_in(1) => 
                           WA(1), RD_in(0) => WA(0), SN => SN, CLK => CLK, RST 
                           => RST, OVF => s_ovf, stall_flag => flag_structHzd, 
                           RD_sel_flag => s_RD_sel2, OUTPUT(31) => output(31), 
                           OUTPUT(30) => output(30), OUTPUT(29) => output(29), 
                           OUTPUT(28) => output(28), OUTPUT(27) => output(27), 
                           OUTPUT(26) => output(26), OUTPUT(25) => output(25), 
                           OUTPUT(24) => output(24), OUTPUT(23) => output(23), 
                           OUTPUT(22) => output(22), OUTPUT(21) => output(21), 
                           OUTPUT(20) => output(20), OUTPUT(19) => output(19), 
                           OUTPUT(18) => output(18), OUTPUT(17) => output(17), 
                           OUTPUT(16) => output(16), OUTPUT(15) => output(15), 
                           OUTPUT(14) => output(14), OUTPUT(13) => output(13), 
                           OUTPUT(12) => output(12), OUTPUT(11) => output(11), 
                           OUTPUT(10) => output(10), OUTPUT(9) => output(9), 
                           OUTPUT(8) => output(8), OUTPUT(7) => output(7), 
                           OUTPUT(6) => output(6), OUTPUT(5) => output(5), 
                           OUTPUT(4) => output(4), OUTPUT(3) => output(3), 
                           OUTPUT(2) => output(2), OUTPUT(1) => output(1), 
                           OUTPUT(0) => output(0), RD_stall(4) => RD_inmul(4), 
                           RD_stall(3) => RD_inmul(3), RD_stall(2) => 
                           RD_inmul(2), RD_stall(1) => RD_inmul(1), RD_stall(0)
                           => RD_inmul(0), RD_out(4) => s_mul_RD_out_4_port, 
                           RD_out(3) => s_mul_RD_out_3_port, RD_out(2) => 
                           s_mul_RD_out_2_port, RD_out(1) => 
                           s_mul_RD_out_1_port, RD_out(0) => 
                           s_mul_RD_out_0_port, H_MULOUT(31) => n_1943, 
                           H_MULOUT(30) => n_1944, H_MULOUT(29) => n_1945, 
                           H_MULOUT(28) => n_1946, H_MULOUT(27) => n_1947, 
                           H_MULOUT(26) => n_1948, H_MULOUT(25) => n_1949, 
                           H_MULOUT(24) => n_1950, H_MULOUT(23) => n_1951, 
                           H_MULOUT(22) => n_1952, H_MULOUT(21) => n_1953, 
                           H_MULOUT(20) => n_1954, H_MULOUT(19) => n_1955, 
                           H_MULOUT(18) => n_1956, H_MULOUT(17) => n_1957, 
                           H_MULOUT(16) => n_1958, H_MULOUT(15) => n_1959, 
                           H_MULOUT(14) => n_1960, H_MULOUT(13) => n_1961, 
                           H_MULOUT(12) => n_1962, H_MULOUT(11) => n_1963, 
                           H_MULOUT(10) => n_1964, H_MULOUT(9) => n_1965, 
                           H_MULOUT(8) => n_1966, H_MULOUT(7) => n_1967, 
                           H_MULOUT(6) => n_1968, H_MULOUT(5) => n_1969, 
                           H_MULOUT(4) => n_1970, H_MULOUT(3) => n_1971, 
                           H_MULOUT(2) => n_1972, H_MULOUT(1) => n_1973, 
                           H_MULOUT(0) => n_1974);
   RD_MUX2 : MUX21_GENERIC_NBIT5_1 port map( A(4) => s_ALU_RD_4_port, A(3) => 
                           s_ALU_RD_3_port, A(2) => s_ALU_RD_2_port, A(1) => 
                           s_ALU_RD_1_port, A(0) => s_ALU_RD_0_port, B(4) => 
                           s_mul_RD_out_4_port, B(3) => s_mul_RD_out_3_port, 
                           B(2) => s_mul_RD_out_2_port, B(1) => 
                           s_mul_RD_out_1_port, B(0) => s_mul_RD_out_0_port, 
                           SEL => s_RD_sel2, Y(4) => WAout(4), Y(3) => WAout(3)
                           , Y(2) => WAout(2), Y(1) => WAout(1), Y(0) => 
                           WAout(0));
   U2 : AND2_X1 port map( A1 => s_ovf, A2 => SN, ZN => OVF);
   U3 : AND4_X1 port map( A1 => ALU3, A2 => ALU2, A3 => ALU1, A4 => ALU0, ZN =>
                           N4);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity DEC is

   port( instr : in std_logic_vector (31 downto 0);  RST : in std_logic;  
         RFdata_in : in std_logic_vector (31 downto 0);  RFWA : in 
         std_logic_vector (4 downto 0);  NPC_in : in std_logic_vector (31 
         downto 0);  EXE_RD : in std_logic_vector (4 downto 0);  Ld : in 
         std_logic;  ALU_regout : in std_logic_vector (31 downto 0);  MEM_RD, 
         WB_RD, RD_inmul : in std_logic_vector (4 downto 0);  flag_structHzd, 
         flag_ismul, RF1, RF2, WF1, EN1 : in std_logic;  opcode : out 
         std_logic_vector (5 downto 0);  func : out std_logic_vector (10 downto
         0);  IMM, RA, RB : out std_logic_vector (31 downto 0);  RSA, RSB, RD :
         out std_logic_vector (4 downto 0);  stall_NPC : out std_logic_vector 
         (31 downto 0);  PC_sel, dec_flag : out std_logic;  NPC_jump : out 
         std_logic_vector (31 downto 0));

end DEC;

architecture SYN_Behavioral of DEC is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component register_file_NBIT32_NREG32
      port( RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
            ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
            std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component 
      stall_detection_unit_op_code_size6_func_size11_PC_reg_size32_reg_file_size32
      port( opcode : in std_logic_vector (5 downto 0);  RSA, RSB, RD : in 
            std_logic_vector (4 downto 0);  FUNC : in std_logic_vector (10 
            downto 0);  EXE_RD : in std_logic_vector (4 downto 0);  NPC_in : in
            std_logic_vector (31 downto 0);  Ld : in std_logic;  RD_inmul : in 
            std_logic_vector (4 downto 0);  flag_structHzd, flag_ismul : in 
            std_logic;  opcode_out : out std_logic_vector (5 downto 0);  RD_out
            : out std_logic_vector (4 downto 0);  FUNC_out : out 
            std_logic_vector (10 downto 0);  NPC_out : out std_logic_vector (31
            downto 0);  PC_sel : out std_logic);
   end component;
   
   component MUX21_GENERIC_NBIT32_3
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component jump_logic_WORD_size32_NREG32_reg_file_size32
      port( opcode : in std_logic_vector (5 downto 0);  RSA, WB_RD, MEM_RD : in
            std_logic_vector (4 downto 0);  Rega, ALU_out, MEM_out : in 
            std_logic_vector (31 downto 0);  Rega_new : out std_logic_vector 
            (31 downto 0);  mux_s, flag : out std_logic);
   end component;
   
   component P4_ADDER_NBIT32_0
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  S :
            out std_logic_vector (31 downto 0);  Cout, ovf : out std_logic);
   end component;
   
   component dec_logic_WORD_size32_NREG32
      port( instr, NPC_in : in std_logic_vector (31 downto 0);  opcode : out 
            std_logic_vector (5 downto 0);  RS1, RS2, RD : out std_logic_vector
            (4 downto 0);  FUNC : out std_logic_vector (10 downto 0);  IMM : 
            out std_logic_vector (15 downto 0);  IMM26 : out std_logic_vector 
            (25 downto 0));
   end component;
   
   signal X_Logic0_port, opcode_5_port, opcode_4_port, opcode_3_port, 
      opcode_2_port, opcode_1_port, opcode_0_port, IMM_31_port, IMM_15_port, 
      IMM_14_port, IMM_13_port, IMM_12_port, IMM_11_port, IMM_10_port, 
      IMM_9_port, IMM_8_port, IMM_7_port, IMM_6_port, IMM_5_port, IMM_4_port, 
      IMM_3_port, IMM_2_port, IMM_1_port, IMM_0_port, RA_31_port, RA_30_port, 
      RA_29_port, RA_28_port, RA_27_port, RA_26_port, RA_25_port, RA_24_port, 
      RA_23_port, RA_22_port, RA_21_port, RA_20_port, RA_19_port, RA_18_port, 
      RA_17_port, RA_16_port, RA_15_port, RA_14_port, RA_13_port, RA_12_port, 
      RA_11_port, RA_10_port, RA_9_port, RA_8_port, RA_7_port, RA_6_port, 
      RA_5_port, RA_4_port, RA_3_port, RA_2_port, RA_1_port, RA_0_port, 
      RSA_4_port, RSA_3_port, RSA_2_port, RSA_1_port, RSA_0_port, RSB_4_port, 
      RSB_3_port, RSB_2_port, RSB_1_port, RSB_0_port, s_opcode_5_port, 
      s_opcode_4_port, s_opcode_3_port, s_opcode_2_port, s_opcode_1_port, 
      s_opcode_0_port, s_FUNC_10_port, s_FUNC_9_port, s_FUNC_8_port, 
      s_FUNC_7_port, s_FUNC_6_port, s_FUNC_5_port, s_FUNC_4_port, s_FUNC_3_port
      , s_FUNC_2_port, s_FUNC_1_port, s_FUNC_0_port, s_RD_4_port, s_RD_3_port, 
      s_RD_2_port, s_RD_1_port, s_RD_0_port, s_IMM26_25_port, s_IMM26_24_port, 
      s_IMM26_23_port, s_IMM26_22_port, s_IMM26_21_port, s_IMM26_20_port, 
      s_IMM26_19_port, s_IMM26_18_port, s_IMM26_17_port, s_IMM26_16_port, 
      s_IMM26_15_port, s_IMM26_14_port, s_IMM26_13_port, s_IMM26_12_port, 
      s_IMM26_11_port, s_IMM26_10_port, s_IMM26_9_port, s_IMM26_8_port, 
      s_IMM26_7_port, s_IMM26_6_port, s_IMM26_5_port, s_IMM26_4_port, 
      s_IMM26_3_port, s_IMM26_2_port, s_IMM26_1_port, s_IMM26_0_port, 
      adder_out_31_port, adder_out_30_port, adder_out_29_port, 
      adder_out_28_port, adder_out_27_port, adder_out_26_port, 
      adder_out_25_port, adder_out_24_port, adder_out_23_port, 
      adder_out_22_port, adder_out_21_port, adder_out_20_port, 
      adder_out_19_port, adder_out_18_port, adder_out_17_port, 
      adder_out_16_port, adder_out_15_port, adder_out_14_port, 
      adder_out_13_port, adder_out_12_port, adder_out_11_port, 
      adder_out_10_port, adder_out_9_port, adder_out_8_port, adder_out_7_port, 
      adder_out_6_port, adder_out_5_port, adder_out_4_port, adder_out_3_port, 
      adder_out_2_port, adder_out_1_port, adder_out_0_port, s_Rega_new_31_port,
      s_Rega_new_30_port, s_Rega_new_29_port, s_Rega_new_28_port, 
      s_Rega_new_27_port, s_Rega_new_26_port, s_Rega_new_25_port, 
      s_Rega_new_24_port, s_Rega_new_23_port, s_Rega_new_22_port, 
      s_Rega_new_21_port, s_Rega_new_20_port, s_Rega_new_19_port, 
      s_Rega_new_18_port, s_Rega_new_17_port, s_Rega_new_16_port, 
      s_Rega_new_15_port, s_Rega_new_14_port, s_Rega_new_13_port, 
      s_Rega_new_12_port, s_Rega_new_11_port, s_Rega_new_10_port, 
      s_Rega_new_9_port, s_Rega_new_8_port, s_Rega_new_7_port, 
      s_Rega_new_6_port, s_Rega_new_5_port, s_Rega_new_4_port, 
      s_Rega_new_3_port, s_Rega_new_2_port, s_Rega_new_1_port, 
      s_Rega_new_0_port, mux_select, n3, n4, n5, n6, n7, n1, n2, n8, n9, n_1975
      , n_1976 : std_logic;

begin
   opcode <= ( opcode_5_port, opcode_4_port, opcode_3_port, opcode_2_port, 
      opcode_1_port, opcode_0_port );
   IMM <= ( IMM_31_port, IMM_31_port, IMM_31_port, IMM_31_port, IMM_31_port, 
      IMM_31_port, IMM_31_port, IMM_31_port, IMM_31_port, IMM_31_port, 
      IMM_31_port, IMM_31_port, IMM_31_port, IMM_31_port, IMM_31_port, 
      IMM_31_port, IMM_15_port, IMM_14_port, IMM_13_port, IMM_12_port, 
      IMM_11_port, IMM_10_port, IMM_9_port, IMM_8_port, IMM_7_port, IMM_6_port,
      IMM_5_port, IMM_4_port, IMM_3_port, IMM_2_port, IMM_1_port, IMM_0_port );
   RA <= ( RA_31_port, RA_30_port, RA_29_port, RA_28_port, RA_27_port, 
      RA_26_port, RA_25_port, RA_24_port, RA_23_port, RA_22_port, RA_21_port, 
      RA_20_port, RA_19_port, RA_18_port, RA_17_port, RA_16_port, RA_15_port, 
      RA_14_port, RA_13_port, RA_12_port, RA_11_port, RA_10_port, RA_9_port, 
      RA_8_port, RA_7_port, RA_6_port, RA_5_port, RA_4_port, RA_3_port, 
      RA_2_port, RA_1_port, RA_0_port );
   RSA <= ( RSA_4_port, RSA_3_port, RSA_2_port, RSA_1_port, RSA_0_port );
   RSB <= ( RSB_4_port, RSB_3_port, RSB_2_port, RSB_1_port, RSB_0_port );
   
   X_Logic0_port <= '0';
   decode_logic : dec_logic_WORD_size32_NREG32 port map( instr(31) => instr(31)
                           , instr(30) => instr(30), instr(29) => instr(29), 
                           instr(28) => instr(28), instr(27) => instr(27), 
                           instr(26) => instr(26), instr(25) => instr(25), 
                           instr(24) => instr(24), instr(23) => instr(23), 
                           instr(22) => instr(22), instr(21) => instr(21), 
                           instr(20) => instr(20), instr(19) => instr(19), 
                           instr(18) => instr(18), instr(17) => instr(17), 
                           instr(16) => instr(16), instr(15) => instr(15), 
                           instr(14) => instr(14), instr(13) => instr(13), 
                           instr(12) => instr(12), instr(11) => instr(11), 
                           instr(10) => instr(10), instr(9) => instr(9), 
                           instr(8) => instr(8), instr(7) => instr(7), instr(6)
                           => instr(6), instr(5) => instr(5), instr(4) => 
                           instr(4), instr(3) => instr(3), instr(2) => instr(2)
                           , instr(1) => instr(1), instr(0) => instr(0), 
                           NPC_in(31) => NPC_in(31), NPC_in(30) => NPC_in(30), 
                           NPC_in(29) => NPC_in(29), NPC_in(28) => NPC_in(28), 
                           NPC_in(27) => NPC_in(27), NPC_in(26) => NPC_in(26), 
                           NPC_in(25) => NPC_in(25), NPC_in(24) => NPC_in(24), 
                           NPC_in(23) => NPC_in(23), NPC_in(22) => NPC_in(22), 
                           NPC_in(21) => NPC_in(21), NPC_in(20) => NPC_in(20), 
                           NPC_in(19) => NPC_in(19), NPC_in(18) => NPC_in(18), 
                           NPC_in(17) => NPC_in(17), NPC_in(16) => NPC_in(16), 
                           NPC_in(15) => NPC_in(15), NPC_in(14) => NPC_in(14), 
                           NPC_in(13) => NPC_in(13), NPC_in(12) => NPC_in(12), 
                           NPC_in(11) => NPC_in(11), NPC_in(10) => NPC_in(10), 
                           NPC_in(9) => NPC_in(9), NPC_in(8) => NPC_in(8), 
                           NPC_in(7) => NPC_in(7), NPC_in(6) => NPC_in(6), 
                           NPC_in(5) => NPC_in(5), NPC_in(4) => NPC_in(4), 
                           NPC_in(3) => NPC_in(3), NPC_in(2) => NPC_in(2), 
                           NPC_in(1) => NPC_in(1), NPC_in(0) => NPC_in(0), 
                           opcode(5) => s_opcode_5_port, opcode(4) => 
                           s_opcode_4_port, opcode(3) => s_opcode_3_port, 
                           opcode(2) => s_opcode_2_port, opcode(1) => 
                           s_opcode_1_port, opcode(0) => s_opcode_0_port, 
                           RS1(4) => RSA_4_port, RS1(3) => RSA_3_port, RS1(2) 
                           => RSA_2_port, RS1(1) => RSA_1_port, RS1(0) => 
                           RSA_0_port, RS2(4) => RSB_4_port, RS2(3) => 
                           RSB_3_port, RS2(2) => RSB_2_port, RS2(1) => 
                           RSB_1_port, RS2(0) => RSB_0_port, RD(4) => 
                           s_RD_4_port, RD(3) => s_RD_3_port, RD(2) => 
                           s_RD_2_port, RD(1) => s_RD_1_port, RD(0) => 
                           s_RD_0_port, FUNC(10) => s_FUNC_10_port, FUNC(9) => 
                           s_FUNC_9_port, FUNC(8) => s_FUNC_8_port, FUNC(7) => 
                           s_FUNC_7_port, FUNC(6) => s_FUNC_6_port, FUNC(5) => 
                           s_FUNC_5_port, FUNC(4) => s_FUNC_4_port, FUNC(3) => 
                           s_FUNC_3_port, FUNC(2) => s_FUNC_2_port, FUNC(1) => 
                           s_FUNC_1_port, FUNC(0) => s_FUNC_0_port, IMM(15) => 
                           IMM_15_port, IMM(14) => IMM_14_port, IMM(13) => 
                           IMM_13_port, IMM(12) => IMM_12_port, IMM(11) => 
                           IMM_11_port, IMM(10) => IMM_10_port, IMM(9) => 
                           IMM_9_port, IMM(8) => IMM_8_port, IMM(7) => 
                           IMM_7_port, IMM(6) => IMM_6_port, IMM(5) => 
                           IMM_5_port, IMM(4) => IMM_4_port, IMM(3) => 
                           IMM_3_port, IMM(2) => IMM_2_port, IMM(1) => 
                           IMM_1_port, IMM(0) => IMM_0_port, IMM26(25) => 
                           s_IMM26_25_port, IMM26(24) => s_IMM26_24_port, 
                           IMM26(23) => s_IMM26_23_port, IMM26(22) => 
                           s_IMM26_22_port, IMM26(21) => s_IMM26_21_port, 
                           IMM26(20) => s_IMM26_20_port, IMM26(19) => 
                           s_IMM26_19_port, IMM26(18) => s_IMM26_18_port, 
                           IMM26(17) => s_IMM26_17_port, IMM26(16) => 
                           s_IMM26_16_port, IMM26(15) => s_IMM26_15_port, 
                           IMM26(14) => s_IMM26_14_port, IMM26(13) => 
                           s_IMM26_13_port, IMM26(12) => s_IMM26_12_port, 
                           IMM26(11) => s_IMM26_11_port, IMM26(10) => 
                           s_IMM26_10_port, IMM26(9) => s_IMM26_9_port, 
                           IMM26(8) => s_IMM26_8_port, IMM26(7) => 
                           s_IMM26_7_port, IMM26(6) => s_IMM26_6_port, IMM26(5)
                           => s_IMM26_5_port, IMM26(4) => s_IMM26_4_port, 
                           IMM26(3) => s_IMM26_3_port, IMM26(2) => 
                           s_IMM26_2_port, IMM26(1) => s_IMM26_1_port, IMM26(0)
                           => s_IMM26_0_port);
   jump_npc_adder : P4_ADDER_NBIT32_0 port map( A(31) => n1, A(30) => n1, A(29)
                           => n1, A(28) => n1, A(27) => n1, A(26) => n2, A(25) 
                           => n2, A(24) => s_IMM26_24_port, A(23) => 
                           s_IMM26_23_port, A(22) => s_IMM26_22_port, A(21) => 
                           s_IMM26_21_port, A(20) => s_IMM26_20_port, A(19) => 
                           s_IMM26_19_port, A(18) => s_IMM26_18_port, A(17) => 
                           s_IMM26_17_port, A(16) => s_IMM26_16_port, A(15) => 
                           s_IMM26_15_port, A(14) => s_IMM26_14_port, A(13) => 
                           s_IMM26_13_port, A(12) => s_IMM26_12_port, A(11) => 
                           s_IMM26_11_port, A(10) => s_IMM26_10_port, A(9) => 
                           s_IMM26_9_port, A(8) => s_IMM26_8_port, A(7) => 
                           s_IMM26_7_port, A(6) => s_IMM26_6_port, A(5) => 
                           s_IMM26_5_port, A(4) => s_IMM26_4_port, A(3) => 
                           s_IMM26_3_port, A(2) => s_IMM26_2_port, A(1) => 
                           s_IMM26_1_port, A(0) => s_IMM26_0_port, B(31) => 
                           NPC_in(31), B(30) => NPC_in(30), B(29) => NPC_in(29)
                           , B(28) => NPC_in(28), B(27) => NPC_in(27), B(26) =>
                           NPC_in(26), B(25) => NPC_in(25), B(24) => NPC_in(24)
                           , B(23) => NPC_in(23), B(22) => NPC_in(22), B(21) =>
                           NPC_in(21), B(20) => NPC_in(20), B(19) => NPC_in(19)
                           , B(18) => NPC_in(18), B(17) => NPC_in(17), B(16) =>
                           NPC_in(16), B(15) => NPC_in(15), B(14) => NPC_in(14)
                           , B(13) => NPC_in(13), B(12) => NPC_in(12), B(11) =>
                           NPC_in(11), B(10) => NPC_in(10), B(9) => NPC_in(9), 
                           B(8) => NPC_in(8), B(7) => NPC_in(7), B(6) => 
                           NPC_in(6), B(5) => NPC_in(5), B(4) => NPC_in(4), 
                           B(3) => NPC_in(3), B(2) => NPC_in(2), B(1) => 
                           NPC_in(1), B(0) => NPC_in(0), Cin => X_Logic0_port, 
                           S(31) => adder_out_31_port, S(30) => 
                           adder_out_30_port, S(29) => adder_out_29_port, S(28)
                           => adder_out_28_port, S(27) => adder_out_27_port, 
                           S(26) => adder_out_26_port, S(25) => 
                           adder_out_25_port, S(24) => adder_out_24_port, S(23)
                           => adder_out_23_port, S(22) => adder_out_22_port, 
                           S(21) => adder_out_21_port, S(20) => 
                           adder_out_20_port, S(19) => adder_out_19_port, S(18)
                           => adder_out_18_port, S(17) => adder_out_17_port, 
                           S(16) => adder_out_16_port, S(15) => 
                           adder_out_15_port, S(14) => adder_out_14_port, S(13)
                           => adder_out_13_port, S(12) => adder_out_12_port, 
                           S(11) => adder_out_11_port, S(10) => 
                           adder_out_10_port, S(9) => adder_out_9_port, S(8) =>
                           adder_out_8_port, S(7) => adder_out_7_port, S(6) => 
                           adder_out_6_port, S(5) => adder_out_5_port, S(4) => 
                           adder_out_4_port, S(3) => adder_out_3_port, S(2) => 
                           adder_out_2_port, S(1) => adder_out_1_port, S(0) => 
                           adder_out_0_port, Cout => n_1975, ovf => n_1976);
   jmp_logic : jump_logic_WORD_size32_NREG32_reg_file_size32 port map( 
                           opcode(5) => opcode_5_port, opcode(4) => 
                           opcode_4_port, opcode(3) => opcode_3_port, opcode(2)
                           => opcode_2_port, opcode(1) => opcode_1_port, 
                           opcode(0) => opcode_0_port, RSA(4) => RSA_4_port, 
                           RSA(3) => RSA_3_port, RSA(2) => RSA_2_port, RSA(1) 
                           => RSA_1_port, RSA(0) => RSA_0_port, WB_RD(4) => 
                           WB_RD(4), WB_RD(3) => WB_RD(3), WB_RD(2) => WB_RD(2)
                           , WB_RD(1) => WB_RD(1), WB_RD(0) => WB_RD(0), 
                           MEM_RD(4) => MEM_RD(4), MEM_RD(3) => MEM_RD(3), 
                           MEM_RD(2) => MEM_RD(2), MEM_RD(1) => MEM_RD(1), 
                           MEM_RD(0) => MEM_RD(0), Rega(31) => RA_31_port, 
                           Rega(30) => RA_30_port, Rega(29) => RA_29_port, 
                           Rega(28) => RA_28_port, Rega(27) => RA_27_port, 
                           Rega(26) => RA_26_port, Rega(25) => RA_25_port, 
                           Rega(24) => RA_24_port, Rega(23) => RA_23_port, 
                           Rega(22) => RA_22_port, Rega(21) => RA_21_port, 
                           Rega(20) => RA_20_port, Rega(19) => RA_19_port, 
                           Rega(18) => RA_18_port, Rega(17) => RA_17_port, 
                           Rega(16) => RA_16_port, Rega(15) => RA_15_port, 
                           Rega(14) => RA_14_port, Rega(13) => RA_13_port, 
                           Rega(12) => RA_12_port, Rega(11) => RA_11_port, 
                           Rega(10) => RA_10_port, Rega(9) => RA_9_port, 
                           Rega(8) => RA_8_port, Rega(7) => RA_7_port, Rega(6) 
                           => RA_6_port, Rega(5) => RA_5_port, Rega(4) => 
                           RA_4_port, Rega(3) => RA_3_port, Rega(2) => 
                           RA_2_port, Rega(1) => RA_1_port, Rega(0) => 
                           RA_0_port, ALU_out(31) => ALU_regout(31), 
                           ALU_out(30) => ALU_regout(30), ALU_out(29) => 
                           ALU_regout(29), ALU_out(28) => ALU_regout(28), 
                           ALU_out(27) => ALU_regout(27), ALU_out(26) => 
                           ALU_regout(26), ALU_out(25) => ALU_regout(25), 
                           ALU_out(24) => ALU_regout(24), ALU_out(23) => 
                           ALU_regout(23), ALU_out(22) => ALU_regout(22), 
                           ALU_out(21) => ALU_regout(21), ALU_out(20) => 
                           ALU_regout(20), ALU_out(19) => ALU_regout(19), 
                           ALU_out(18) => ALU_regout(18), ALU_out(17) => 
                           ALU_regout(17), ALU_out(16) => ALU_regout(16), 
                           ALU_out(15) => ALU_regout(15), ALU_out(14) => 
                           ALU_regout(14), ALU_out(13) => ALU_regout(13), 
                           ALU_out(12) => ALU_regout(12), ALU_out(11) => 
                           ALU_regout(11), ALU_out(10) => ALU_regout(10), 
                           ALU_out(9) => ALU_regout(9), ALU_out(8) => 
                           ALU_regout(8), ALU_out(7) => ALU_regout(7), 
                           ALU_out(6) => ALU_regout(6), ALU_out(5) => 
                           ALU_regout(5), ALU_out(4) => ALU_regout(4), 
                           ALU_out(3) => ALU_regout(3), ALU_out(2) => 
                           ALU_regout(2), ALU_out(1) => ALU_regout(1), 
                           ALU_out(0) => ALU_regout(0), MEM_out(31) => 
                           RFdata_in(31), MEM_out(30) => RFdata_in(30), 
                           MEM_out(29) => RFdata_in(29), MEM_out(28) => 
                           RFdata_in(28), MEM_out(27) => RFdata_in(27), 
                           MEM_out(26) => RFdata_in(26), MEM_out(25) => 
                           RFdata_in(25), MEM_out(24) => RFdata_in(24), 
                           MEM_out(23) => RFdata_in(23), MEM_out(22) => 
                           RFdata_in(22), MEM_out(21) => RFdata_in(21), 
                           MEM_out(20) => RFdata_in(20), MEM_out(19) => 
                           RFdata_in(19), MEM_out(18) => RFdata_in(18), 
                           MEM_out(17) => RFdata_in(17), MEM_out(16) => 
                           RFdata_in(16), MEM_out(15) => RFdata_in(15), 
                           MEM_out(14) => RFdata_in(14), MEM_out(13) => 
                           RFdata_in(13), MEM_out(12) => RFdata_in(12), 
                           MEM_out(11) => RFdata_in(11), MEM_out(10) => 
                           RFdata_in(10), MEM_out(9) => RFdata_in(9), 
                           MEM_out(8) => RFdata_in(8), MEM_out(7) => 
                           RFdata_in(7), MEM_out(6) => RFdata_in(6), MEM_out(5)
                           => RFdata_in(5), MEM_out(4) => RFdata_in(4), 
                           MEM_out(3) => RFdata_in(3), MEM_out(2) => 
                           RFdata_in(2), MEM_out(1) => RFdata_in(1), MEM_out(0)
                           => RFdata_in(0), Rega_new(31) => s_Rega_new_31_port,
                           Rega_new(30) => s_Rega_new_30_port, Rega_new(29) => 
                           s_Rega_new_29_port, Rega_new(28) => 
                           s_Rega_new_28_port, Rega_new(27) => 
                           s_Rega_new_27_port, Rega_new(26) => 
                           s_Rega_new_26_port, Rega_new(25) => 
                           s_Rega_new_25_port, Rega_new(24) => 
                           s_Rega_new_24_port, Rega_new(23) => 
                           s_Rega_new_23_port, Rega_new(22) => 
                           s_Rega_new_22_port, Rega_new(21) => 
                           s_Rega_new_21_port, Rega_new(20) => 
                           s_Rega_new_20_port, Rega_new(19) => 
                           s_Rega_new_19_port, Rega_new(18) => 
                           s_Rega_new_18_port, Rega_new(17) => 
                           s_Rega_new_17_port, Rega_new(16) => 
                           s_Rega_new_16_port, Rega_new(15) => 
                           s_Rega_new_15_port, Rega_new(14) => 
                           s_Rega_new_14_port, Rega_new(13) => 
                           s_Rega_new_13_port, Rega_new(12) => 
                           s_Rega_new_12_port, Rega_new(11) => 
                           s_Rega_new_11_port, Rega_new(10) => 
                           s_Rega_new_10_port, Rega_new(9) => s_Rega_new_9_port
                           , Rega_new(8) => s_Rega_new_8_port, Rega_new(7) => 
                           s_Rega_new_7_port, Rega_new(6) => s_Rega_new_6_port,
                           Rega_new(5) => s_Rega_new_5_port, Rega_new(4) => 
                           s_Rega_new_4_port, Rega_new(3) => s_Rega_new_3_port,
                           Rega_new(2) => s_Rega_new_2_port, Rega_new(1) => 
                           s_Rega_new_1_port, Rega_new(0) => s_Rega_new_0_port,
                           mux_s => mux_select, flag => dec_flag);
   MUX : MUX21_GENERIC_NBIT32_3 port map( A(31) => adder_out_31_port, A(30) => 
                           adder_out_30_port, A(29) => adder_out_29_port, A(28)
                           => adder_out_28_port, A(27) => adder_out_27_port, 
                           A(26) => adder_out_26_port, A(25) => 
                           adder_out_25_port, A(24) => adder_out_24_port, A(23)
                           => adder_out_23_port, A(22) => adder_out_22_port, 
                           A(21) => adder_out_21_port, A(20) => 
                           adder_out_20_port, A(19) => adder_out_19_port, A(18)
                           => adder_out_18_port, A(17) => adder_out_17_port, 
                           A(16) => adder_out_16_port, A(15) => 
                           adder_out_15_port, A(14) => adder_out_14_port, A(13)
                           => adder_out_13_port, A(12) => adder_out_12_port, 
                           A(11) => adder_out_11_port, A(10) => 
                           adder_out_10_port, A(9) => adder_out_9_port, A(8) =>
                           adder_out_8_port, A(7) => adder_out_7_port, A(6) => 
                           adder_out_6_port, A(5) => adder_out_5_port, A(4) => 
                           adder_out_4_port, A(3) => adder_out_3_port, A(2) => 
                           adder_out_2_port, A(1) => adder_out_1_port, A(0) => 
                           adder_out_0_port, B(31) => s_Rega_new_31_port, B(30)
                           => s_Rega_new_30_port, B(29) => s_Rega_new_29_port, 
                           B(28) => s_Rega_new_28_port, B(27) => 
                           s_Rega_new_27_port, B(26) => s_Rega_new_26_port, 
                           B(25) => s_Rega_new_25_port, B(24) => 
                           s_Rega_new_24_port, B(23) => s_Rega_new_23_port, 
                           B(22) => s_Rega_new_22_port, B(21) => 
                           s_Rega_new_21_port, B(20) => s_Rega_new_20_port, 
                           B(19) => s_Rega_new_19_port, B(18) => 
                           s_Rega_new_18_port, B(17) => s_Rega_new_17_port, 
                           B(16) => s_Rega_new_16_port, B(15) => 
                           s_Rega_new_15_port, B(14) => s_Rega_new_14_port, 
                           B(13) => s_Rega_new_13_port, B(12) => 
                           s_Rega_new_12_port, B(11) => s_Rega_new_11_port, 
                           B(10) => s_Rega_new_10_port, B(9) => 
                           s_Rega_new_9_port, B(8) => s_Rega_new_8_port, B(7) 
                           => s_Rega_new_7_port, B(6) => s_Rega_new_6_port, 
                           B(5) => s_Rega_new_5_port, B(4) => s_Rega_new_4_port
                           , B(3) => s_Rega_new_3_port, B(2) => 
                           s_Rega_new_2_port, B(1) => s_Rega_new_1_port, B(0) 
                           => s_Rega_new_0_port, SEL => mux_select, Y(31) => 
                           NPC_jump(31), Y(30) => NPC_jump(30), Y(29) => 
                           NPC_jump(29), Y(28) => NPC_jump(28), Y(27) => 
                           NPC_jump(27), Y(26) => NPC_jump(26), Y(25) => 
                           NPC_jump(25), Y(24) => NPC_jump(24), Y(23) => 
                           NPC_jump(23), Y(22) => NPC_jump(22), Y(21) => 
                           NPC_jump(21), Y(20) => NPC_jump(20), Y(19) => 
                           NPC_jump(19), Y(18) => NPC_jump(18), Y(17) => 
                           NPC_jump(17), Y(16) => NPC_jump(16), Y(15) => 
                           NPC_jump(15), Y(14) => NPC_jump(14), Y(13) => 
                           NPC_jump(13), Y(12) => NPC_jump(12), Y(11) => 
                           NPC_jump(11), Y(10) => NPC_jump(10), Y(9) => 
                           NPC_jump(9), Y(8) => NPC_jump(8), Y(7) => 
                           NPC_jump(7), Y(6) => NPC_jump(6), Y(5) => 
                           NPC_jump(5), Y(4) => NPC_jump(4), Y(3) => 
                           NPC_jump(3), Y(2) => NPC_jump(2), Y(1) => 
                           NPC_jump(1), Y(0) => NPC_jump(0));
   SDU : 
                           stall_detection_unit_op_code_size6_func_size11_PC_reg_size32_reg_file_size32 
                           port map( opcode(5) => s_opcode_5_port, opcode(4) =>
                           s_opcode_4_port, opcode(3) => s_opcode_3_port, 
                           opcode(2) => s_opcode_2_port, opcode(1) => 
                           s_opcode_1_port, opcode(0) => s_opcode_0_port, 
                           RSA(4) => RSA_4_port, RSA(3) => RSA_3_port, RSA(2) 
                           => RSA_2_port, RSA(1) => RSA_1_port, RSA(0) => 
                           RSA_0_port, RSB(4) => RSB_4_port, RSB(3) => 
                           RSB_3_port, RSB(2) => RSB_2_port, RSB(1) => 
                           RSB_1_port, RSB(0) => RSB_0_port, RD(4) => 
                           s_RD_4_port, RD(3) => s_RD_3_port, RD(2) => 
                           s_RD_2_port, RD(1) => s_RD_1_port, RD(0) => 
                           s_RD_0_port, FUNC(10) => s_FUNC_10_port, FUNC(9) => 
                           s_FUNC_9_port, FUNC(8) => s_FUNC_8_port, FUNC(7) => 
                           s_FUNC_7_port, FUNC(6) => s_FUNC_6_port, FUNC(5) => 
                           s_FUNC_5_port, FUNC(4) => s_FUNC_4_port, FUNC(3) => 
                           s_FUNC_3_port, FUNC(2) => s_FUNC_2_port, FUNC(1) => 
                           s_FUNC_1_port, FUNC(0) => s_FUNC_0_port, EXE_RD(4) 
                           => EXE_RD(4), EXE_RD(3) => EXE_RD(3), EXE_RD(2) => 
                           EXE_RD(2), EXE_RD(1) => EXE_RD(1), EXE_RD(0) => 
                           EXE_RD(0), NPC_in(31) => NPC_in(31), NPC_in(30) => 
                           NPC_in(30), NPC_in(29) => NPC_in(29), NPC_in(28) => 
                           NPC_in(28), NPC_in(27) => NPC_in(27), NPC_in(26) => 
                           NPC_in(26), NPC_in(25) => NPC_in(25), NPC_in(24) => 
                           NPC_in(24), NPC_in(23) => NPC_in(23), NPC_in(22) => 
                           NPC_in(22), NPC_in(21) => NPC_in(21), NPC_in(20) => 
                           NPC_in(20), NPC_in(19) => NPC_in(19), NPC_in(18) => 
                           NPC_in(18), NPC_in(17) => NPC_in(17), NPC_in(16) => 
                           NPC_in(16), NPC_in(15) => NPC_in(15), NPC_in(14) => 
                           NPC_in(14), NPC_in(13) => NPC_in(13), NPC_in(12) => 
                           NPC_in(12), NPC_in(11) => NPC_in(11), NPC_in(10) => 
                           NPC_in(10), NPC_in(9) => NPC_in(9), NPC_in(8) => 
                           NPC_in(8), NPC_in(7) => NPC_in(7), NPC_in(6) => 
                           NPC_in(6), NPC_in(5) => NPC_in(5), NPC_in(4) => 
                           NPC_in(4), NPC_in(3) => NPC_in(3), NPC_in(2) => 
                           NPC_in(2), NPC_in(1) => NPC_in(1), NPC_in(0) => 
                           NPC_in(0), Ld => Ld, RD_inmul(4) => RD_inmul(4), 
                           RD_inmul(3) => RD_inmul(3), RD_inmul(2) => 
                           RD_inmul(2), RD_inmul(1) => RD_inmul(1), RD_inmul(0)
                           => RD_inmul(0), flag_structHzd => flag_structHzd, 
                           flag_ismul => flag_ismul, opcode_out(5) => 
                           opcode_5_port, opcode_out(4) => opcode_4_port, 
                           opcode_out(3) => opcode_3_port, opcode_out(2) => 
                           opcode_2_port, opcode_out(1) => opcode_1_port, 
                           opcode_out(0) => opcode_0_port, RD_out(4) => RD(4), 
                           RD_out(3) => RD(3), RD_out(2) => RD(2), RD_out(1) =>
                           RD(1), RD_out(0) => RD(0), FUNC_out(10) => func(10),
                           FUNC_out(9) => func(9), FUNC_out(8) => func(8), 
                           FUNC_out(7) => func(7), FUNC_out(6) => func(6), 
                           FUNC_out(5) => func(5), FUNC_out(4) => func(4), 
                           FUNC_out(3) => func(3), FUNC_out(2) => func(2), 
                           FUNC_out(1) => func(1), FUNC_out(0) => func(0), 
                           NPC_out(31) => stall_NPC(31), NPC_out(30) => 
                           stall_NPC(30), NPC_out(29) => stall_NPC(29), 
                           NPC_out(28) => stall_NPC(28), NPC_out(27) => 
                           stall_NPC(27), NPC_out(26) => stall_NPC(26), 
                           NPC_out(25) => stall_NPC(25), NPC_out(24) => 
                           stall_NPC(24), NPC_out(23) => stall_NPC(23), 
                           NPC_out(22) => stall_NPC(22), NPC_out(21) => 
                           stall_NPC(21), NPC_out(20) => stall_NPC(20), 
                           NPC_out(19) => stall_NPC(19), NPC_out(18) => 
                           stall_NPC(18), NPC_out(17) => stall_NPC(17), 
                           NPC_out(16) => stall_NPC(16), NPC_out(15) => 
                           stall_NPC(15), NPC_out(14) => stall_NPC(14), 
                           NPC_out(13) => stall_NPC(13), NPC_out(12) => 
                           stall_NPC(12), NPC_out(11) => stall_NPC(11), 
                           NPC_out(10) => stall_NPC(10), NPC_out(9) => 
                           stall_NPC(9), NPC_out(8) => stall_NPC(8), NPC_out(7)
                           => stall_NPC(7), NPC_out(6) => stall_NPC(6), 
                           NPC_out(5) => stall_NPC(5), NPC_out(4) => 
                           stall_NPC(4), NPC_out(3) => stall_NPC(3), NPC_out(2)
                           => stall_NPC(2), NPC_out(1) => stall_NPC(1), 
                           NPC_out(0) => stall_NPC(0), PC_sel => PC_sel);
   REG_FILE : register_file_NBIT32_NREG32 port map( RESET => RST, ENABLE => EN1
                           , RD1 => RF1, RD2 => RF2, WR => WF1, ADD_WR(4) => 
                           RFWA(4), ADD_WR(3) => RFWA(3), ADD_WR(2) => RFWA(2),
                           ADD_WR(1) => RFWA(1), ADD_WR(0) => RFWA(0), 
                           ADD_RD1(4) => RSA_4_port, ADD_RD1(3) => RSA_3_port, 
                           ADD_RD1(2) => RSA_2_port, ADD_RD1(1) => RSA_1_port, 
                           ADD_RD1(0) => RSA_0_port, ADD_RD2(4) => RSB_4_port, 
                           ADD_RD2(3) => RSB_3_port, ADD_RD2(2) => RSB_2_port, 
                           ADD_RD2(1) => RSB_1_port, ADD_RD2(0) => RSB_0_port, 
                           DATAIN(31) => RFdata_in(31), DATAIN(30) => 
                           RFdata_in(30), DATAIN(29) => RFdata_in(29), 
                           DATAIN(28) => RFdata_in(28), DATAIN(27) => 
                           RFdata_in(27), DATAIN(26) => RFdata_in(26), 
                           DATAIN(25) => RFdata_in(25), DATAIN(24) => 
                           RFdata_in(24), DATAIN(23) => RFdata_in(23), 
                           DATAIN(22) => RFdata_in(22), DATAIN(21) => 
                           RFdata_in(21), DATAIN(20) => RFdata_in(20), 
                           DATAIN(19) => RFdata_in(19), DATAIN(18) => 
                           RFdata_in(18), DATAIN(17) => RFdata_in(17), 
                           DATAIN(16) => RFdata_in(16), DATAIN(15) => 
                           RFdata_in(15), DATAIN(14) => RFdata_in(14), 
                           DATAIN(13) => RFdata_in(13), DATAIN(12) => 
                           RFdata_in(12), DATAIN(11) => RFdata_in(11), 
                           DATAIN(10) => RFdata_in(10), DATAIN(9) => 
                           RFdata_in(9), DATAIN(8) => RFdata_in(8), DATAIN(7) 
                           => RFdata_in(7), DATAIN(6) => RFdata_in(6), 
                           DATAIN(5) => RFdata_in(5), DATAIN(4) => RFdata_in(4)
                           , DATAIN(3) => RFdata_in(3), DATAIN(2) => 
                           RFdata_in(2), DATAIN(1) => RFdata_in(1), DATAIN(0) 
                           => RFdata_in(0), OUT1(31) => RA_31_port, OUT1(30) =>
                           RA_30_port, OUT1(29) => RA_29_port, OUT1(28) => 
                           RA_28_port, OUT1(27) => RA_27_port, OUT1(26) => 
                           RA_26_port, OUT1(25) => RA_25_port, OUT1(24) => 
                           RA_24_port, OUT1(23) => RA_23_port, OUT1(22) => 
                           RA_22_port, OUT1(21) => RA_21_port, OUT1(20) => 
                           RA_20_port, OUT1(19) => RA_19_port, OUT1(18) => 
                           RA_18_port, OUT1(17) => RA_17_port, OUT1(16) => 
                           RA_16_port, OUT1(15) => RA_15_port, OUT1(14) => 
                           RA_14_port, OUT1(13) => RA_13_port, OUT1(12) => 
                           RA_12_port, OUT1(11) => RA_11_port, OUT1(10) => 
                           RA_10_port, OUT1(9) => RA_9_port, OUT1(8) => 
                           RA_8_port, OUT1(7) => RA_7_port, OUT1(6) => 
                           RA_6_port, OUT1(5) => RA_5_port, OUT1(4) => 
                           RA_4_port, OUT1(3) => RA_3_port, OUT1(2) => 
                           RA_2_port, OUT1(1) => RA_1_port, OUT1(0) => 
                           RA_0_port, OUT2(31) => RB(31), OUT2(30) => RB(30), 
                           OUT2(29) => RB(29), OUT2(28) => RB(28), OUT2(27) => 
                           RB(27), OUT2(26) => RB(26), OUT2(25) => RB(25), 
                           OUT2(24) => RB(24), OUT2(23) => RB(23), OUT2(22) => 
                           RB(22), OUT2(21) => RB(21), OUT2(20) => RB(20), 
                           OUT2(19) => RB(19), OUT2(18) => RB(18), OUT2(17) => 
                           RB(17), OUT2(16) => RB(16), OUT2(15) => RB(15), 
                           OUT2(14) => RB(14), OUT2(13) => RB(13), OUT2(12) => 
                           RB(12), OUT2(11) => RB(11), OUT2(10) => RB(10), 
                           OUT2(9) => RB(9), OUT2(8) => RB(8), OUT2(7) => RB(7)
                           , OUT2(6) => RB(6), OUT2(5) => RB(5), OUT2(4) => 
                           RB(4), OUT2(3) => RB(3), OUT2(2) => RB(2), OUT2(1) 
                           => RB(1), OUT2(0) => RB(0));
   U2 : AND2_X1 port map( A1 => IMM_15_port, A2 => n3, ZN => IMM_31_port);
   U3 : NAND4_X1 port map( A1 => n4, A2 => s_opcode_3_port, A3 => n5, A4 => n6,
                           ZN => n3);
   U4 : NAND2_X1 port map( A1 => n7, A2 => n8, ZN => n5);
   U5 : INV_X1 port map( A => s_opcode_2_port, ZN => n8);
   U6 : BUF_X2 port map( A => s_IMM26_25_port, Z => n1);
   U7 : BUF_X1 port map( A => s_IMM26_25_port, Z => n2);
   U8 : XNOR2_X1 port map( A => s_opcode_4_port, B => s_opcode_5_port, ZN => n4
                           );
   U9 : OAI211_X1 port map( C1 => s_opcode_0_port, C2 => s_opcode_4_port, A => 
                           s_opcode_1_port, B => s_opcode_2_port, ZN => n6);
   U10 : OAI22_X1 port map( A1 => s_opcode_0_port, A2 => s_opcode_4_port, B1 =>
                           s_opcode_1_port, B2 => n9, ZN => n7);
   U11 : INV_X1 port map( A => s_opcode_4_port, ZN => n9);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity FETCH is

   port( PC, hazard_PC : in std_logic_vector (31 downto 0);  PC_sel : in 
         std_logic;  IRAM_addr, NPC : out std_logic_vector (31 downto 0));

end FETCH;

architecture SYN_Behavioral of FETCH is

   component FETCH_DW01_add_0
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   component MUX21_GENERIC_NBIT32_4
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   signal IRAM_addr_31_port, IRAM_addr_30_port, IRAM_addr_29_port, 
      IRAM_addr_28_port, IRAM_addr_27_port, IRAM_addr_26_port, 
      IRAM_addr_25_port, IRAM_addr_24_port, IRAM_addr_23_port, 
      IRAM_addr_22_port, IRAM_addr_21_port, IRAM_addr_20_port, 
      IRAM_addr_19_port, IRAM_addr_18_port, IRAM_addr_17_port, 
      IRAM_addr_16_port, IRAM_addr_15_port, IRAM_addr_14_port, 
      IRAM_addr_13_port, IRAM_addr_12_port, IRAM_addr_11_port, 
      IRAM_addr_10_port, IRAM_addr_9_port, IRAM_addr_8_port, IRAM_addr_7_port, 
      IRAM_addr_6_port, IRAM_addr_5_port, IRAM_addr_4_port, IRAM_addr_3_port, 
      IRAM_addr_2_port, IRAM_addr_1_port, IRAM_addr_0_port, n1, n2, n3, n_1977 
      : std_logic;

begin
   IRAM_addr <= ( IRAM_addr_31_port, IRAM_addr_30_port, IRAM_addr_29_port, 
      IRAM_addr_28_port, IRAM_addr_27_port, IRAM_addr_26_port, 
      IRAM_addr_25_port, IRAM_addr_24_port, IRAM_addr_23_port, 
      IRAM_addr_22_port, IRAM_addr_21_port, IRAM_addr_20_port, 
      IRAM_addr_19_port, IRAM_addr_18_port, IRAM_addr_17_port, 
      IRAM_addr_16_port, IRAM_addr_15_port, IRAM_addr_14_port, 
      IRAM_addr_13_port, IRAM_addr_12_port, IRAM_addr_11_port, 
      IRAM_addr_10_port, IRAM_addr_9_port, IRAM_addr_8_port, IRAM_addr_7_port, 
      IRAM_addr_6_port, IRAM_addr_5_port, IRAM_addr_4_port, IRAM_addr_3_port, 
      IRAM_addr_2_port, IRAM_addr_1_port, IRAM_addr_0_port );
   
   n1 <= '0';
   n2 <= '1';
   n3 <= '0';
   MUX : MUX21_GENERIC_NBIT32_4 port map( A(31) => PC(31), A(30) => PC(30), 
                           A(29) => PC(29), A(28) => PC(28), A(27) => PC(27), 
                           A(26) => PC(26), A(25) => PC(25), A(24) => PC(24), 
                           A(23) => PC(23), A(22) => PC(22), A(21) => PC(21), 
                           A(20) => PC(20), A(19) => PC(19), A(18) => PC(18), 
                           A(17) => PC(17), A(16) => PC(16), A(15) => PC(15), 
                           A(14) => PC(14), A(13) => PC(13), A(12) => PC(12), 
                           A(11) => PC(11), A(10) => PC(10), A(9) => PC(9), 
                           A(8) => PC(8), A(7) => PC(7), A(6) => PC(6), A(5) =>
                           PC(5), A(4) => PC(4), A(3) => PC(3), A(2) => PC(2), 
                           A(1) => PC(1), A(0) => PC(0), B(31) => hazard_PC(31)
                           , B(30) => hazard_PC(30), B(29) => hazard_PC(29), 
                           B(28) => hazard_PC(28), B(27) => hazard_PC(27), 
                           B(26) => hazard_PC(26), B(25) => hazard_PC(25), 
                           B(24) => hazard_PC(24), B(23) => hazard_PC(23), 
                           B(22) => hazard_PC(22), B(21) => hazard_PC(21), 
                           B(20) => hazard_PC(20), B(19) => hazard_PC(19), 
                           B(18) => hazard_PC(18), B(17) => hazard_PC(17), 
                           B(16) => hazard_PC(16), B(15) => hazard_PC(15), 
                           B(14) => hazard_PC(14), B(13) => hazard_PC(13), 
                           B(12) => hazard_PC(12), B(11) => hazard_PC(11), 
                           B(10) => hazard_PC(10), B(9) => hazard_PC(9), B(8) 
                           => hazard_PC(8), B(7) => hazard_PC(7), B(6) => 
                           hazard_PC(6), B(5) => hazard_PC(5), B(4) => 
                           hazard_PC(4), B(3) => hazard_PC(3), B(2) => 
                           hazard_PC(2), B(1) => hazard_PC(1), B(0) => 
                           hazard_PC(0), SEL => PC_sel, Y(31) => 
                           IRAM_addr_31_port, Y(30) => IRAM_addr_30_port, Y(29)
                           => IRAM_addr_29_port, Y(28) => IRAM_addr_28_port, 
                           Y(27) => IRAM_addr_27_port, Y(26) => 
                           IRAM_addr_26_port, Y(25) => IRAM_addr_25_port, Y(24)
                           => IRAM_addr_24_port, Y(23) => IRAM_addr_23_port, 
                           Y(22) => IRAM_addr_22_port, Y(21) => 
                           IRAM_addr_21_port, Y(20) => IRAM_addr_20_port, Y(19)
                           => IRAM_addr_19_port, Y(18) => IRAM_addr_18_port, 
                           Y(17) => IRAM_addr_17_port, Y(16) => 
                           IRAM_addr_16_port, Y(15) => IRAM_addr_15_port, Y(14)
                           => IRAM_addr_14_port, Y(13) => IRAM_addr_13_port, 
                           Y(12) => IRAM_addr_12_port, Y(11) => 
                           IRAM_addr_11_port, Y(10) => IRAM_addr_10_port, Y(9) 
                           => IRAM_addr_9_port, Y(8) => IRAM_addr_8_port, Y(7) 
                           => IRAM_addr_7_port, Y(6) => IRAM_addr_6_port, Y(5) 
                           => IRAM_addr_5_port, Y(4) => IRAM_addr_4_port, Y(3) 
                           => IRAM_addr_3_port, Y(2) => IRAM_addr_2_port, Y(1) 
                           => IRAM_addr_1_port, Y(0) => IRAM_addr_0_port);
   add_37 : FETCH_DW01_add_0 port map( A(31) => IRAM_addr_31_port, A(30) => 
                           IRAM_addr_30_port, A(29) => IRAM_addr_29_port, A(28)
                           => IRAM_addr_28_port, A(27) => IRAM_addr_27_port, 
                           A(26) => IRAM_addr_26_port, A(25) => 
                           IRAM_addr_25_port, A(24) => IRAM_addr_24_port, A(23)
                           => IRAM_addr_23_port, A(22) => IRAM_addr_22_port, 
                           A(21) => IRAM_addr_21_port, A(20) => 
                           IRAM_addr_20_port, A(19) => IRAM_addr_19_port, A(18)
                           => IRAM_addr_18_port, A(17) => IRAM_addr_17_port, 
                           A(16) => IRAM_addr_16_port, A(15) => 
                           IRAM_addr_15_port, A(14) => IRAM_addr_14_port, A(13)
                           => IRAM_addr_13_port, A(12) => IRAM_addr_12_port, 
                           A(11) => IRAM_addr_11_port, A(10) => 
                           IRAM_addr_10_port, A(9) => IRAM_addr_9_port, A(8) =>
                           IRAM_addr_8_port, A(7) => IRAM_addr_7_port, A(6) => 
                           IRAM_addr_6_port, A(5) => IRAM_addr_5_port, A(4) => 
                           IRAM_addr_4_port, A(3) => IRAM_addr_3_port, A(2) => 
                           IRAM_addr_2_port, A(1) => IRAM_addr_1_port, A(0) => 
                           IRAM_addr_0_port, B(31) => n3, B(30) => n3, B(29) =>
                           n3, B(28) => n3, B(27) => n3, B(26) => n3, B(25) => 
                           n3, B(24) => n3, B(23) => n3, B(22) => n3, B(21) => 
                           n3, B(20) => n3, B(19) => n3, B(18) => n3, B(17) => 
                           n3, B(16) => n3, B(15) => n3, B(14) => n3, B(13) => 
                           n3, B(12) => n3, B(11) => n3, B(10) => n3, B(9) => 
                           n3, B(8) => n3, B(7) => n3, B(6) => n3, B(5) => n3, 
                           B(4) => n3, B(3) => n3, B(2) => n2, B(1) => n1, B(0)
                           => n1, CI => n3, SUM(31) => NPC(31), SUM(30) => 
                           NPC(30), SUM(29) => NPC(29), SUM(28) => NPC(28), 
                           SUM(27) => NPC(27), SUM(26) => NPC(26), SUM(25) => 
                           NPC(25), SUM(24) => NPC(24), SUM(23) => NPC(23), 
                           SUM(22) => NPC(22), SUM(21) => NPC(21), SUM(20) => 
                           NPC(20), SUM(19) => NPC(19), SUM(18) => NPC(18), 
                           SUM(17) => NPC(17), SUM(16) => NPC(16), SUM(15) => 
                           NPC(15), SUM(14) => NPC(14), SUM(13) => NPC(13), 
                           SUM(12) => NPC(12), SUM(11) => NPC(11), SUM(10) => 
                           NPC(10), SUM(9) => NPC(9), SUM(8) => NPC(8), SUM(7) 
                           => NPC(7), SUM(6) => NPC(6), SUM(5) => NPC(5), 
                           SUM(4) => NPC(4), SUM(3) => NPC(3), SUM(2) => NPC(2)
                           , SUM(1) => NPC(1), SUM(0) => NPC(0), CO => n_1977);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity MUX21_GENERIC_NBIT32_0 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end MUX21_GENERIC_NBIT32_0;

architecture SYN_structural of MUX21_GENERIC_NBIT32_0 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX21_563
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_564
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_565
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_566
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_567
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_568
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_569
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_570
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_571
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_572
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_573
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_574
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_575
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_576
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_577
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_578
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_579
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_580
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_581
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_582
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_583
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_584
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_585
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_586
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_587
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_588
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_589
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_590
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_591
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_592
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_593
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   component MUX21_0
      port( A, B, S : in std_logic;  Y : out std_logic);
   end component;
   
   signal n1, n2, n3 : std_logic;

begin
   
   MUXES_0 : MUX21_0 port map( A => A(0), B => B(0), S => n3, Y => Y(0));
   MUXES_1 : MUX21_593 port map( A => A(1), B => B(1), S => n1, Y => Y(1));
   MUXES_2 : MUX21_592 port map( A => A(2), B => B(2), S => n1, Y => Y(2));
   MUXES_3 : MUX21_591 port map( A => A(3), B => B(3), S => n1, Y => Y(3));
   MUXES_4 : MUX21_590 port map( A => A(4), B => B(4), S => n1, Y => Y(4));
   MUXES_5 : MUX21_589 port map( A => A(5), B => B(5), S => n1, Y => Y(5));
   MUXES_6 : MUX21_588 port map( A => A(6), B => B(6), S => n1, Y => Y(6));
   MUXES_7 : MUX21_587 port map( A => A(7), B => B(7), S => n1, Y => Y(7));
   MUXES_8 : MUX21_586 port map( A => A(8), B => B(8), S => n1, Y => Y(8));
   MUXES_9 : MUX21_585 port map( A => A(9), B => B(9), S => n1, Y => Y(9));
   MUXES_10 : MUX21_584 port map( A => A(10), B => B(10), S => n1, Y => Y(10));
   MUXES_11 : MUX21_583 port map( A => A(11), B => B(11), S => n1, Y => Y(11));
   MUXES_12 : MUX21_582 port map( A => A(12), B => B(12), S => n1, Y => Y(12));
   MUXES_13 : MUX21_581 port map( A => A(13), B => B(13), S => n2, Y => Y(13));
   MUXES_14 : MUX21_580 port map( A => A(14), B => B(14), S => n2, Y => Y(14));
   MUXES_15 : MUX21_579 port map( A => A(15), B => B(15), S => n2, Y => Y(15));
   MUXES_16 : MUX21_578 port map( A => A(16), B => B(16), S => n2, Y => Y(16));
   MUXES_17 : MUX21_577 port map( A => A(17), B => B(17), S => n2, Y => Y(17));
   MUXES_18 : MUX21_576 port map( A => A(18), B => B(18), S => n2, Y => Y(18));
   MUXES_19 : MUX21_575 port map( A => A(19), B => B(19), S => n2, Y => Y(19));
   MUXES_20 : MUX21_574 port map( A => A(20), B => B(20), S => n2, Y => Y(20));
   MUXES_21 : MUX21_573 port map( A => A(21), B => B(21), S => n2, Y => Y(21));
   MUXES_22 : MUX21_572 port map( A => A(22), B => B(22), S => n2, Y => Y(22));
   MUXES_23 : MUX21_571 port map( A => A(23), B => B(23), S => n2, Y => Y(23));
   MUXES_24 : MUX21_570 port map( A => A(24), B => B(24), S => n2, Y => Y(24));
   MUXES_25 : MUX21_569 port map( A => A(25), B => B(25), S => n3, Y => Y(25));
   MUXES_26 : MUX21_568 port map( A => A(26), B => B(26), S => n3, Y => Y(26));
   MUXES_27 : MUX21_567 port map( A => A(27), B => B(27), S => n3, Y => Y(27));
   MUXES_28 : MUX21_566 port map( A => A(28), B => B(28), S => n3, Y => Y(28));
   MUXES_29 : MUX21_565 port map( A => A(29), B => B(29), S => n3, Y => Y(29));
   MUXES_30 : MUX21_564 port map( A => A(30), B => B(30), S => n3, Y => Y(30));
   MUXES_31 : MUX21_563 port map( A => A(31), B => B(31), S => n3, Y => Y(31));
   U1 : BUF_X1 port map( A => SEL, Z => n2);
   U2 : BUF_X1 port map( A => SEL, Z => n1);
   U3 : BUF_X1 port map( A => SEL, Z => n3);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity DataPath_MEM_SIZE128_WORD_size32_NREG32 is

   port( CLK, RST, RF1, RF2, EN1, S1, S2, ALU3, ALU2, ALU1, ALU0, SN, LnS, BHU1
         , BHU0, Wrd, EN3, S3, WF1, Ld : in std_logic;  instr : in 
         std_logic_vector (31 downto 0);  IRAM_addr : out std_logic_vector (31 
         downto 0);  DRAM_data_out : in std_logic_vector (31 downto 0);  
         MMU_out : out std_logic_vector (1 downto 0);  DRAM_addr : out 
         std_logic_vector (8 downto 0);  DRAM_data_in : out std_logic_vector 
         (31 downto 0);  opcode : out std_logic_vector (5 downto 0);  func : 
         out std_logic_vector (10 downto 0);  OVF : out std_logic);

end DataPath_MEM_SIZE128_WORD_size32_NREG32;

architecture SYN_Structural of DataPath_MEM_SIZE128_WORD_size32_NREG32 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFS_X1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFS_X2
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component WB
      port( mem_out, alu_out : in std_logic_vector (31 downto 0);  S3 : in 
            std_logic;  output : out std_logic_vector (31 downto 0));
   end component;
   
   component MEM_MEMORY_SIZE128
      port( CLK, RST : in std_logic;  ALUout, MEout : in std_logic_vector (31 
            downto 0);  RDin : in std_logic_vector (4 downto 0);  DRAM_data_out
            : in std_logic_vector (31 downto 0);  LnS, Wrd, BHU1, BHU0, EN3 : 
            in std_logic;  DRAM_addr : out std_logic_vector (8 downto 0);  
            DRAM_data_in : out std_logic_vector (31 downto 0);  MMU_out : out 
            std_logic_vector (1 downto 0);  output, alu_out : out 
            std_logic_vector (31 downto 0);  RDout : out std_logic_vector (4 
            downto 0));
   end component;
   
   component EXE
      port( CLK, RST : in std_logic;  IMM, RA, RB : in std_logic_vector (31 
            downto 0);  WA, RSA, RSB : in std_logic_vector (4 downto 0);  
            ALU_outmem, WB_out : in std_logic_vector (31 downto 0);  MEM_RD, 
            WB_RD : in std_logic_vector (4 downto 0);  LD_EN, WB_EN, S1, S2, 
            ALU3, ALU2, ALU1, ALU0, SN : in std_logic;  RD_inmul : out 
            std_logic_vector (4 downto 0);  flag_structHzd, flag_ismul, OVF : 
            out std_logic;  output, ME : out std_logic_vector (31 downto 0);  
            WAout : out std_logic_vector (4 downto 0));
   end component;
   
   component DEC
      port( instr : in std_logic_vector (31 downto 0);  RST : in std_logic;  
            RFdata_in : in std_logic_vector (31 downto 0);  RFWA : in 
            std_logic_vector (4 downto 0);  NPC_in : in std_logic_vector (31 
            downto 0);  EXE_RD : in std_logic_vector (4 downto 0);  Ld : in 
            std_logic;  ALU_regout : in std_logic_vector (31 downto 0);  MEM_RD
            , WB_RD, RD_inmul : in std_logic_vector (4 downto 0);  
            flag_structHzd, flag_ismul, RF1, RF2, WF1, EN1 : in std_logic;  
            opcode : out std_logic_vector (5 downto 0);  func : out 
            std_logic_vector (10 downto 0);  IMM, RA, RB : out std_logic_vector
            (31 downto 0);  RSA, RSB, RD : out std_logic_vector (4 downto 0);  
            stall_NPC : out std_logic_vector (31 downto 0);  PC_sel, dec_flag :
            out std_logic;  NPC_jump : out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT32_5
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component FETCH
      port( PC, hazard_PC : in std_logic_vector (31 downto 0);  PC_sel : in 
            std_logic;  IRAM_addr, NPC : out std_logic_vector (31 downto 0));
   end component;
   
   component MUX21_GENERIC_NBIT32_0
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, PC_reg_31_port, PC_reg_30_port, 
      PC_reg_29_port, PC_reg_28_port, PC_reg_27_port, PC_reg_26_port, 
      PC_reg_25_port, PC_reg_24_port, PC_reg_23_port, PC_reg_22_port, 
      PC_reg_21_port, PC_reg_20_port, PC_reg_19_port, PC_reg_18_port, 
      PC_reg_17_port, PC_reg_16_port, PC_reg_15_port, PC_reg_14_port, 
      PC_reg_13_port, PC_reg_12_port, PC_reg_11_port, PC_reg_10_port, 
      PC_reg_9_port, PC_reg_8_port, PC_reg_7_port, PC_reg_6_port, PC_reg_5_port
      , PC_reg_4_port, PC_reg_3_port, PC_reg_2_port, PC_reg_1_port, 
      PC_reg_0_port, NPC_reg_31_port, NPC_reg_30_port, NPC_reg_29_port, 
      NPC_reg_28_port, NPC_reg_27_port, NPC_reg_26_port, NPC_reg_25_port, 
      NPC_reg_24_port, NPC_reg_23_port, NPC_reg_22_port, NPC_reg_21_port, 
      NPC_reg_20_port, NPC_reg_19_port, NPC_reg_18_port, NPC_reg_17_port, 
      NPC_reg_16_port, NPC_reg_15_port, NPC_reg_14_port, NPC_reg_13_port, 
      NPC_reg_12_port, NPC_reg_11_port, NPC_reg_10_port, NPC_reg_9_port, 
      NPC_reg_8_port, NPC_reg_7_port, NPC_reg_6_port, NPC_reg_5_port, 
      NPC_reg_4_port, NPC_reg_3_port, NPC_reg_2_port, NPC_reg_1_port, 
      NPC_reg_0_port, IR_reg_31_port, IR_reg_30_port, IR_reg_29_port, 
      IR_reg_28_port, IR_reg_27_port, IR_reg_26_port, IR_reg_25_port, 
      IR_reg_24_port, IR_reg_23_port, IR_reg_22_port, IR_reg_21_port, 
      IR_reg_20_port, IR_reg_19_port, IR_reg_18_port, IR_reg_17_port, 
      IR_reg_16_port, IR_reg_15_port, IR_reg_14_port, IR_reg_13_port, 
      IR_reg_12_port, IR_reg_11_port, IR_reg_10_port, IR_reg_9_port, 
      IR_reg_8_port, IR_reg_7_port, IR_reg_6_port, IR_reg_5_port, IR_reg_4_port
      , IR_reg_3_port, IR_reg_2_port, IR_reg_1_port, IR_reg_0_port, 
      Imm_reg_31_port, Imm_reg_30_port, Imm_reg_29_port, Imm_reg_28_port, 
      Imm_reg_27_port, Imm_reg_26_port, Imm_reg_25_port, Imm_reg_24_port, 
      Imm_reg_23_port, Imm_reg_22_port, Imm_reg_21_port, Imm_reg_20_port, 
      Imm_reg_19_port, Imm_reg_18_port, Imm_reg_17_port, Imm_reg_16_port, 
      Imm_reg_15_port, Imm_reg_14_port, Imm_reg_13_port, Imm_reg_12_port, 
      Imm_reg_11_port, Imm_reg_10_port, Imm_reg_9_port, Imm_reg_8_port, 
      Imm_reg_7_port, Imm_reg_6_port, Imm_reg_5_port, Imm_reg_4_port, 
      Imm_reg_3_port, Imm_reg_2_port, Imm_reg_1_port, Imm_reg_0_port, 
      RA_reg_31_port, RA_reg_30_port, RA_reg_29_port, RA_reg_28_port, 
      RA_reg_27_port, RA_reg_26_port, RA_reg_25_port, RA_reg_24_port, 
      RA_reg_23_port, RA_reg_22_port, RA_reg_21_port, RA_reg_20_port, 
      RA_reg_19_port, RA_reg_18_port, RA_reg_17_port, RA_reg_16_port, 
      RA_reg_15_port, RA_reg_14_port, RA_reg_13_port, RA_reg_12_port, 
      RA_reg_11_port, RA_reg_10_port, RA_reg_9_port, RA_reg_8_port, 
      RA_reg_7_port, RA_reg_6_port, RA_reg_5_port, RA_reg_4_port, RA_reg_3_port
      , RA_reg_2_port, RA_reg_1_port, RA_reg_0_port, RB_reg_31_port, 
      RB_reg_30_port, RB_reg_29_port, RB_reg_28_port, RB_reg_27_port, 
      RB_reg_26_port, RB_reg_25_port, RB_reg_24_port, RB_reg_23_port, 
      RB_reg_22_port, RB_reg_21_port, RB_reg_20_port, RB_reg_19_port, 
      RB_reg_18_port, RB_reg_17_port, RB_reg_16_port, RB_reg_15_port, 
      RB_reg_14_port, RB_reg_13_port, RB_reg_12_port, RB_reg_11_port, 
      RB_reg_10_port, RB_reg_9_port, RB_reg_8_port, RB_reg_7_port, 
      RB_reg_6_port, RB_reg_5_port, RB_reg_4_port, RB_reg_3_port, RB_reg_2_port
      , RB_reg_1_port, RB_reg_0_port, RSA_reg_4_port, RSA_reg_3_port, 
      RSA_reg_2_port, RSA_reg_1_port, RSA_reg_0_port, RSB_reg_4_port, 
      RSB_reg_3_port, RSB_reg_2_port, RSB_reg_1_port, RSB_reg_0_port, 
      RD_regexe_4_port, RD_regexe_3_port, RD_regexe_2_port, RD_regexe_1_port, 
      RD_regexe_0_port, ALU_reg_31_port, ALU_reg_30_port, ALU_reg_29_port, 
      ALU_reg_28_port, ALU_reg_27_port, ALU_reg_26_port, ALU_reg_25_port, 
      ALU_reg_24_port, ALU_reg_23_port, ALU_reg_22_port, ALU_reg_21_port, 
      ALU_reg_20_port, ALU_reg_19_port, ALU_reg_18_port, ALU_reg_17_port, 
      ALU_reg_16_port, ALU_reg_15_port, ALU_reg_14_port, ALU_reg_13_port, 
      ALU_reg_12_port, ALU_reg_11_port, ALU_reg_10_port, ALU_reg_9_port, 
      ALU_reg_8_port, ALU_reg_7_port, ALU_reg_6_port, ALU_reg_5_port, 
      ALU_reg_4_port, ALU_reg_3_port, ALU_reg_2_port, ALU_reg_1_port, 
      ALU_reg_0_port, ME_reg_31_port, ME_reg_30_port, ME_reg_29_port, 
      ME_reg_28_port, ME_reg_27_port, ME_reg_26_port, ME_reg_25_port, 
      ME_reg_24_port, ME_reg_23_port, ME_reg_22_port, ME_reg_21_port, 
      ME_reg_20_port, ME_reg_19_port, ME_reg_18_port, ME_reg_17_port, 
      ME_reg_16_port, ME_reg_15_port, ME_reg_14_port, ME_reg_13_port, 
      ME_reg_12_port, ME_reg_11_port, ME_reg_10_port, ME_reg_9_port, 
      ME_reg_8_port, ME_reg_7_port, ME_reg_6_port, ME_reg_5_port, ME_reg_4_port
      , ME_reg_3_port, ME_reg_2_port, ME_reg_1_port, ME_reg_0_port, 
      RD_regmem_4_port, RD_regmem_3_port, RD_regmem_2_port, RD_regmem_1_port, 
      RD_regmem_0_port, LMD_reg_31_port, LMD_reg_30_port, LMD_reg_29_port, 
      LMD_reg_28_port, LMD_reg_27_port, LMD_reg_26_port, LMD_reg_25_port, 
      LMD_reg_24_port, LMD_reg_23_port, LMD_reg_22_port, LMD_reg_21_port, 
      LMD_reg_20_port, LMD_reg_19_port, LMD_reg_18_port, LMD_reg_17_port, 
      LMD_reg_16_port, LMD_reg_15_port, LMD_reg_14_port, LMD_reg_13_port, 
      LMD_reg_12_port, LMD_reg_11_port, LMD_reg_10_port, LMD_reg_9_port, 
      LMD_reg_8_port, LMD_reg_7_port, LMD_reg_6_port, LMD_reg_5_port, 
      LMD_reg_4_port, LMD_reg_3_port, LMD_reg_2_port, LMD_reg_1_port, 
      LMD_reg_0_port, ALU_regmem_31_port, ALU_regmem_30_port, 
      ALU_regmem_29_port, ALU_regmem_28_port, ALU_regmem_27_port, 
      ALU_regmem_26_port, ALU_regmem_25_port, ALU_regmem_24_port, 
      ALU_regmem_23_port, ALU_regmem_22_port, ALU_regmem_21_port, 
      ALU_regmem_20_port, ALU_regmem_19_port, ALU_regmem_18_port, 
      ALU_regmem_17_port, ALU_regmem_16_port, ALU_regmem_15_port, 
      ALU_regmem_14_port, ALU_regmem_13_port, ALU_regmem_12_port, 
      ALU_regmem_11_port, ALU_regmem_10_port, ALU_regmem_9_port, 
      ALU_regmem_8_port, ALU_regmem_7_port, ALU_regmem_6_port, 
      ALU_regmem_5_port, ALU_regmem_4_port, ALU_regmem_3_port, 
      ALU_regmem_2_port, ALU_regmem_1_port, ALU_regmem_0_port, RD_regwb_4_port,
      RD_regwb_3_port, RD_regwb_2_port, RD_regwb_1_port, RD_regwb_0_port, 
      PC_muxout_31_port, PC_muxout_30_port, PC_muxout_29_port, 
      PC_muxout_28_port, PC_muxout_27_port, PC_muxout_26_port, 
      PC_muxout_25_port, PC_muxout_24_port, PC_muxout_23_port, 
      PC_muxout_22_port, PC_muxout_21_port, PC_muxout_20_port, 
      PC_muxout_19_port, PC_muxout_18_port, PC_muxout_17_port, 
      PC_muxout_16_port, PC_muxout_15_port, PC_muxout_14_port, 
      PC_muxout_13_port, PC_muxout_12_port, PC_muxout_11_port, 
      PC_muxout_10_port, PC_muxout_9_port, PC_muxout_8_port, PC_muxout_7_port, 
      PC_muxout_6_port, PC_muxout_5_port, PC_muxout_4_port, PC_muxout_3_port, 
      PC_muxout_2_port, PC_muxout_1_port, PC_muxout_0_port, 
      NPC_fetchout_31_port, NPC_fetchout_30_port, NPC_fetchout_29_port, 
      NPC_fetchout_28_port, NPC_fetchout_27_port, NPC_fetchout_26_port, 
      NPC_fetchout_25_port, NPC_fetchout_24_port, NPC_fetchout_23_port, 
      NPC_fetchout_22_port, NPC_fetchout_21_port, NPC_fetchout_20_port, 
      NPC_fetchout_19_port, NPC_fetchout_18_port, NPC_fetchout_17_port, 
      NPC_fetchout_16_port, NPC_fetchout_15_port, NPC_fetchout_14_port, 
      NPC_fetchout_13_port, NPC_fetchout_12_port, NPC_fetchout_11_port, 
      NPC_fetchout_10_port, NPC_fetchout_9_port, NPC_fetchout_8_port, 
      NPC_fetchout_7_port, NPC_fetchout_6_port, NPC_fetchout_5_port, 
      NPC_fetchout_4_port, NPC_fetchout_3_port, NPC_fetchout_2_port, 
      NPC_fetchout_1_port, NPC_fetchout_0_port, NOP_MUX_OUT_31_port, 
      NOP_MUX_OUT_30_port, NOP_MUX_OUT_29_port, NOP_MUX_OUT_28_port, 
      NOP_MUX_OUT_27_port, NOP_MUX_OUT_26_port, NOP_MUX_OUT_25_port, 
      NOP_MUX_OUT_24_port, NOP_MUX_OUT_23_port, NOP_MUX_OUT_22_port, 
      NOP_MUX_OUT_21_port, NOP_MUX_OUT_20_port, NOP_MUX_OUT_19_port, 
      NOP_MUX_OUT_18_port, NOP_MUX_OUT_17_port, NOP_MUX_OUT_16_port, 
      NOP_MUX_OUT_15_port, NOP_MUX_OUT_14_port, NOP_MUX_OUT_13_port, 
      NOP_MUX_OUT_12_port, NOP_MUX_OUT_11_port, NOP_MUX_OUT_10_port, 
      NOP_MUX_OUT_9_port, NOP_MUX_OUT_8_port, NOP_MUX_OUT_7_port, 
      NOP_MUX_OUT_6_port, NOP_MUX_OUT_5_port, NOP_MUX_OUT_4_port, 
      NOP_MUX_OUT_3_port, NOP_MUX_OUT_2_port, NOP_MUX_OUT_1_port, 
      NOP_MUX_OUT_0_port, IMM_decout_31_port, IMM_decout_30_port, 
      IMM_decout_29_port, IMM_decout_28_port, IMM_decout_27_port, 
      IMM_decout_26_port, IMM_decout_25_port, IMM_decout_24_port, 
      IMM_decout_23_port, IMM_decout_22_port, IMM_decout_21_port, 
      IMM_decout_20_port, IMM_decout_19_port, IMM_decout_18_port, 
      IMM_decout_17_port, IMM_decout_16_port, IMM_decout_15_port, 
      IMM_decout_14_port, IMM_decout_13_port, IMM_decout_12_port, 
      IMM_decout_11_port, IMM_decout_10_port, IMM_decout_9_port, 
      IMM_decout_8_port, IMM_decout_7_port, IMM_decout_6_port, 
      IMM_decout_5_port, IMM_decout_4_port, IMM_decout_3_port, 
      IMM_decout_2_port, IMM_decout_1_port, IMM_decout_0_port, 
      RA_decout_31_port, RA_decout_30_port, RA_decout_29_port, 
      RA_decout_28_port, RA_decout_27_port, RA_decout_26_port, 
      RA_decout_25_port, RA_decout_24_port, RA_decout_23_port, 
      RA_decout_22_port, RA_decout_21_port, RA_decout_20_port, 
      RA_decout_19_port, RA_decout_18_port, RA_decout_17_port, 
      RA_decout_16_port, RA_decout_15_port, RA_decout_14_port, 
      RA_decout_13_port, RA_decout_12_port, RA_decout_11_port, 
      RA_decout_10_port, RA_decout_9_port, RA_decout_8_port, RA_decout_7_port, 
      RA_decout_6_port, RA_decout_5_port, RA_decout_4_port, RA_decout_3_port, 
      RA_decout_2_port, RA_decout_1_port, RA_decout_0_port, RB_decout_31_port, 
      RB_decout_30_port, RB_decout_29_port, RB_decout_28_port, 
      RB_decout_27_port, RB_decout_26_port, RB_decout_25_port, 
      RB_decout_24_port, RB_decout_23_port, RB_decout_22_port, 
      RB_decout_21_port, RB_decout_20_port, RB_decout_19_port, 
      RB_decout_18_port, RB_decout_17_port, RB_decout_16_port, 
      RB_decout_15_port, RB_decout_14_port, RB_decout_13_port, 
      RB_decout_12_port, RB_decout_11_port, RB_decout_10_port, RB_decout_9_port
      , RB_decout_8_port, RB_decout_7_port, RB_decout_6_port, RB_decout_5_port,
      RB_decout_4_port, RB_decout_3_port, RB_decout_2_port, RB_decout_1_port, 
      RB_decout_0_port, RD_decout_4_port, RD_decout_3_port, RD_decout_2_port, 
      RD_decout_1_port, RD_decout_0_port, RSA_decout_4_port, RSA_decout_3_port,
      RSA_decout_2_port, RSA_decout_1_port, RSA_decout_0_port, 
      RSB_decout_4_port, RSB_decout_3_port, RSB_decout_2_port, 
      RSB_decout_1_port, RSB_decout_0_port, ALU_exeout_31_port, 
      ALU_exeout_30_port, ALU_exeout_29_port, ALU_exeout_28_port, 
      ALU_exeout_27_port, ALU_exeout_26_port, ALU_exeout_25_port, 
      ALU_exeout_24_port, ALU_exeout_23_port, ALU_exeout_22_port, 
      ALU_exeout_21_port, ALU_exeout_20_port, ALU_exeout_19_port, 
      ALU_exeout_18_port, ALU_exeout_17_port, ALU_exeout_16_port, 
      ALU_exeout_15_port, ALU_exeout_14_port, ALU_exeout_13_port, 
      ALU_exeout_12_port, ALU_exeout_11_port, ALU_exeout_10_port, 
      ALU_exeout_9_port, ALU_exeout_8_port, ALU_exeout_7_port, 
      ALU_exeout_6_port, ALU_exeout_5_port, ALU_exeout_4_port, 
      ALU_exeout_3_port, ALU_exeout_2_port, ALU_exeout_1_port, 
      ALU_exeout_0_port, ME_exeout_31_port, ME_exeout_30_port, 
      ME_exeout_29_port, ME_exeout_28_port, ME_exeout_27_port, 
      ME_exeout_26_port, ME_exeout_25_port, ME_exeout_24_port, 
      ME_exeout_23_port, ME_exeout_22_port, ME_exeout_21_port, 
      ME_exeout_20_port, ME_exeout_19_port, ME_exeout_18_port, 
      ME_exeout_17_port, ME_exeout_16_port, ME_exeout_15_port, 
      ME_exeout_14_port, ME_exeout_13_port, ME_exeout_12_port, 
      ME_exeout_11_port, ME_exeout_10_port, ME_exeout_9_port, ME_exeout_8_port,
      ME_exeout_7_port, ME_exeout_6_port, ME_exeout_5_port, ME_exeout_4_port, 
      ME_exeout_3_port, ME_exeout_2_port, ME_exeout_1_port, ME_exeout_0_port, 
      RD_exeout_4_port, RD_exeout_3_port, RD_exeout_2_port, RD_exeout_1_port, 
      RD_exeout_0_port, mem_out_31_port, mem_out_30_port, mem_out_29_port, 
      mem_out_28_port, mem_out_27_port, mem_out_26_port, mem_out_25_port, 
      mem_out_24_port, mem_out_23_port, mem_out_22_port, mem_out_21_port, 
      mem_out_20_port, mem_out_19_port, mem_out_18_port, mem_out_17_port, 
      mem_out_16_port, mem_out_15_port, mem_out_14_port, mem_out_13_port, 
      mem_out_12_port, mem_out_11_port, mem_out_10_port, mem_out_9_port, 
      mem_out_8_port, mem_out_7_port, mem_out_6_port, mem_out_5_port, 
      mem_out_4_port, mem_out_3_port, mem_out_2_port, mem_out_1_port, 
      mem_out_0_port, ALU_memout_31_port, ALU_memout_30_port, 
      ALU_memout_29_port, ALU_memout_28_port, ALU_memout_27_port, 
      ALU_memout_26_port, ALU_memout_25_port, ALU_memout_24_port, 
      ALU_memout_23_port, ALU_memout_22_port, ALU_memout_21_port, 
      ALU_memout_20_port, ALU_memout_19_port, ALU_memout_18_port, 
      ALU_memout_17_port, ALU_memout_16_port, ALU_memout_15_port, 
      ALU_memout_14_port, ALU_memout_13_port, ALU_memout_12_port, 
      ALU_memout_11_port, ALU_memout_10_port, ALU_memout_9_port, 
      ALU_memout_8_port, ALU_memout_7_port, ALU_memout_6_port, 
      ALU_memout_5_port, ALU_memout_4_port, ALU_memout_3_port, 
      ALU_memout_2_port, ALU_memout_1_port, ALU_memout_0_port, RD_memout_4_port
      , RD_memout_3_port, RD_memout_2_port, RD_memout_1_port, RD_memout_0_port,
      s_NPC_jump_31_port, s_NPC_jump_30_port, s_NPC_jump_29_port, 
      s_NPC_jump_28_port, s_NPC_jump_27_port, s_NPC_jump_26_port, 
      s_NPC_jump_25_port, s_NPC_jump_24_port, s_NPC_jump_23_port, 
      s_NPC_jump_22_port, s_NPC_jump_21_port, s_NPC_jump_20_port, 
      s_NPC_jump_19_port, s_NPC_jump_18_port, s_NPC_jump_17_port, 
      s_NPC_jump_16_port, s_NPC_jump_15_port, s_NPC_jump_14_port, 
      s_NPC_jump_13_port, s_NPC_jump_12_port, s_NPC_jump_11_port, 
      s_NPC_jump_10_port, s_NPC_jump_9_port, s_NPC_jump_8_port, 
      s_NPC_jump_7_port, s_NPC_jump_6_port, s_NPC_jump_5_port, 
      s_NPC_jump_4_port, s_NPC_jump_3_port, s_NPC_jump_2_port, 
      s_NPC_jump_1_port, s_NPC_jump_0_port, flag_signal, hazard_NPC_31_port, 
      hazard_NPC_30_port, hazard_NPC_29_port, hazard_NPC_28_port, 
      hazard_NPC_27_port, hazard_NPC_26_port, hazard_NPC_25_port, 
      hazard_NPC_24_port, hazard_NPC_23_port, hazard_NPC_22_port, 
      hazard_NPC_21_port, hazard_NPC_20_port, hazard_NPC_19_port, 
      hazard_NPC_18_port, hazard_NPC_17_port, hazard_NPC_16_port, 
      hazard_NPC_15_port, hazard_NPC_14_port, hazard_NPC_13_port, 
      hazard_NPC_12_port, hazard_NPC_11_port, hazard_NPC_10_port, 
      hazard_NPC_9_port, hazard_NPC_8_port, hazard_NPC_7_port, 
      hazard_NPC_6_port, hazard_NPC_5_port, hazard_NPC_4_port, 
      hazard_NPC_3_port, hazard_NPC_2_port, hazard_NPC_1_port, 
      hazard_NPC_0_port, hazard_NPC_sel, WB_data_31_port, WB_data_30_port, 
      WB_data_29_port, WB_data_28_port, WB_data_27_port, WB_data_26_port, 
      WB_data_25_port, WB_data_24_port, WB_data_23_port, WB_data_22_port, 
      WB_data_21_port, WB_data_20_port, WB_data_19_port, WB_data_18_port, 
      WB_data_17_port, WB_data_16_port, WB_data_15_port, WB_data_14_port, 
      WB_data_13_port, WB_data_12_port, WB_data_11_port, WB_data_10_port, 
      WB_data_9_port, WB_data_8_port, WB_data_7_port, WB_data_6_port, 
      WB_data_5_port, WB_data_4_port, WB_data_3_port, WB_data_2_port, 
      WB_data_1_port, WB_data_0_port, s_RD_inmul_4_port, s_RD_inmul_3_port, 
      s_RD_inmul_2_port, s_RD_inmul_1_port, s_RD_inmul_0_port, s_flag_structHzd
      , s_flag_ismul, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n_1978
      , n_1979, n_1980, n_1981, n_1982, n_1983, n_1984, n_1985, n_1986, n_1987,
      n_1988, n_1989, n_1990, n_1991, n_1992, n_1993, n_1994, n_1995, n_1996, 
      n_1997, n_1998, n_1999, n_2000, n_2001, n_2002, n_2003, n_2004, n_2005, 
      n_2006, n_2007, n_2008, n_2009, n_2010, n_2011, n_2012, n_2013, n_2014, 
      n_2015, n_2016, n_2017, n_2018, n_2019, n_2020, n_2021, n_2022, n_2023, 
      n_2024, n_2025, n_2026, n_2027, n_2028, n_2029, n_2030, n_2031, n_2032, 
      n_2033, n_2034, n_2035, n_2036, n_2037, n_2038, n_2039, n_2040, n_2041, 
      n_2042, n_2043, n_2044, n_2045, n_2046, n_2047, n_2048, n_2049, n_2050, 
      n_2051, n_2052, n_2053, n_2054, n_2055, n_2056, n_2057, n_2058, n_2059, 
      n_2060, n_2061, n_2062, n_2063, n_2064, n_2065, n_2066, n_2067, n_2068, 
      n_2069, n_2070, n_2071, n_2072, n_2073, n_2074, n_2075, n_2076, n_2077, 
      n_2078, n_2079, n_2080, n_2081, n_2082, n_2083, n_2084, n_2085, n_2086, 
      n_2087, n_2088, n_2089, n_2090, n_2091, n_2092, n_2093, n_2094, n_2095, 
      n_2096, n_2097, n_2098, n_2099, n_2100, n_2101, n_2102, n_2103, n_2104, 
      n_2105, n_2106, n_2107, n_2108, n_2109, n_2110, n_2111, n_2112, n_2113, 
      n_2114, n_2115, n_2116, n_2117, n_2118, n_2119, n_2120, n_2121, n_2122, 
      n_2123, n_2124, n_2125, n_2126, n_2127, n_2128, n_2129, n_2130, n_2131, 
      n_2132, n_2133, n_2134, n_2135, n_2136, n_2137, n_2138, n_2139, n_2140, 
      n_2141, n_2142, n_2143, n_2144, n_2145, n_2146, n_2147, n_2148, n_2149, 
      n_2150, n_2151, n_2152, n_2153, n_2154, n_2155, n_2156, n_2157, n_2158, 
      n_2159, n_2160, n_2161, n_2162, n_2163, n_2164, n_2165, n_2166, n_2167, 
      n_2168, n_2169, n_2170, n_2171, n_2172, n_2173, n_2174, n_2175, n_2176, 
      n_2177, n_2178, n_2179, n_2180, n_2181, n_2182, n_2183, n_2184, n_2185, 
      n_2186, n_2187, n_2188, n_2189, n_2190, n_2191, n_2192, n_2193, n_2194, 
      n_2195, n_2196, n_2197, n_2198, n_2199, n_2200, n_2201, n_2202, n_2203, 
      n_2204, n_2205, n_2206, n_2207, n_2208, n_2209, n_2210, n_2211, n_2212, 
      n_2213, n_2214, n_2215, n_2216, n_2217, n_2218, n_2219, n_2220, n_2221, 
      n_2222, n_2223, n_2224, n_2225, n_2226, n_2227, n_2228, n_2229, n_2230, 
      n_2231, n_2232, n_2233, n_2234, n_2235, n_2236, n_2237, n_2238, n_2239, 
      n_2240, n_2241, n_2242, n_2243, n_2244, n_2245, n_2246, n_2247, n_2248, 
      n_2249, n_2250, n_2251, n_2252, n_2253, n_2254, n_2255, n_2256, n_2257, 
      n_2258, n_2259, n_2260, n_2261, n_2262, n_2263, n_2264, n_2265, n_2266, 
      n_2267, n_2268, n_2269, n_2270, n_2271, n_2272, n_2273, n_2274, n_2275, 
      n_2276, n_2277, n_2278, n_2279, n_2280, n_2281, n_2282, n_2283, n_2284, 
      n_2285, n_2286, n_2287, n_2288, n_2289, n_2290, n_2291, n_2292, n_2293, 
      n_2294, n_2295, n_2296, n_2297, n_2298, n_2299, n_2300, n_2301, n_2302, 
      n_2303, n_2304, n_2305, n_2306, n_2307, n_2308, n_2309, n_2310, n_2311, 
      n_2312, n_2313, n_2314, n_2315, n_2316, n_2317, n_2318, n_2319, n_2320, 
      n_2321, n_2322 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   ALU_regmem_reg_0_inst : DFFR_X1 port map( D => ALU_memout_0_port, CK => CLK,
                           RN => n8, Q => ALU_regmem_0_port, QN => n_1978);
   IR_reg_reg_0_inst : DFFR_X1 port map( D => NOP_MUX_OUT_0_port, CK => CLK, RN
                           => n4, Q => IR_reg_0_port, QN => n_1979);
   IR_reg_reg_1_inst : DFFR_X1 port map( D => NOP_MUX_OUT_1_port, CK => CLK, RN
                           => n8, Q => IR_reg_1_port, QN => n_1980);
   IR_reg_reg_2_inst : DFFR_X1 port map( D => NOP_MUX_OUT_2_port, CK => CLK, RN
                           => n8, Q => IR_reg_2_port, QN => n_1981);
   IR_reg_reg_3_inst : DFFR_X1 port map( D => NOP_MUX_OUT_3_port, CK => CLK, RN
                           => n8, Q => IR_reg_3_port, QN => n_1982);
   IR_reg_reg_4_inst : DFFR_X1 port map( D => NOP_MUX_OUT_4_port, CK => CLK, RN
                           => n8, Q => IR_reg_4_port, QN => n_1983);
   IR_reg_reg_5_inst : DFFR_X1 port map( D => NOP_MUX_OUT_5_port, CK => CLK, RN
                           => n8, Q => IR_reg_5_port, QN => n_1984);
   IR_reg_reg_6_inst : DFFR_X1 port map( D => NOP_MUX_OUT_6_port, CK => CLK, RN
                           => n8, Q => IR_reg_6_port, QN => n_1985);
   IR_reg_reg_7_inst : DFFR_X1 port map( D => NOP_MUX_OUT_7_port, CK => CLK, RN
                           => n8, Q => IR_reg_7_port, QN => n_1986);
   IR_reg_reg_8_inst : DFFR_X1 port map( D => NOP_MUX_OUT_8_port, CK => CLK, RN
                           => n8, Q => IR_reg_8_port, QN => n_1987);
   IR_reg_reg_9_inst : DFFR_X1 port map( D => NOP_MUX_OUT_9_port, CK => CLK, RN
                           => n8, Q => IR_reg_9_port, QN => n_1988);
   IR_reg_reg_10_inst : DFFR_X1 port map( D => NOP_MUX_OUT_10_port, CK => CLK, 
                           RN => n8, Q => IR_reg_10_port, QN => n_1989);
   IR_reg_reg_11_inst : DFFR_X1 port map( D => NOP_MUX_OUT_11_port, CK => CLK, 
                           RN => n8, Q => IR_reg_11_port, QN => n_1990);
   IR_reg_reg_12_inst : DFFR_X1 port map( D => NOP_MUX_OUT_12_port, CK => CLK, 
                           RN => n8, Q => IR_reg_12_port, QN => n_1991);
   IR_reg_reg_13_inst : DFFR_X1 port map( D => NOP_MUX_OUT_13_port, CK => CLK, 
                           RN => n7, Q => IR_reg_13_port, QN => n_1992);
   IR_reg_reg_14_inst : DFFR_X1 port map( D => NOP_MUX_OUT_14_port, CK => CLK, 
                           RN => n7, Q => IR_reg_14_port, QN => n_1993);
   IR_reg_reg_15_inst : DFFR_X1 port map( D => NOP_MUX_OUT_15_port, CK => CLK, 
                           RN => n7, Q => IR_reg_15_port, QN => n_1994);
   IR_reg_reg_16_inst : DFFR_X1 port map( D => NOP_MUX_OUT_16_port, CK => CLK, 
                           RN => n7, Q => IR_reg_16_port, QN => n_1995);
   IR_reg_reg_17_inst : DFFR_X1 port map( D => NOP_MUX_OUT_17_port, CK => CLK, 
                           RN => n7, Q => IR_reg_17_port, QN => n_1996);
   IR_reg_reg_18_inst : DFFR_X1 port map( D => NOP_MUX_OUT_18_port, CK => CLK, 
                           RN => n7, Q => IR_reg_18_port, QN => n_1997);
   IR_reg_reg_19_inst : DFFR_X1 port map( D => NOP_MUX_OUT_19_port, CK => CLK, 
                           RN => n7, Q => IR_reg_19_port, QN => n_1998);
   IR_reg_reg_20_inst : DFFR_X1 port map( D => NOP_MUX_OUT_20_port, CK => CLK, 
                           RN => n7, Q => IR_reg_20_port, QN => n_1999);
   IR_reg_reg_21_inst : DFFR_X1 port map( D => NOP_MUX_OUT_21_port, CK => CLK, 
                           RN => n7, Q => IR_reg_21_port, QN => n_2000);
   IR_reg_reg_22_inst : DFFR_X1 port map( D => NOP_MUX_OUT_22_port, CK => CLK, 
                           RN => n7, Q => IR_reg_22_port, QN => n_2001);
   IR_reg_reg_23_inst : DFFR_X1 port map( D => NOP_MUX_OUT_23_port, CK => CLK, 
                           RN => n7, Q => IR_reg_23_port, QN => n_2002);
   IR_reg_reg_24_inst : DFFR_X1 port map( D => NOP_MUX_OUT_24_port, CK => CLK, 
                           RN => n7, Q => IR_reg_24_port, QN => n_2003);
   IR_reg_reg_25_inst : DFFR_X1 port map( D => NOP_MUX_OUT_25_port, CK => CLK, 
                           RN => n7, Q => IR_reg_25_port, QN => n_2004);
   IR_reg_reg_26_inst : DFFS_X1 port map( D => NOP_MUX_OUT_26_port, CK => CLK, 
                           SN => n12, Q => IR_reg_26_port, QN => n_2005);
   IR_reg_reg_27_inst : DFFR_X1 port map( D => NOP_MUX_OUT_27_port, CK => CLK, 
                           RN => n7, Q => IR_reg_27_port, QN => n_2006);
   IR_reg_reg_29_inst : DFFR_X1 port map( D => NOP_MUX_OUT_29_port, CK => CLK, 
                           RN => n7, Q => IR_reg_29_port, QN => n_2007);
   IR_reg_reg_31_inst : DFFR_X1 port map( D => NOP_MUX_OUT_31_port, CK => CLK, 
                           RN => n7, Q => IR_reg_31_port, QN => n_2008);
   NPC_reg_reg_0_inst : DFFR_X1 port map( D => NPC_fetchout_0_port, CK => CLK, 
                           RN => n7, Q => NPC_reg_0_port, QN => n_2009);
   NPC_reg_reg_1_inst : DFFR_X1 port map( D => NPC_fetchout_1_port, CK => CLK, 
                           RN => n7, Q => NPC_reg_1_port, QN => n_2010);
   NPC_reg_reg_2_inst : DFFR_X1 port map( D => NPC_fetchout_2_port, CK => CLK, 
                           RN => n7, Q => NPC_reg_2_port, QN => n_2011);
   NPC_reg_reg_3_inst : DFFR_X1 port map( D => NPC_fetchout_3_port, CK => CLK, 
                           RN => n7, Q => NPC_reg_3_port, QN => n_2012);
   NPC_reg_reg_4_inst : DFFR_X1 port map( D => NPC_fetchout_4_port, CK => CLK, 
                           RN => n7, Q => NPC_reg_4_port, QN => n_2013);
   NPC_reg_reg_5_inst : DFFR_X1 port map( D => NPC_fetchout_5_port, CK => CLK, 
                           RN => n7, Q => NPC_reg_5_port, QN => n_2014);
   NPC_reg_reg_6_inst : DFFR_X1 port map( D => NPC_fetchout_6_port, CK => CLK, 
                           RN => n7, Q => NPC_reg_6_port, QN => n_2015);
   NPC_reg_reg_7_inst : DFFR_X1 port map( D => NPC_fetchout_7_port, CK => CLK, 
                           RN => n7, Q => NPC_reg_7_port, QN => n_2016);
   NPC_reg_reg_8_inst : DFFR_X1 port map( D => NPC_fetchout_8_port, CK => CLK, 
                           RN => n7, Q => NPC_reg_8_port, QN => n_2017);
   NPC_reg_reg_9_inst : DFFR_X1 port map( D => NPC_fetchout_9_port, CK => CLK, 
                           RN => n7, Q => NPC_reg_9_port, QN => n_2018);
   NPC_reg_reg_10_inst : DFFR_X1 port map( D => NPC_fetchout_10_port, CK => CLK
                           , RN => n7, Q => NPC_reg_10_port, QN => n_2019);
   NPC_reg_reg_11_inst : DFFR_X1 port map( D => NPC_fetchout_11_port, CK => CLK
                           , RN => n7, Q => NPC_reg_11_port, QN => n_2020);
   NPC_reg_reg_12_inst : DFFR_X1 port map( D => NPC_fetchout_12_port, CK => CLK
                           , RN => n7, Q => NPC_reg_12_port, QN => n_2021);
   NPC_reg_reg_13_inst : DFFR_X1 port map( D => NPC_fetchout_13_port, CK => CLK
                           , RN => n7, Q => NPC_reg_13_port, QN => n_2022);
   NPC_reg_reg_14_inst : DFFR_X1 port map( D => NPC_fetchout_14_port, CK => CLK
                           , RN => n7, Q => NPC_reg_14_port, QN => n_2023);
   NPC_reg_reg_15_inst : DFFR_X1 port map( D => NPC_fetchout_15_port, CK => CLK
                           , RN => n7, Q => NPC_reg_15_port, QN => n_2024);
   NPC_reg_reg_16_inst : DFFR_X1 port map( D => NPC_fetchout_16_port, CK => CLK
                           , RN => n7, Q => NPC_reg_16_port, QN => n_2025);
   NPC_reg_reg_17_inst : DFFR_X1 port map( D => NPC_fetchout_17_port, CK => CLK
                           , RN => n7, Q => NPC_reg_17_port, QN => n_2026);
   NPC_reg_reg_18_inst : DFFR_X1 port map( D => NPC_fetchout_18_port, CK => CLK
                           , RN => n7, Q => NPC_reg_18_port, QN => n_2027);
   NPC_reg_reg_19_inst : DFFR_X1 port map( D => NPC_fetchout_19_port, CK => CLK
                           , RN => n7, Q => NPC_reg_19_port, QN => n_2028);
   NPC_reg_reg_20_inst : DFFR_X1 port map( D => NPC_fetchout_20_port, CK => CLK
                           , RN => n7, Q => NPC_reg_20_port, QN => n_2029);
   NPC_reg_reg_21_inst : DFFR_X1 port map( D => NPC_fetchout_21_port, CK => CLK
                           , RN => n7, Q => NPC_reg_21_port, QN => n_2030);
   NPC_reg_reg_22_inst : DFFR_X1 port map( D => NPC_fetchout_22_port, CK => CLK
                           , RN => n7, Q => NPC_reg_22_port, QN => n_2031);
   NPC_reg_reg_23_inst : DFFR_X1 port map( D => NPC_fetchout_23_port, CK => CLK
                           , RN => n7, Q => NPC_reg_23_port, QN => n_2032);
   NPC_reg_reg_24_inst : DFFR_X1 port map( D => NPC_fetchout_24_port, CK => CLK
                           , RN => n7, Q => NPC_reg_24_port, QN => n_2033);
   NPC_reg_reg_25_inst : DFFR_X1 port map( D => NPC_fetchout_25_port, CK => CLK
                           , RN => n7, Q => NPC_reg_25_port, QN => n_2034);
   NPC_reg_reg_26_inst : DFFR_X1 port map( D => NPC_fetchout_26_port, CK => CLK
                           , RN => n6, Q => NPC_reg_26_port, QN => n_2035);
   NPC_reg_reg_27_inst : DFFR_X1 port map( D => NPC_fetchout_27_port, CK => CLK
                           , RN => n6, Q => NPC_reg_27_port, QN => n_2036);
   NPC_reg_reg_28_inst : DFFR_X1 port map( D => NPC_fetchout_28_port, CK => CLK
                           , RN => n6, Q => NPC_reg_28_port, QN => n_2037);
   NPC_reg_reg_29_inst : DFFR_X1 port map( D => NPC_fetchout_29_port, CK => CLK
                           , RN => n6, Q => NPC_reg_29_port, QN => n_2038);
   NPC_reg_reg_30_inst : DFFR_X1 port map( D => NPC_fetchout_30_port, CK => CLK
                           , RN => n6, Q => NPC_reg_30_port, QN => n_2039);
   NPC_reg_reg_31_inst : DFFR_X1 port map( D => NPC_fetchout_31_port, CK => CLK
                           , RN => n6, Q => NPC_reg_31_port, QN => n_2040);
   PC_reg_reg_0_inst : DFFR_X1 port map( D => PC_muxout_0_port, CK => CLK, RN 
                           => n6, Q => PC_reg_0_port, QN => n_2041);
   PC_reg_reg_1_inst : DFFR_X1 port map( D => PC_muxout_1_port, CK => CLK, RN 
                           => n6, Q => PC_reg_1_port, QN => n_2042);
   PC_reg_reg_2_inst : DFFR_X1 port map( D => PC_muxout_2_port, CK => CLK, RN 
                           => n6, Q => PC_reg_2_port, QN => n_2043);
   PC_reg_reg_3_inst : DFFR_X1 port map( D => PC_muxout_3_port, CK => CLK, RN 
                           => n6, Q => PC_reg_3_port, QN => n_2044);
   PC_reg_reg_4_inst : DFFR_X1 port map( D => PC_muxout_4_port, CK => CLK, RN 
                           => n6, Q => PC_reg_4_port, QN => n_2045);
   PC_reg_reg_5_inst : DFFR_X1 port map( D => PC_muxout_5_port, CK => CLK, RN 
                           => n6, Q => PC_reg_5_port, QN => n_2046);
   PC_reg_reg_6_inst : DFFR_X1 port map( D => PC_muxout_6_port, CK => CLK, RN 
                           => n6, Q => PC_reg_6_port, QN => n_2047);
   PC_reg_reg_7_inst : DFFR_X1 port map( D => PC_muxout_7_port, CK => CLK, RN 
                           => n6, Q => PC_reg_7_port, QN => n_2048);
   PC_reg_reg_8_inst : DFFR_X1 port map( D => PC_muxout_8_port, CK => CLK, RN 
                           => n6, Q => PC_reg_8_port, QN => n_2049);
   PC_reg_reg_9_inst : DFFR_X1 port map( D => PC_muxout_9_port, CK => CLK, RN 
                           => n6, Q => PC_reg_9_port, QN => n_2050);
   PC_reg_reg_10_inst : DFFR_X1 port map( D => PC_muxout_10_port, CK => CLK, RN
                           => n6, Q => PC_reg_10_port, QN => n_2051);
   PC_reg_reg_11_inst : DFFR_X1 port map( D => PC_muxout_11_port, CK => CLK, RN
                           => n6, Q => PC_reg_11_port, QN => n_2052);
   PC_reg_reg_12_inst : DFFR_X1 port map( D => PC_muxout_12_port, CK => CLK, RN
                           => n6, Q => PC_reg_12_port, QN => n_2053);
   PC_reg_reg_13_inst : DFFR_X1 port map( D => PC_muxout_13_port, CK => CLK, RN
                           => n6, Q => PC_reg_13_port, QN => n_2054);
   PC_reg_reg_14_inst : DFFR_X1 port map( D => PC_muxout_14_port, CK => CLK, RN
                           => n6, Q => PC_reg_14_port, QN => n_2055);
   PC_reg_reg_15_inst : DFFR_X1 port map( D => PC_muxout_15_port, CK => CLK, RN
                           => n6, Q => PC_reg_15_port, QN => n_2056);
   PC_reg_reg_16_inst : DFFR_X1 port map( D => PC_muxout_16_port, CK => CLK, RN
                           => n6, Q => PC_reg_16_port, QN => n_2057);
   PC_reg_reg_17_inst : DFFR_X1 port map( D => PC_muxout_17_port, CK => CLK, RN
                           => n6, Q => PC_reg_17_port, QN => n_2058);
   PC_reg_reg_18_inst : DFFR_X1 port map( D => PC_muxout_18_port, CK => CLK, RN
                           => n6, Q => PC_reg_18_port, QN => n_2059);
   PC_reg_reg_19_inst : DFFR_X1 port map( D => PC_muxout_19_port, CK => CLK, RN
                           => n6, Q => PC_reg_19_port, QN => n_2060);
   PC_reg_reg_20_inst : DFFR_X1 port map( D => PC_muxout_20_port, CK => CLK, RN
                           => n6, Q => PC_reg_20_port, QN => n_2061);
   PC_reg_reg_21_inst : DFFR_X1 port map( D => PC_muxout_21_port, CK => CLK, RN
                           => n6, Q => PC_reg_21_port, QN => n_2062);
   PC_reg_reg_22_inst : DFFR_X1 port map( D => PC_muxout_22_port, CK => CLK, RN
                           => n6, Q => PC_reg_22_port, QN => n_2063);
   PC_reg_reg_23_inst : DFFR_X1 port map( D => PC_muxout_23_port, CK => CLK, RN
                           => n6, Q => PC_reg_23_port, QN => n_2064);
   PC_reg_reg_24_inst : DFFR_X1 port map( D => PC_muxout_24_port, CK => CLK, RN
                           => n6, Q => PC_reg_24_port, QN => n_2065);
   PC_reg_reg_25_inst : DFFR_X1 port map( D => PC_muxout_25_port, CK => CLK, RN
                           => n6, Q => PC_reg_25_port, QN => n_2066);
   PC_reg_reg_26_inst : DFFR_X1 port map( D => PC_muxout_26_port, CK => CLK, RN
                           => n6, Q => PC_reg_26_port, QN => n_2067);
   PC_reg_reg_27_inst : DFFR_X1 port map( D => PC_muxout_27_port, CK => CLK, RN
                           => n6, Q => PC_reg_27_port, QN => n_2068);
   PC_reg_reg_28_inst : DFFR_X1 port map( D => PC_muxout_28_port, CK => CLK, RN
                           => n6, Q => PC_reg_28_port, QN => n_2069);
   PC_reg_reg_29_inst : DFFR_X1 port map( D => PC_muxout_29_port, CK => CLK, RN
                           => n6, Q => PC_reg_29_port, QN => n_2070);
   PC_reg_reg_30_inst : DFFR_X1 port map( D => PC_muxout_30_port, CK => CLK, RN
                           => n6, Q => PC_reg_30_port, QN => n_2071);
   PC_reg_reg_31_inst : DFFR_X1 port map( D => PC_muxout_31_port, CK => CLK, RN
                           => n6, Q => PC_reg_31_port, QN => n_2072);
   RD_regexe_reg_0_inst : DFFR_X1 port map( D => RD_decout_0_port, CK => CLK, 
                           RN => n6, Q => RD_regexe_0_port, QN => n_2073);
   RD_regexe_reg_1_inst : DFFR_X1 port map( D => RD_decout_1_port, CK => CLK, 
                           RN => n6, Q => RD_regexe_1_port, QN => n_2074);
   RD_regexe_reg_2_inst : DFFR_X1 port map( D => RD_decout_2_port, CK => CLK, 
                           RN => n6, Q => RD_regexe_2_port, QN => n_2075);
   RD_regexe_reg_3_inst : DFFR_X1 port map( D => RD_decout_3_port, CK => CLK, 
                           RN => n5, Q => RD_regexe_3_port, QN => n_2076);
   RD_regexe_reg_4_inst : DFFR_X1 port map( D => RD_decout_4_port, CK => CLK, 
                           RN => n5, Q => RD_regexe_4_port, QN => n_2077);
   RSB_reg_reg_0_inst : DFFR_X1 port map( D => RSB_decout_0_port, CK => CLK, RN
                           => n5, Q => RSB_reg_0_port, QN => n_2078);
   RSB_reg_reg_1_inst : DFFR_X1 port map( D => RSB_decout_1_port, CK => CLK, RN
                           => n5, Q => RSB_reg_1_port, QN => n_2079);
   RSB_reg_reg_2_inst : DFFR_X1 port map( D => RSB_decout_2_port, CK => CLK, RN
                           => n5, Q => RSB_reg_2_port, QN => n_2080);
   RSB_reg_reg_3_inst : DFFR_X1 port map( D => RSB_decout_3_port, CK => CLK, RN
                           => n5, Q => RSB_reg_3_port, QN => n_2081);
   RSB_reg_reg_4_inst : DFFR_X1 port map( D => RSB_decout_4_port, CK => CLK, RN
                           => n5, Q => RSB_reg_4_port, QN => n_2082);
   RSA_reg_reg_0_inst : DFFR_X1 port map( D => RSA_decout_0_port, CK => CLK, RN
                           => n5, Q => RSA_reg_0_port, QN => n_2083);
   RSA_reg_reg_1_inst : DFFR_X1 port map( D => RSA_decout_1_port, CK => CLK, RN
                           => n5, Q => RSA_reg_1_port, QN => n_2084);
   RSA_reg_reg_2_inst : DFFR_X1 port map( D => RSA_decout_2_port, CK => CLK, RN
                           => n5, Q => RSA_reg_2_port, QN => n_2085);
   RSA_reg_reg_3_inst : DFFR_X1 port map( D => RSA_decout_3_port, CK => CLK, RN
                           => n5, Q => RSA_reg_3_port, QN => n_2086);
   RSA_reg_reg_4_inst : DFFR_X1 port map( D => RSA_decout_4_port, CK => CLK, RN
                           => n5, Q => RSA_reg_4_port, QN => n_2087);
   RB_reg_reg_0_inst : DFFR_X1 port map( D => RB_decout_0_port, CK => CLK, RN 
                           => n5, Q => RB_reg_0_port, QN => n_2088);
   RB_reg_reg_1_inst : DFFR_X1 port map( D => RB_decout_1_port, CK => CLK, RN 
                           => n5, Q => RB_reg_1_port, QN => n_2089);
   RB_reg_reg_2_inst : DFFR_X1 port map( D => RB_decout_2_port, CK => CLK, RN 
                           => n5, Q => RB_reg_2_port, QN => n_2090);
   RB_reg_reg_3_inst : DFFR_X1 port map( D => RB_decout_3_port, CK => CLK, RN 
                           => n5, Q => RB_reg_3_port, QN => n_2091);
   RB_reg_reg_4_inst : DFFR_X1 port map( D => RB_decout_4_port, CK => CLK, RN 
                           => n5, Q => RB_reg_4_port, QN => n_2092);
   RB_reg_reg_5_inst : DFFR_X1 port map( D => RB_decout_5_port, CK => CLK, RN 
                           => n5, Q => RB_reg_5_port, QN => n_2093);
   RB_reg_reg_6_inst : DFFR_X1 port map( D => RB_decout_6_port, CK => CLK, RN 
                           => n5, Q => RB_reg_6_port, QN => n_2094);
   RB_reg_reg_7_inst : DFFR_X1 port map( D => RB_decout_7_port, CK => CLK, RN 
                           => n5, Q => RB_reg_7_port, QN => n_2095);
   RB_reg_reg_8_inst : DFFR_X1 port map( D => RB_decout_8_port, CK => CLK, RN 
                           => n5, Q => RB_reg_8_port, QN => n_2096);
   RB_reg_reg_9_inst : DFFR_X1 port map( D => RB_decout_9_port, CK => CLK, RN 
                           => n5, Q => RB_reg_9_port, QN => n_2097);
   RB_reg_reg_10_inst : DFFR_X1 port map( D => RB_decout_10_port, CK => CLK, RN
                           => n5, Q => RB_reg_10_port, QN => n_2098);
   RB_reg_reg_11_inst : DFFR_X1 port map( D => RB_decout_11_port, CK => CLK, RN
                           => n5, Q => RB_reg_11_port, QN => n_2099);
   RB_reg_reg_12_inst : DFFR_X1 port map( D => RB_decout_12_port, CK => CLK, RN
                           => n5, Q => RB_reg_12_port, QN => n_2100);
   RB_reg_reg_13_inst : DFFR_X1 port map( D => RB_decout_13_port, CK => CLK, RN
                           => n5, Q => RB_reg_13_port, QN => n_2101);
   RB_reg_reg_14_inst : DFFR_X1 port map( D => RB_decout_14_port, CK => CLK, RN
                           => n5, Q => RB_reg_14_port, QN => n_2102);
   RB_reg_reg_15_inst : DFFR_X1 port map( D => RB_decout_15_port, CK => CLK, RN
                           => n5, Q => RB_reg_15_port, QN => n_2103);
   RB_reg_reg_16_inst : DFFR_X1 port map( D => RB_decout_16_port, CK => CLK, RN
                           => n5, Q => RB_reg_16_port, QN => n_2104);
   RB_reg_reg_17_inst : DFFR_X1 port map( D => RB_decout_17_port, CK => CLK, RN
                           => n5, Q => RB_reg_17_port, QN => n_2105);
   RB_reg_reg_18_inst : DFFR_X1 port map( D => RB_decout_18_port, CK => CLK, RN
                           => n5, Q => RB_reg_18_port, QN => n_2106);
   RB_reg_reg_19_inst : DFFR_X1 port map( D => RB_decout_19_port, CK => CLK, RN
                           => n5, Q => RB_reg_19_port, QN => n_2107);
   RB_reg_reg_20_inst : DFFR_X1 port map( D => RB_decout_20_port, CK => CLK, RN
                           => n5, Q => RB_reg_20_port, QN => n_2108);
   RB_reg_reg_21_inst : DFFR_X1 port map( D => RB_decout_21_port, CK => CLK, RN
                           => n5, Q => RB_reg_21_port, QN => n_2109);
   RB_reg_reg_22_inst : DFFR_X1 port map( D => RB_decout_22_port, CK => CLK, RN
                           => n5, Q => RB_reg_22_port, QN => n_2110);
   RB_reg_reg_23_inst : DFFR_X1 port map( D => RB_decout_23_port, CK => CLK, RN
                           => n5, Q => RB_reg_23_port, QN => n_2111);
   RB_reg_reg_24_inst : DFFR_X1 port map( D => RB_decout_24_port, CK => CLK, RN
                           => n5, Q => RB_reg_24_port, QN => n_2112);
   RB_reg_reg_25_inst : DFFR_X1 port map( D => RB_decout_25_port, CK => CLK, RN
                           => n5, Q => RB_reg_25_port, QN => n_2113);
   RB_reg_reg_26_inst : DFFR_X1 port map( D => RB_decout_26_port, CK => CLK, RN
                           => n5, Q => RB_reg_26_port, QN => n_2114);
   RB_reg_reg_27_inst : DFFR_X1 port map( D => RB_decout_27_port, CK => CLK, RN
                           => n5, Q => RB_reg_27_port, QN => n_2115);
   RB_reg_reg_28_inst : DFFR_X1 port map( D => RB_decout_28_port, CK => CLK, RN
                           => n5, Q => RB_reg_28_port, QN => n_2116);
   RB_reg_reg_29_inst : DFFR_X1 port map( D => RB_decout_29_port, CK => CLK, RN
                           => n5, Q => RB_reg_29_port, QN => n_2117);
   RB_reg_reg_30_inst : DFFR_X1 port map( D => RB_decout_30_port, CK => CLK, RN
                           => n4, Q => RB_reg_30_port, QN => n_2118);
   RB_reg_reg_31_inst : DFFR_X1 port map( D => RB_decout_31_port, CK => CLK, RN
                           => n4, Q => RB_reg_31_port, QN => n_2119);
   RA_reg_reg_0_inst : DFFR_X1 port map( D => RA_decout_0_port, CK => CLK, RN 
                           => n4, Q => RA_reg_0_port, QN => n_2120);
   RA_reg_reg_1_inst : DFFR_X1 port map( D => RA_decout_1_port, CK => CLK, RN 
                           => n4, Q => RA_reg_1_port, QN => n_2121);
   RA_reg_reg_2_inst : DFFR_X1 port map( D => RA_decout_2_port, CK => CLK, RN 
                           => n4, Q => RA_reg_2_port, QN => n_2122);
   RA_reg_reg_3_inst : DFFR_X1 port map( D => RA_decout_3_port, CK => CLK, RN 
                           => n4, Q => RA_reg_3_port, QN => n_2123);
   RA_reg_reg_4_inst : DFFR_X1 port map( D => RA_decout_4_port, CK => CLK, RN 
                           => n4, Q => RA_reg_4_port, QN => n_2124);
   RA_reg_reg_5_inst : DFFR_X1 port map( D => RA_decout_5_port, CK => CLK, RN 
                           => n4, Q => RA_reg_5_port, QN => n_2125);
   RA_reg_reg_6_inst : DFFR_X1 port map( D => RA_decout_6_port, CK => CLK, RN 
                           => n4, Q => RA_reg_6_port, QN => n_2126);
   RA_reg_reg_7_inst : DFFR_X1 port map( D => RA_decout_7_port, CK => CLK, RN 
                           => n4, Q => RA_reg_7_port, QN => n_2127);
   RA_reg_reg_8_inst : DFFR_X1 port map( D => RA_decout_8_port, CK => CLK, RN 
                           => n4, Q => RA_reg_8_port, QN => n_2128);
   RA_reg_reg_9_inst : DFFR_X1 port map( D => RA_decout_9_port, CK => CLK, RN 
                           => n4, Q => RA_reg_9_port, QN => n_2129);
   RA_reg_reg_10_inst : DFFR_X1 port map( D => RA_decout_10_port, CK => CLK, RN
                           => n4, Q => RA_reg_10_port, QN => n_2130);
   RA_reg_reg_11_inst : DFFR_X1 port map( D => RA_decout_11_port, CK => CLK, RN
                           => n4, Q => RA_reg_11_port, QN => n_2131);
   RA_reg_reg_12_inst : DFFR_X1 port map( D => RA_decout_12_port, CK => CLK, RN
                           => n4, Q => RA_reg_12_port, QN => n_2132);
   RA_reg_reg_13_inst : DFFR_X1 port map( D => RA_decout_13_port, CK => CLK, RN
                           => n4, Q => RA_reg_13_port, QN => n_2133);
   RA_reg_reg_14_inst : DFFR_X1 port map( D => RA_decout_14_port, CK => CLK, RN
                           => n4, Q => RA_reg_14_port, QN => n_2134);
   RA_reg_reg_15_inst : DFFR_X1 port map( D => RA_decout_15_port, CK => CLK, RN
                           => n4, Q => RA_reg_15_port, QN => n_2135);
   RA_reg_reg_16_inst : DFFR_X1 port map( D => RA_decout_16_port, CK => CLK, RN
                           => n4, Q => RA_reg_16_port, QN => n_2136);
   RA_reg_reg_17_inst : DFFR_X1 port map( D => RA_decout_17_port, CK => CLK, RN
                           => n4, Q => RA_reg_17_port, QN => n_2137);
   RA_reg_reg_18_inst : DFFR_X1 port map( D => RA_decout_18_port, CK => CLK, RN
                           => n4, Q => RA_reg_18_port, QN => n_2138);
   RA_reg_reg_19_inst : DFFR_X1 port map( D => RA_decout_19_port, CK => CLK, RN
                           => n4, Q => RA_reg_19_port, QN => n_2139);
   RA_reg_reg_20_inst : DFFR_X1 port map( D => RA_decout_20_port, CK => CLK, RN
                           => n4, Q => RA_reg_20_port, QN => n_2140);
   RA_reg_reg_21_inst : DFFR_X1 port map( D => RA_decout_21_port, CK => CLK, RN
                           => n4, Q => RA_reg_21_port, QN => n_2141);
   RA_reg_reg_22_inst : DFFR_X1 port map( D => RA_decout_22_port, CK => CLK, RN
                           => n4, Q => RA_reg_22_port, QN => n_2142);
   RA_reg_reg_23_inst : DFFR_X1 port map( D => RA_decout_23_port, CK => CLK, RN
                           => n4, Q => RA_reg_23_port, QN => n_2143);
   RA_reg_reg_24_inst : DFFR_X1 port map( D => RA_decout_24_port, CK => CLK, RN
                           => n4, Q => RA_reg_24_port, QN => n_2144);
   RA_reg_reg_25_inst : DFFR_X1 port map( D => RA_decout_25_port, CK => CLK, RN
                           => n4, Q => RA_reg_25_port, QN => n_2145);
   RA_reg_reg_26_inst : DFFR_X1 port map( D => RA_decout_26_port, CK => CLK, RN
                           => n4, Q => RA_reg_26_port, QN => n_2146);
   RA_reg_reg_27_inst : DFFR_X1 port map( D => RA_decout_27_port, CK => CLK, RN
                           => n4, Q => RA_reg_27_port, QN => n_2147);
   RA_reg_reg_28_inst : DFFR_X1 port map( D => RA_decout_28_port, CK => CLK, RN
                           => n4, Q => RA_reg_28_port, QN => n_2148);
   RA_reg_reg_29_inst : DFFR_X1 port map( D => RA_decout_29_port, CK => CLK, RN
                           => n4, Q => RA_reg_29_port, QN => n_2149);
   RA_reg_reg_30_inst : DFFR_X1 port map( D => RA_decout_30_port, CK => CLK, RN
                           => n6, Q => RA_reg_30_port, QN => n_2150);
   RA_reg_reg_31_inst : DFFR_X1 port map( D => RA_decout_31_port, CK => CLK, RN
                           => n12, Q => RA_reg_31_port, QN => n_2151);
   Imm_reg_reg_0_inst : DFFR_X1 port map( D => IMM_decout_0_port, CK => CLK, RN
                           => n12, Q => Imm_reg_0_port, QN => n_2152);
   Imm_reg_reg_1_inst : DFFR_X1 port map( D => IMM_decout_1_port, CK => CLK, RN
                           => n12, Q => Imm_reg_1_port, QN => n_2153);
   Imm_reg_reg_2_inst : DFFR_X1 port map( D => IMM_decout_2_port, CK => CLK, RN
                           => n12, Q => Imm_reg_2_port, QN => n_2154);
   Imm_reg_reg_3_inst : DFFR_X1 port map( D => IMM_decout_3_port, CK => CLK, RN
                           => n12, Q => Imm_reg_3_port, QN => n_2155);
   Imm_reg_reg_4_inst : DFFR_X1 port map( D => IMM_decout_4_port, CK => CLK, RN
                           => n12, Q => Imm_reg_4_port, QN => n_2156);
   Imm_reg_reg_5_inst : DFFR_X1 port map( D => IMM_decout_5_port, CK => CLK, RN
                           => n12, Q => Imm_reg_5_port, QN => n_2157);
   Imm_reg_reg_6_inst : DFFR_X1 port map( D => IMM_decout_6_port, CK => CLK, RN
                           => n12, Q => Imm_reg_6_port, QN => n_2158);
   Imm_reg_reg_7_inst : DFFR_X1 port map( D => IMM_decout_7_port, CK => CLK, RN
                           => n12, Q => Imm_reg_7_port, QN => n_2159);
   Imm_reg_reg_8_inst : DFFR_X1 port map( D => IMM_decout_8_port, CK => CLK, RN
                           => n12, Q => Imm_reg_8_port, QN => n_2160);
   Imm_reg_reg_9_inst : DFFR_X1 port map( D => IMM_decout_9_port, CK => CLK, RN
                           => n12, Q => Imm_reg_9_port, QN => n_2161);
   Imm_reg_reg_10_inst : DFFR_X1 port map( D => IMM_decout_10_port, CK => CLK, 
                           RN => n12, Q => Imm_reg_10_port, QN => n_2162);
   Imm_reg_reg_11_inst : DFFR_X1 port map( D => IMM_decout_11_port, CK => CLK, 
                           RN => n11, Q => Imm_reg_11_port, QN => n_2163);
   Imm_reg_reg_12_inst : DFFR_X1 port map( D => IMM_decout_12_port, CK => CLK, 
                           RN => n12, Q => Imm_reg_12_port, QN => n_2164);
   Imm_reg_reg_13_inst : DFFR_X1 port map( D => IMM_decout_13_port, CK => CLK, 
                           RN => n12, Q => Imm_reg_13_port, QN => n_2165);
   Imm_reg_reg_14_inst : DFFR_X1 port map( D => IMM_decout_14_port, CK => CLK, 
                           RN => n11, Q => Imm_reg_14_port, QN => n_2166);
   Imm_reg_reg_15_inst : DFFR_X1 port map( D => IMM_decout_15_port, CK => CLK, 
                           RN => n12, Q => Imm_reg_15_port, QN => n_2167);
   Imm_reg_reg_16_inst : DFFR_X1 port map( D => IMM_decout_16_port, CK => CLK, 
                           RN => n11, Q => Imm_reg_16_port, QN => n_2168);
   Imm_reg_reg_17_inst : DFFR_X1 port map( D => IMM_decout_17_port, CK => CLK, 
                           RN => n11, Q => Imm_reg_17_port, QN => n_2169);
   Imm_reg_reg_18_inst : DFFR_X1 port map( D => IMM_decout_18_port, CK => CLK, 
                           RN => n11, Q => Imm_reg_18_port, QN => n_2170);
   Imm_reg_reg_19_inst : DFFR_X1 port map( D => IMM_decout_19_port, CK => CLK, 
                           RN => n11, Q => Imm_reg_19_port, QN => n_2171);
   Imm_reg_reg_20_inst : DFFR_X1 port map( D => IMM_decout_20_port, CK => CLK, 
                           RN => n11, Q => Imm_reg_20_port, QN => n_2172);
   Imm_reg_reg_21_inst : DFFR_X1 port map( D => IMM_decout_21_port, CK => CLK, 
                           RN => n11, Q => Imm_reg_21_port, QN => n_2173);
   Imm_reg_reg_22_inst : DFFR_X1 port map( D => IMM_decout_22_port, CK => CLK, 
                           RN => n11, Q => Imm_reg_22_port, QN => n_2174);
   Imm_reg_reg_23_inst : DFFR_X1 port map( D => IMM_decout_23_port, CK => CLK, 
                           RN => n11, Q => Imm_reg_23_port, QN => n_2175);
   Imm_reg_reg_24_inst : DFFR_X1 port map( D => IMM_decout_24_port, CK => CLK, 
                           RN => n11, Q => Imm_reg_24_port, QN => n_2176);
   Imm_reg_reg_25_inst : DFFR_X1 port map( D => IMM_decout_25_port, CK => CLK, 
                           RN => n11, Q => Imm_reg_25_port, QN => n_2177);
   Imm_reg_reg_26_inst : DFFR_X1 port map( D => IMM_decout_26_port, CK => CLK, 
                           RN => n11, Q => Imm_reg_26_port, QN => n_2178);
   Imm_reg_reg_27_inst : DFFR_X1 port map( D => IMM_decout_27_port, CK => CLK, 
                           RN => n11, Q => Imm_reg_27_port, QN => n_2179);
   Imm_reg_reg_28_inst : DFFR_X1 port map( D => IMM_decout_28_port, CK => CLK, 
                           RN => n11, Q => Imm_reg_28_port, QN => n_2180);
   Imm_reg_reg_29_inst : DFFR_X1 port map( D => IMM_decout_29_port, CK => CLK, 
                           RN => n11, Q => Imm_reg_29_port, QN => n_2181);
   Imm_reg_reg_30_inst : DFFR_X1 port map( D => IMM_decout_30_port, CK => CLK, 
                           RN => n11, Q => Imm_reg_30_port, QN => n_2182);
   Imm_reg_reg_31_inst : DFFR_X1 port map( D => IMM_decout_31_port, CK => CLK, 
                           RN => n11, Q => Imm_reg_31_port, QN => n_2183);
   RD_regmem_reg_0_inst : DFFR_X1 port map( D => RD_exeout_0_port, CK => CLK, 
                           RN => n11, Q => RD_regmem_0_port, QN => n_2184);
   RD_regmem_reg_1_inst : DFFR_X1 port map( D => RD_exeout_1_port, CK => CLK, 
                           RN => n11, Q => RD_regmem_1_port, QN => n_2185);
   RD_regmem_reg_2_inst : DFFR_X1 port map( D => RD_exeout_2_port, CK => CLK, 
                           RN => n11, Q => RD_regmem_2_port, QN => n_2186);
   RD_regmem_reg_3_inst : DFFR_X1 port map( D => RD_exeout_3_port, CK => CLK, 
                           RN => n11, Q => RD_regmem_3_port, QN => n_2187);
   RD_regmem_reg_4_inst : DFFR_X1 port map( D => RD_exeout_4_port, CK => CLK, 
                           RN => n11, Q => RD_regmem_4_port, QN => n_2188);
   ME_reg_reg_0_inst : DFFR_X1 port map( D => ME_exeout_0_port, CK => CLK, RN 
                           => n11, Q => ME_reg_0_port, QN => n_2189);
   ME_reg_reg_1_inst : DFFR_X1 port map( D => ME_exeout_1_port, CK => CLK, RN 
                           => n11, Q => ME_reg_1_port, QN => n_2190);
   ME_reg_reg_2_inst : DFFR_X1 port map( D => ME_exeout_2_port, CK => CLK, RN 
                           => n11, Q => ME_reg_2_port, QN => n_2191);
   ME_reg_reg_3_inst : DFFR_X1 port map( D => ME_exeout_3_port, CK => CLK, RN 
                           => n11, Q => ME_reg_3_port, QN => n_2192);
   ME_reg_reg_4_inst : DFFR_X1 port map( D => ME_exeout_4_port, CK => CLK, RN 
                           => n11, Q => ME_reg_4_port, QN => n_2193);
   ME_reg_reg_5_inst : DFFR_X1 port map( D => ME_exeout_5_port, CK => CLK, RN 
                           => n11, Q => ME_reg_5_port, QN => n_2194);
   ME_reg_reg_6_inst : DFFR_X1 port map( D => ME_exeout_6_port, CK => CLK, RN 
                           => n11, Q => ME_reg_6_port, QN => n_2195);
   ME_reg_reg_7_inst : DFFR_X1 port map( D => ME_exeout_7_port, CK => CLK, RN 
                           => n11, Q => ME_reg_7_port, QN => n_2196);
   ME_reg_reg_8_inst : DFFR_X1 port map( D => ME_exeout_8_port, CK => CLK, RN 
                           => n11, Q => ME_reg_8_port, QN => n_2197);
   ME_reg_reg_9_inst : DFFR_X1 port map( D => ME_exeout_9_port, CK => CLK, RN 
                           => n11, Q => ME_reg_9_port, QN => n_2198);
   ME_reg_reg_10_inst : DFFR_X1 port map( D => ME_exeout_10_port, CK => CLK, RN
                           => n11, Q => ME_reg_10_port, QN => n_2199);
   ME_reg_reg_11_inst : DFFR_X1 port map( D => ME_exeout_11_port, CK => CLK, RN
                           => n11, Q => ME_reg_11_port, QN => n_2200);
   ME_reg_reg_12_inst : DFFR_X1 port map( D => ME_exeout_12_port, CK => CLK, RN
                           => n11, Q => ME_reg_12_port, QN => n_2201);
   ME_reg_reg_13_inst : DFFR_X1 port map( D => ME_exeout_13_port, CK => CLK, RN
                           => n11, Q => ME_reg_13_port, QN => n_2202);
   ME_reg_reg_14_inst : DFFR_X1 port map( D => ME_exeout_14_port, CK => CLK, RN
                           => n11, Q => ME_reg_14_port, QN => n_2203);
   ME_reg_reg_15_inst : DFFR_X1 port map( D => ME_exeout_15_port, CK => CLK, RN
                           => n11, Q => ME_reg_15_port, QN => n_2204);
   ME_reg_reg_16_inst : DFFR_X1 port map( D => ME_exeout_16_port, CK => CLK, RN
                           => n11, Q => ME_reg_16_port, QN => n_2205);
   ME_reg_reg_17_inst : DFFR_X1 port map( D => ME_exeout_17_port, CK => CLK, RN
                           => n11, Q => ME_reg_17_port, QN => n_2206);
   ME_reg_reg_18_inst : DFFR_X1 port map( D => ME_exeout_18_port, CK => CLK, RN
                           => n11, Q => ME_reg_18_port, QN => n_2207);
   ME_reg_reg_19_inst : DFFR_X1 port map( D => ME_exeout_19_port, CK => CLK, RN
                           => n10, Q => ME_reg_19_port, QN => n_2208);
   ME_reg_reg_20_inst : DFFR_X1 port map( D => ME_exeout_20_port, CK => CLK, RN
                           => n10, Q => ME_reg_20_port, QN => n_2209);
   ME_reg_reg_21_inst : DFFR_X1 port map( D => ME_exeout_21_port, CK => CLK, RN
                           => n10, Q => ME_reg_21_port, QN => n_2210);
   ME_reg_reg_22_inst : DFFR_X1 port map( D => ME_exeout_22_port, CK => CLK, RN
                           => n10, Q => ME_reg_22_port, QN => n_2211);
   ME_reg_reg_23_inst : DFFR_X1 port map( D => ME_exeout_23_port, CK => CLK, RN
                           => n10, Q => ME_reg_23_port, QN => n_2212);
   ME_reg_reg_24_inst : DFFR_X1 port map( D => ME_exeout_24_port, CK => CLK, RN
                           => n10, Q => ME_reg_24_port, QN => n_2213);
   ME_reg_reg_25_inst : DFFR_X1 port map( D => ME_exeout_25_port, CK => CLK, RN
                           => n10, Q => ME_reg_25_port, QN => n_2214);
   ME_reg_reg_26_inst : DFFR_X1 port map( D => ME_exeout_26_port, CK => CLK, RN
                           => n10, Q => ME_reg_26_port, QN => n_2215);
   ME_reg_reg_27_inst : DFFR_X1 port map( D => ME_exeout_27_port, CK => CLK, RN
                           => n10, Q => ME_reg_27_port, QN => n_2216);
   ME_reg_reg_28_inst : DFFR_X1 port map( D => ME_exeout_28_port, CK => CLK, RN
                           => n10, Q => ME_reg_28_port, QN => n_2217);
   ME_reg_reg_29_inst : DFFR_X1 port map( D => ME_exeout_29_port, CK => CLK, RN
                           => n10, Q => ME_reg_29_port, QN => n_2218);
   ME_reg_reg_30_inst : DFFR_X1 port map( D => ME_exeout_30_port, CK => CLK, RN
                           => n10, Q => ME_reg_30_port, QN => n_2219);
   ME_reg_reg_31_inst : DFFR_X1 port map( D => ME_exeout_31_port, CK => CLK, RN
                           => n10, Q => ME_reg_31_port, QN => n_2220);
   ALU_reg_reg_0_inst : DFFR_X1 port map( D => ALU_exeout_0_port, CK => CLK, RN
                           => n10, Q => ALU_reg_0_port, QN => n_2221);
   ALU_reg_reg_1_inst : DFFR_X1 port map( D => ALU_exeout_1_port, CK => CLK, RN
                           => n10, Q => ALU_reg_1_port, QN => n_2222);
   ALU_reg_reg_2_inst : DFFR_X1 port map( D => ALU_exeout_2_port, CK => CLK, RN
                           => n10, Q => ALU_reg_2_port, QN => n_2223);
   ALU_reg_reg_3_inst : DFFR_X1 port map( D => ALU_exeout_3_port, CK => CLK, RN
                           => n10, Q => ALU_reg_3_port, QN => n_2224);
   ALU_reg_reg_4_inst : DFFR_X1 port map( D => ALU_exeout_4_port, CK => CLK, RN
                           => n10, Q => ALU_reg_4_port, QN => n_2225);
   ALU_reg_reg_5_inst : DFFR_X1 port map( D => ALU_exeout_5_port, CK => CLK, RN
                           => n10, Q => ALU_reg_5_port, QN => n_2226);
   ALU_reg_reg_6_inst : DFFR_X1 port map( D => ALU_exeout_6_port, CK => CLK, RN
                           => n10, Q => ALU_reg_6_port, QN => n_2227);
   ALU_reg_reg_7_inst : DFFR_X1 port map( D => ALU_exeout_7_port, CK => CLK, RN
                           => n10, Q => ALU_reg_7_port, QN => n_2228);
   ALU_reg_reg_8_inst : DFFR_X1 port map( D => ALU_exeout_8_port, CK => CLK, RN
                           => n10, Q => ALU_reg_8_port, QN => n_2229);
   ALU_reg_reg_9_inst : DFFR_X1 port map( D => ALU_exeout_9_port, CK => CLK, RN
                           => n10, Q => ALU_reg_9_port, QN => n_2230);
   ALU_reg_reg_10_inst : DFFR_X1 port map( D => ALU_exeout_10_port, CK => CLK, 
                           RN => n10, Q => ALU_reg_10_port, QN => n_2231);
   ALU_reg_reg_11_inst : DFFR_X1 port map( D => ALU_exeout_11_port, CK => CLK, 
                           RN => n10, Q => ALU_reg_11_port, QN => n_2232);
   ALU_reg_reg_12_inst : DFFR_X1 port map( D => ALU_exeout_12_port, CK => CLK, 
                           RN => n10, Q => ALU_reg_12_port, QN => n_2233);
   ALU_reg_reg_13_inst : DFFR_X1 port map( D => ALU_exeout_13_port, CK => CLK, 
                           RN => n10, Q => ALU_reg_13_port, QN => n_2234);
   ALU_reg_reg_14_inst : DFFR_X1 port map( D => ALU_exeout_14_port, CK => CLK, 
                           RN => n10, Q => ALU_reg_14_port, QN => n_2235);
   ALU_reg_reg_15_inst : DFFR_X1 port map( D => ALU_exeout_15_port, CK => CLK, 
                           RN => n10, Q => ALU_reg_15_port, QN => n_2236);
   ALU_reg_reg_16_inst : DFFR_X1 port map( D => ALU_exeout_16_port, CK => CLK, 
                           RN => n10, Q => ALU_reg_16_port, QN => n_2237);
   ALU_reg_reg_17_inst : DFFR_X1 port map( D => ALU_exeout_17_port, CK => CLK, 
                           RN => n10, Q => ALU_reg_17_port, QN => n_2238);
   ALU_reg_reg_18_inst : DFFR_X1 port map( D => ALU_exeout_18_port, CK => CLK, 
                           RN => n10, Q => ALU_reg_18_port, QN => n_2239);
   ALU_reg_reg_19_inst : DFFR_X1 port map( D => ALU_exeout_19_port, CK => CLK, 
                           RN => n10, Q => ALU_reg_19_port, QN => n_2240);
   ALU_reg_reg_20_inst : DFFR_X1 port map( D => ALU_exeout_20_port, CK => CLK, 
                           RN => n10, Q => ALU_reg_20_port, QN => n_2241);
   ALU_reg_reg_21_inst : DFFR_X1 port map( D => ALU_exeout_21_port, CK => CLK, 
                           RN => n10, Q => ALU_reg_21_port, QN => n_2242);
   ALU_reg_reg_22_inst : DFFR_X1 port map( D => ALU_exeout_22_port, CK => CLK, 
                           RN => n10, Q => ALU_reg_22_port, QN => n_2243);
   ALU_reg_reg_23_inst : DFFR_X1 port map( D => ALU_exeout_23_port, CK => CLK, 
                           RN => n10, Q => ALU_reg_23_port, QN => n_2244);
   ALU_reg_reg_24_inst : DFFR_X1 port map( D => ALU_exeout_24_port, CK => CLK, 
                           RN => n10, Q => ALU_reg_24_port, QN => n_2245);
   ALU_reg_reg_25_inst : DFFR_X1 port map( D => ALU_exeout_25_port, CK => CLK, 
                           RN => n10, Q => ALU_reg_25_port, QN => n_2246);
   ALU_reg_reg_26_inst : DFFR_X1 port map( D => ALU_exeout_26_port, CK => CLK, 
                           RN => n10, Q => ALU_reg_26_port, QN => n_2247);
   ALU_reg_reg_27_inst : DFFR_X1 port map( D => ALU_exeout_27_port, CK => CLK, 
                           RN => n10, Q => ALU_reg_27_port, QN => n_2248);
   ALU_reg_reg_28_inst : DFFR_X1 port map( D => ALU_exeout_28_port, CK => CLK, 
                           RN => n9, Q => ALU_reg_28_port, QN => n_2249);
   ALU_reg_reg_29_inst : DFFR_X1 port map( D => ALU_exeout_29_port, CK => CLK, 
                           RN => n9, Q => ALU_reg_29_port, QN => n_2250);
   ALU_reg_reg_30_inst : DFFR_X1 port map( D => ALU_exeout_30_port, CK => CLK, 
                           RN => n9, Q => ALU_reg_30_port, QN => n_2251);
   ALU_reg_reg_31_inst : DFFR_X1 port map( D => ALU_exeout_31_port, CK => CLK, 
                           RN => n9, Q => ALU_reg_31_port, QN => n_2252);
   RD_regwb_reg_0_inst : DFFR_X1 port map( D => RD_memout_0_port, CK => CLK, RN
                           => n9, Q => RD_regwb_0_port, QN => n_2253);
   RD_regwb_reg_1_inst : DFFR_X1 port map( D => RD_memout_1_port, CK => CLK, RN
                           => n9, Q => RD_regwb_1_port, QN => n_2254);
   RD_regwb_reg_2_inst : DFFR_X1 port map( D => RD_memout_2_port, CK => CLK, RN
                           => n9, Q => RD_regwb_2_port, QN => n_2255);
   RD_regwb_reg_3_inst : DFFR_X1 port map( D => RD_memout_3_port, CK => CLK, RN
                           => n9, Q => RD_regwb_3_port, QN => n_2256);
   RD_regwb_reg_4_inst : DFFR_X1 port map( D => RD_memout_4_port, CK => CLK, RN
                           => n9, Q => RD_regwb_4_port, QN => n_2257);
   ALU_regmem_reg_1_inst : DFFR_X1 port map( D => ALU_memout_1_port, CK => CLK,
                           RN => n9, Q => ALU_regmem_1_port, QN => n_2258);
   ALU_regmem_reg_2_inst : DFFR_X1 port map( D => ALU_memout_2_port, CK => CLK,
                           RN => n9, Q => ALU_regmem_2_port, QN => n_2259);
   ALU_regmem_reg_3_inst : DFFR_X1 port map( D => ALU_memout_3_port, CK => CLK,
                           RN => n9, Q => ALU_regmem_3_port, QN => n_2260);
   ALU_regmem_reg_4_inst : DFFR_X1 port map( D => ALU_memout_4_port, CK => CLK,
                           RN => n9, Q => ALU_regmem_4_port, QN => n_2261);
   ALU_regmem_reg_5_inst : DFFR_X1 port map( D => ALU_memout_5_port, CK => CLK,
                           RN => n9, Q => ALU_regmem_5_port, QN => n_2262);
   ALU_regmem_reg_6_inst : DFFR_X1 port map( D => ALU_memout_6_port, CK => CLK,
                           RN => n9, Q => ALU_regmem_6_port, QN => n_2263);
   ALU_regmem_reg_7_inst : DFFR_X1 port map( D => ALU_memout_7_port, CK => CLK,
                           RN => n9, Q => ALU_regmem_7_port, QN => n_2264);
   ALU_regmem_reg_8_inst : DFFR_X1 port map( D => ALU_memout_8_port, CK => CLK,
                           RN => n9, Q => ALU_regmem_8_port, QN => n_2265);
   ALU_regmem_reg_9_inst : DFFR_X1 port map( D => ALU_memout_9_port, CK => CLK,
                           RN => n9, Q => ALU_regmem_9_port, QN => n_2266);
   ALU_regmem_reg_10_inst : DFFR_X1 port map( D => ALU_memout_10_port, CK => 
                           CLK, RN => n9, Q => ALU_regmem_10_port, QN => n_2267
                           );
   ALU_regmem_reg_11_inst : DFFR_X1 port map( D => ALU_memout_11_port, CK => 
                           CLK, RN => n9, Q => ALU_regmem_11_port, QN => n_2268
                           );
   ALU_regmem_reg_12_inst : DFFR_X1 port map( D => ALU_memout_12_port, CK => 
                           CLK, RN => n9, Q => ALU_regmem_12_port, QN => n_2269
                           );
   ALU_regmem_reg_13_inst : DFFR_X1 port map( D => ALU_memout_13_port, CK => 
                           CLK, RN => n9, Q => ALU_regmem_13_port, QN => n_2270
                           );
   ALU_regmem_reg_14_inst : DFFR_X1 port map( D => ALU_memout_14_port, CK => 
                           CLK, RN => n9, Q => ALU_regmem_14_port, QN => n_2271
                           );
   ALU_regmem_reg_15_inst : DFFR_X1 port map( D => ALU_memout_15_port, CK => 
                           CLK, RN => n9, Q => ALU_regmem_15_port, QN => n_2272
                           );
   ALU_regmem_reg_16_inst : DFFR_X1 port map( D => ALU_memout_16_port, CK => 
                           CLK, RN => n9, Q => ALU_regmem_16_port, QN => n_2273
                           );
   ALU_regmem_reg_17_inst : DFFR_X1 port map( D => ALU_memout_17_port, CK => 
                           CLK, RN => n9, Q => ALU_regmem_17_port, QN => n_2274
                           );
   ALU_regmem_reg_18_inst : DFFR_X1 port map( D => ALU_memout_18_port, CK => 
                           CLK, RN => n9, Q => ALU_regmem_18_port, QN => n_2275
                           );
   ALU_regmem_reg_19_inst : DFFR_X1 port map( D => ALU_memout_19_port, CK => 
                           CLK, RN => n9, Q => ALU_regmem_19_port, QN => n_2276
                           );
   ALU_regmem_reg_20_inst : DFFR_X1 port map( D => ALU_memout_20_port, CK => 
                           CLK, RN => n9, Q => ALU_regmem_20_port, QN => n_2277
                           );
   ALU_regmem_reg_21_inst : DFFR_X1 port map( D => ALU_memout_21_port, CK => 
                           CLK, RN => n9, Q => ALU_regmem_21_port, QN => n_2278
                           );
   ALU_regmem_reg_22_inst : DFFR_X1 port map( D => ALU_memout_22_port, CK => 
                           CLK, RN => n9, Q => ALU_regmem_22_port, QN => n_2279
                           );
   ALU_regmem_reg_23_inst : DFFR_X1 port map( D => ALU_memout_23_port, CK => 
                           CLK, RN => n9, Q => ALU_regmem_23_port, QN => n_2280
                           );
   ALU_regmem_reg_24_inst : DFFR_X1 port map( D => ALU_memout_24_port, CK => 
                           CLK, RN => n9, Q => ALU_regmem_24_port, QN => n_2281
                           );
   ALU_regmem_reg_25_inst : DFFR_X1 port map( D => ALU_memout_25_port, CK => 
                           CLK, RN => n10, Q => ALU_regmem_25_port, QN => 
                           n_2282);
   ALU_regmem_reg_26_inst : DFFR_X1 port map( D => ALU_memout_26_port, CK => 
                           CLK, RN => n9, Q => ALU_regmem_26_port, QN => n_2283
                           );
   ALU_regmem_reg_27_inst : DFFR_X1 port map( D => ALU_memout_27_port, CK => 
                           CLK, RN => n9, Q => ALU_regmem_27_port, QN => n_2284
                           );
   ALU_regmem_reg_28_inst : DFFR_X1 port map( D => ALU_memout_28_port, CK => 
                           CLK, RN => n9, Q => ALU_regmem_28_port, QN => n_2285
                           );
   ALU_regmem_reg_29_inst : DFFR_X1 port map( D => ALU_memout_29_port, CK => 
                           CLK, RN => n9, Q => ALU_regmem_29_port, QN => n_2286
                           );
   ALU_regmem_reg_30_inst : DFFR_X1 port map( D => ALU_memout_30_port, CK => 
                           CLK, RN => n9, Q => ALU_regmem_30_port, QN => n_2287
                           );
   ALU_regmem_reg_31_inst : DFFR_X1 port map( D => ALU_memout_31_port, CK => 
                           CLK, RN => n9, Q => ALU_regmem_31_port, QN => n_2288
                           );
   LMD_reg_reg_0_inst : DFFR_X1 port map( D => mem_out_0_port, CK => CLK, RN =>
                           n9, Q => LMD_reg_0_port, QN => n_2289);
   LMD_reg_reg_1_inst : DFFR_X1 port map( D => mem_out_1_port, CK => CLK, RN =>
                           n9, Q => LMD_reg_1_port, QN => n_2290);
   LMD_reg_reg_2_inst : DFFR_X1 port map( D => mem_out_2_port, CK => CLK, RN =>
                           n9, Q => LMD_reg_2_port, QN => n_2291);
   LMD_reg_reg_3_inst : DFFR_X1 port map( D => mem_out_3_port, CK => CLK, RN =>
                           n8, Q => LMD_reg_3_port, QN => n_2292);
   LMD_reg_reg_4_inst : DFFR_X1 port map( D => mem_out_4_port, CK => CLK, RN =>
                           n8, Q => LMD_reg_4_port, QN => n_2293);
   LMD_reg_reg_5_inst : DFFR_X1 port map( D => mem_out_5_port, CK => CLK, RN =>
                           n8, Q => LMD_reg_5_port, QN => n_2294);
   LMD_reg_reg_6_inst : DFFR_X1 port map( D => mem_out_6_port, CK => CLK, RN =>
                           n8, Q => LMD_reg_6_port, QN => n_2295);
   LMD_reg_reg_7_inst : DFFR_X1 port map( D => mem_out_7_port, CK => CLK, RN =>
                           n8, Q => LMD_reg_7_port, QN => n_2296);
   LMD_reg_reg_8_inst : DFFR_X1 port map( D => mem_out_8_port, CK => CLK, RN =>
                           n8, Q => LMD_reg_8_port, QN => n_2297);
   LMD_reg_reg_9_inst : DFFR_X1 port map( D => mem_out_9_port, CK => CLK, RN =>
                           n8, Q => LMD_reg_9_port, QN => n_2298);
   LMD_reg_reg_10_inst : DFFR_X1 port map( D => mem_out_10_port, CK => CLK, RN 
                           => n8, Q => LMD_reg_10_port, QN => n_2299);
   LMD_reg_reg_11_inst : DFFR_X1 port map( D => mem_out_11_port, CK => CLK, RN 
                           => n8, Q => LMD_reg_11_port, QN => n_2300);
   LMD_reg_reg_12_inst : DFFR_X1 port map( D => mem_out_12_port, CK => CLK, RN 
                           => n8, Q => LMD_reg_12_port, QN => n_2301);
   LMD_reg_reg_13_inst : DFFR_X1 port map( D => mem_out_13_port, CK => CLK, RN 
                           => n8, Q => LMD_reg_13_port, QN => n_2302);
   LMD_reg_reg_14_inst : DFFR_X1 port map( D => mem_out_14_port, CK => CLK, RN 
                           => n8, Q => LMD_reg_14_port, QN => n_2303);
   LMD_reg_reg_15_inst : DFFR_X1 port map( D => mem_out_15_port, CK => CLK, RN 
                           => n8, Q => LMD_reg_15_port, QN => n_2304);
   LMD_reg_reg_16_inst : DFFR_X1 port map( D => mem_out_16_port, CK => CLK, RN 
                           => n8, Q => LMD_reg_16_port, QN => n_2305);
   LMD_reg_reg_17_inst : DFFR_X1 port map( D => mem_out_17_port, CK => CLK, RN 
                           => n8, Q => LMD_reg_17_port, QN => n_2306);
   LMD_reg_reg_18_inst : DFFR_X1 port map( D => mem_out_18_port, CK => CLK, RN 
                           => n8, Q => LMD_reg_18_port, QN => n_2307);
   LMD_reg_reg_19_inst : DFFR_X1 port map( D => mem_out_19_port, CK => CLK, RN 
                           => n8, Q => LMD_reg_19_port, QN => n_2308);
   LMD_reg_reg_20_inst : DFFR_X1 port map( D => mem_out_20_port, CK => CLK, RN 
                           => n8, Q => LMD_reg_20_port, QN => n_2309);
   LMD_reg_reg_21_inst : DFFR_X1 port map( D => mem_out_21_port, CK => CLK, RN 
                           => n8, Q => LMD_reg_21_port, QN => n_2310);
   LMD_reg_reg_22_inst : DFFR_X1 port map( D => mem_out_22_port, CK => CLK, RN 
                           => n8, Q => LMD_reg_22_port, QN => n_2311);
   LMD_reg_reg_23_inst : DFFR_X1 port map( D => mem_out_23_port, CK => CLK, RN 
                           => n8, Q => LMD_reg_23_port, QN => n_2312);
   LMD_reg_reg_24_inst : DFFR_X1 port map( D => mem_out_24_port, CK => CLK, RN 
                           => n8, Q => LMD_reg_24_port, QN => n_2313);
   LMD_reg_reg_25_inst : DFFR_X1 port map( D => mem_out_25_port, CK => CLK, RN 
                           => n8, Q => LMD_reg_25_port, QN => n_2314);
   LMD_reg_reg_26_inst : DFFR_X1 port map( D => mem_out_26_port, CK => CLK, RN 
                           => n8, Q => LMD_reg_26_port, QN => n_2315);
   LMD_reg_reg_27_inst : DFFR_X1 port map( D => mem_out_27_port, CK => CLK, RN 
                           => n8, Q => LMD_reg_27_port, QN => n_2316);
   LMD_reg_reg_28_inst : DFFR_X1 port map( D => mem_out_28_port, CK => CLK, RN 
                           => n8, Q => LMD_reg_28_port, QN => n_2317);
   LMD_reg_reg_29_inst : DFFR_X1 port map( D => mem_out_29_port, CK => CLK, RN 
                           => n8, Q => LMD_reg_29_port, QN => n_2318);
   LMD_reg_reg_30_inst : DFFR_X1 port map( D => mem_out_30_port, CK => CLK, RN 
                           => n8, Q => LMD_reg_30_port, QN => n_2319);
   LMD_reg_reg_31_inst : DFFR_X1 port map( D => mem_out_31_port, CK => CLK, RN 
                           => n8, Q => LMD_reg_31_port, QN => n_2320);
   MUX : MUX21_GENERIC_NBIT32_0 port map( A(31) => NPC_fetchout_31_port, A(30) 
                           => NPC_fetchout_30_port, A(29) => 
                           NPC_fetchout_29_port, A(28) => NPC_fetchout_28_port,
                           A(27) => NPC_fetchout_27_port, A(26) => 
                           NPC_fetchout_26_port, A(25) => NPC_fetchout_25_port,
                           A(24) => NPC_fetchout_24_port, A(23) => 
                           NPC_fetchout_23_port, A(22) => NPC_fetchout_22_port,
                           A(21) => NPC_fetchout_21_port, A(20) => 
                           NPC_fetchout_20_port, A(19) => NPC_fetchout_19_port,
                           A(18) => NPC_fetchout_18_port, A(17) => 
                           NPC_fetchout_17_port, A(16) => NPC_fetchout_16_port,
                           A(15) => NPC_fetchout_15_port, A(14) => 
                           NPC_fetchout_14_port, A(13) => NPC_fetchout_13_port,
                           A(12) => NPC_fetchout_12_port, A(11) => 
                           NPC_fetchout_11_port, A(10) => NPC_fetchout_10_port,
                           A(9) => NPC_fetchout_9_port, A(8) => 
                           NPC_fetchout_8_port, A(7) => NPC_fetchout_7_port, 
                           A(6) => NPC_fetchout_6_port, A(5) => 
                           NPC_fetchout_5_port, A(4) => NPC_fetchout_4_port, 
                           A(3) => NPC_fetchout_3_port, A(2) => 
                           NPC_fetchout_2_port, A(1) => NPC_fetchout_1_port, 
                           A(0) => NPC_fetchout_0_port, B(31) => 
                           s_NPC_jump_31_port, B(30) => s_NPC_jump_30_port, 
                           B(29) => s_NPC_jump_29_port, B(28) => 
                           s_NPC_jump_28_port, B(27) => s_NPC_jump_27_port, 
                           B(26) => s_NPC_jump_26_port, B(25) => 
                           s_NPC_jump_25_port, B(24) => s_NPC_jump_24_port, 
                           B(23) => s_NPC_jump_23_port, B(22) => 
                           s_NPC_jump_22_port, B(21) => s_NPC_jump_21_port, 
                           B(20) => s_NPC_jump_20_port, B(19) => 
                           s_NPC_jump_19_port, B(18) => s_NPC_jump_18_port, 
                           B(17) => s_NPC_jump_17_port, B(16) => 
                           s_NPC_jump_16_port, B(15) => s_NPC_jump_15_port, 
                           B(14) => s_NPC_jump_14_port, B(13) => 
                           s_NPC_jump_13_port, B(12) => s_NPC_jump_12_port, 
                           B(11) => s_NPC_jump_11_port, B(10) => 
                           s_NPC_jump_10_port, B(9) => s_NPC_jump_9_port, B(8) 
                           => s_NPC_jump_8_port, B(7) => s_NPC_jump_7_port, 
                           B(6) => s_NPC_jump_6_port, B(5) => s_NPC_jump_5_port
                           , B(4) => s_NPC_jump_4_port, B(3) => 
                           s_NPC_jump_3_port, B(2) => s_NPC_jump_2_port, B(1) 
                           => s_NPC_jump_1_port, B(0) => s_NPC_jump_0_port, SEL
                           => flag_signal, Y(31) => PC_muxout_31_port, Y(30) =>
                           PC_muxout_30_port, Y(29) => PC_muxout_29_port, Y(28)
                           => PC_muxout_28_port, Y(27) => PC_muxout_27_port, 
                           Y(26) => PC_muxout_26_port, Y(25) => 
                           PC_muxout_25_port, Y(24) => PC_muxout_24_port, Y(23)
                           => PC_muxout_23_port, Y(22) => PC_muxout_22_port, 
                           Y(21) => PC_muxout_21_port, Y(20) => 
                           PC_muxout_20_port, Y(19) => PC_muxout_19_port, Y(18)
                           => PC_muxout_18_port, Y(17) => PC_muxout_17_port, 
                           Y(16) => PC_muxout_16_port, Y(15) => 
                           PC_muxout_15_port, Y(14) => PC_muxout_14_port, Y(13)
                           => PC_muxout_13_port, Y(12) => PC_muxout_12_port, 
                           Y(11) => PC_muxout_11_port, Y(10) => 
                           PC_muxout_10_port, Y(9) => PC_muxout_9_port, Y(8) =>
                           PC_muxout_8_port, Y(7) => PC_muxout_7_port, Y(6) => 
                           PC_muxout_6_port, Y(5) => PC_muxout_5_port, Y(4) => 
                           PC_muxout_4_port, Y(3) => PC_muxout_3_port, Y(2) => 
                           PC_muxout_2_port, Y(1) => PC_muxout_1_port, Y(0) => 
                           PC_muxout_0_port);
   fetch_stage : FETCH port map( PC(31) => PC_reg_31_port, PC(30) => 
                           PC_reg_30_port, PC(29) => PC_reg_29_port, PC(28) => 
                           PC_reg_28_port, PC(27) => PC_reg_27_port, PC(26) => 
                           PC_reg_26_port, PC(25) => PC_reg_25_port, PC(24) => 
                           PC_reg_24_port, PC(23) => PC_reg_23_port, PC(22) => 
                           PC_reg_22_port, PC(21) => PC_reg_21_port, PC(20) => 
                           PC_reg_20_port, PC(19) => PC_reg_19_port, PC(18) => 
                           PC_reg_18_port, PC(17) => PC_reg_17_port, PC(16) => 
                           PC_reg_16_port, PC(15) => PC_reg_15_port, PC(14) => 
                           PC_reg_14_port, PC(13) => PC_reg_13_port, PC(12) => 
                           PC_reg_12_port, PC(11) => PC_reg_11_port, PC(10) => 
                           PC_reg_10_port, PC(9) => PC_reg_9_port, PC(8) => 
                           PC_reg_8_port, PC(7) => PC_reg_7_port, PC(6) => 
                           PC_reg_6_port, PC(5) => PC_reg_5_port, PC(4) => 
                           PC_reg_4_port, PC(3) => PC_reg_3_port, PC(2) => 
                           PC_reg_2_port, PC(1) => PC_reg_1_port, PC(0) => 
                           PC_reg_0_port, hazard_PC(31) => hazard_NPC_31_port, 
                           hazard_PC(30) => hazard_NPC_30_port, hazard_PC(29) 
                           => hazard_NPC_29_port, hazard_PC(28) => 
                           hazard_NPC_28_port, hazard_PC(27) => 
                           hazard_NPC_27_port, hazard_PC(26) => 
                           hazard_NPC_26_port, hazard_PC(25) => 
                           hazard_NPC_25_port, hazard_PC(24) => 
                           hazard_NPC_24_port, hazard_PC(23) => 
                           hazard_NPC_23_port, hazard_PC(22) => 
                           hazard_NPC_22_port, hazard_PC(21) => 
                           hazard_NPC_21_port, hazard_PC(20) => 
                           hazard_NPC_20_port, hazard_PC(19) => 
                           hazard_NPC_19_port, hazard_PC(18) => 
                           hazard_NPC_18_port, hazard_PC(17) => 
                           hazard_NPC_17_port, hazard_PC(16) => 
                           hazard_NPC_16_port, hazard_PC(15) => 
                           hazard_NPC_15_port, hazard_PC(14) => 
                           hazard_NPC_14_port, hazard_PC(13) => 
                           hazard_NPC_13_port, hazard_PC(12) => 
                           hazard_NPC_12_port, hazard_PC(11) => 
                           hazard_NPC_11_port, hazard_PC(10) => 
                           hazard_NPC_10_port, hazard_PC(9) => 
                           hazard_NPC_9_port, hazard_PC(8) => hazard_NPC_8_port
                           , hazard_PC(7) => hazard_NPC_7_port, hazard_PC(6) =>
                           hazard_NPC_6_port, hazard_PC(5) => hazard_NPC_5_port
                           , hazard_PC(4) => hazard_NPC_4_port, hazard_PC(3) =>
                           hazard_NPC_3_port, hazard_PC(2) => hazard_NPC_2_port
                           , hazard_PC(1) => hazard_NPC_1_port, hazard_PC(0) =>
                           hazard_NPC_0_port, PC_sel => hazard_NPC_sel, 
                           IRAM_addr(31) => IRAM_addr(31), IRAM_addr(30) => 
                           IRAM_addr(30), IRAM_addr(29) => IRAM_addr(29), 
                           IRAM_addr(28) => IRAM_addr(28), IRAM_addr(27) => 
                           IRAM_addr(27), IRAM_addr(26) => IRAM_addr(26), 
                           IRAM_addr(25) => IRAM_addr(25), IRAM_addr(24) => 
                           IRAM_addr(24), IRAM_addr(23) => IRAM_addr(23), 
                           IRAM_addr(22) => IRAM_addr(22), IRAM_addr(21) => 
                           IRAM_addr(21), IRAM_addr(20) => IRAM_addr(20), 
                           IRAM_addr(19) => IRAM_addr(19), IRAM_addr(18) => 
                           IRAM_addr(18), IRAM_addr(17) => IRAM_addr(17), 
                           IRAM_addr(16) => IRAM_addr(16), IRAM_addr(15) => 
                           IRAM_addr(15), IRAM_addr(14) => IRAM_addr(14), 
                           IRAM_addr(13) => IRAM_addr(13), IRAM_addr(12) => 
                           IRAM_addr(12), IRAM_addr(11) => IRAM_addr(11), 
                           IRAM_addr(10) => IRAM_addr(10), IRAM_addr(9) => 
                           IRAM_addr(9), IRAM_addr(8) => IRAM_addr(8), 
                           IRAM_addr(7) => IRAM_addr(7), IRAM_addr(6) => 
                           IRAM_addr(6), IRAM_addr(5) => IRAM_addr(5), 
                           IRAM_addr(4) => IRAM_addr(4), IRAM_addr(3) => 
                           IRAM_addr(3), IRAM_addr(2) => IRAM_addr(2), 
                           IRAM_addr(1) => IRAM_addr(1), IRAM_addr(0) => 
                           IRAM_addr(0), NPC(31) => NPC_fetchout_31_port, 
                           NPC(30) => NPC_fetchout_30_port, NPC(29) => 
                           NPC_fetchout_29_port, NPC(28) => 
                           NPC_fetchout_28_port, NPC(27) => 
                           NPC_fetchout_27_port, NPC(26) => 
                           NPC_fetchout_26_port, NPC(25) => 
                           NPC_fetchout_25_port, NPC(24) => 
                           NPC_fetchout_24_port, NPC(23) => 
                           NPC_fetchout_23_port, NPC(22) => 
                           NPC_fetchout_22_port, NPC(21) => 
                           NPC_fetchout_21_port, NPC(20) => 
                           NPC_fetchout_20_port, NPC(19) => 
                           NPC_fetchout_19_port, NPC(18) => 
                           NPC_fetchout_18_port, NPC(17) => 
                           NPC_fetchout_17_port, NPC(16) => 
                           NPC_fetchout_16_port, NPC(15) => 
                           NPC_fetchout_15_port, NPC(14) => 
                           NPC_fetchout_14_port, NPC(13) => 
                           NPC_fetchout_13_port, NPC(12) => 
                           NPC_fetchout_12_port, NPC(11) => 
                           NPC_fetchout_11_port, NPC(10) => 
                           NPC_fetchout_10_port, NPC(9) => NPC_fetchout_9_port,
                           NPC(8) => NPC_fetchout_8_port, NPC(7) => 
                           NPC_fetchout_7_port, NPC(6) => NPC_fetchout_6_port, 
                           NPC(5) => NPC_fetchout_5_port, NPC(4) => 
                           NPC_fetchout_4_port, NPC(3) => NPC_fetchout_3_port, 
                           NPC(2) => NPC_fetchout_2_port, NPC(1) => 
                           NPC_fetchout_1_port, NPC(0) => NPC_fetchout_0_port);
   NOP_MUX : MUX21_GENERIC_NBIT32_5 port map( A(31) => instr(31), A(30) => 
                           instr(30), A(29) => instr(29), A(28) => instr(28), 
                           A(27) => instr(27), A(26) => instr(26), A(25) => 
                           instr(25), A(24) => instr(24), A(23) => instr(23), 
                           A(22) => instr(22), A(21) => instr(21), A(20) => 
                           instr(20), A(19) => instr(19), A(18) => instr(18), 
                           A(17) => instr(17), A(16) => instr(16), A(15) => 
                           instr(15), A(14) => instr(14), A(13) => instr(13), 
                           A(12) => instr(12), A(11) => instr(11), A(10) => 
                           instr(10), A(9) => instr(9), A(8) => instr(8), A(7) 
                           => instr(7), A(6) => instr(6), A(5) => instr(5), 
                           A(4) => instr(4), A(3) => instr(3), A(2) => instr(2)
                           , A(1) => instr(1), A(0) => instr(0), B(31) => 
                           X_Logic0_port, B(30) => X_Logic1_port, B(29) => 
                           X_Logic0_port, B(28) => X_Logic1_port, B(27) => 
                           X_Logic0_port, B(26) => X_Logic1_port, B(25) => 
                           X_Logic0_port, B(24) => X_Logic0_port, B(23) => 
                           X_Logic0_port, B(22) => X_Logic0_port, B(21) => 
                           X_Logic0_port, B(20) => X_Logic0_port, B(19) => 
                           X_Logic0_port, B(18) => X_Logic0_port, B(17) => 
                           X_Logic0_port, B(16) => X_Logic0_port, B(15) => 
                           X_Logic0_port, B(14) => X_Logic0_port, B(13) => 
                           X_Logic0_port, B(12) => X_Logic0_port, B(11) => 
                           X_Logic0_port, B(10) => X_Logic0_port, B(9) => 
                           X_Logic0_port, B(8) => X_Logic0_port, B(7) => 
                           X_Logic0_port, B(6) => X_Logic0_port, B(5) => 
                           X_Logic0_port, B(4) => X_Logic0_port, B(3) => 
                           X_Logic0_port, B(2) => X_Logic0_port, B(1) => 
                           X_Logic0_port, B(0) => X_Logic0_port, SEL => 
                           flag_signal, Y(31) => NOP_MUX_OUT_31_port, Y(30) => 
                           NOP_MUX_OUT_30_port, Y(29) => NOP_MUX_OUT_29_port, 
                           Y(28) => NOP_MUX_OUT_28_port, Y(27) => 
                           NOP_MUX_OUT_27_port, Y(26) => NOP_MUX_OUT_26_port, 
                           Y(25) => NOP_MUX_OUT_25_port, Y(24) => 
                           NOP_MUX_OUT_24_port, Y(23) => NOP_MUX_OUT_23_port, 
                           Y(22) => NOP_MUX_OUT_22_port, Y(21) => 
                           NOP_MUX_OUT_21_port, Y(20) => NOP_MUX_OUT_20_port, 
                           Y(19) => NOP_MUX_OUT_19_port, Y(18) => 
                           NOP_MUX_OUT_18_port, Y(17) => NOP_MUX_OUT_17_port, 
                           Y(16) => NOP_MUX_OUT_16_port, Y(15) => 
                           NOP_MUX_OUT_15_port, Y(14) => NOP_MUX_OUT_14_port, 
                           Y(13) => NOP_MUX_OUT_13_port, Y(12) => 
                           NOP_MUX_OUT_12_port, Y(11) => NOP_MUX_OUT_11_port, 
                           Y(10) => NOP_MUX_OUT_10_port, Y(9) => 
                           NOP_MUX_OUT_9_port, Y(8) => NOP_MUX_OUT_8_port, Y(7)
                           => NOP_MUX_OUT_7_port, Y(6) => NOP_MUX_OUT_6_port, 
                           Y(5) => NOP_MUX_OUT_5_port, Y(4) => 
                           NOP_MUX_OUT_4_port, Y(3) => NOP_MUX_OUT_3_port, Y(2)
                           => NOP_MUX_OUT_2_port, Y(1) => NOP_MUX_OUT_1_port, 
                           Y(0) => NOP_MUX_OUT_0_port);
   dec_stage : DEC port map( instr(31) => IR_reg_31_port, instr(30) => 
                           IR_reg_30_port, instr(29) => IR_reg_29_port, 
                           instr(28) => IR_reg_28_port, instr(27) => 
                           IR_reg_27_port, instr(26) => IR_reg_26_port, 
                           instr(25) => IR_reg_25_port, instr(24) => 
                           IR_reg_24_port, instr(23) => IR_reg_23_port, 
                           instr(22) => IR_reg_22_port, instr(21) => 
                           IR_reg_21_port, instr(20) => IR_reg_20_port, 
                           instr(19) => IR_reg_19_port, instr(18) => 
                           IR_reg_18_port, instr(17) => IR_reg_17_port, 
                           instr(16) => IR_reg_16_port, instr(15) => 
                           IR_reg_15_port, instr(14) => IR_reg_14_port, 
                           instr(13) => IR_reg_13_port, instr(12) => 
                           IR_reg_12_port, instr(11) => IR_reg_11_port, 
                           instr(10) => IR_reg_10_port, instr(9) => 
                           IR_reg_9_port, instr(8) => IR_reg_8_port, instr(7) 
                           => IR_reg_7_port, instr(6) => IR_reg_6_port, 
                           instr(5) => IR_reg_5_port, instr(4) => IR_reg_4_port
                           , instr(3) => IR_reg_3_port, instr(2) => 
                           IR_reg_2_port, instr(1) => IR_reg_1_port, instr(0) 
                           => IR_reg_0_port, RST => n4, RFdata_in(31) => 
                           WB_data_31_port, RFdata_in(30) => WB_data_30_port, 
                           RFdata_in(29) => WB_data_29_port, RFdata_in(28) => 
                           WB_data_28_port, RFdata_in(27) => WB_data_27_port, 
                           RFdata_in(26) => WB_data_26_port, RFdata_in(25) => 
                           WB_data_25_port, RFdata_in(24) => WB_data_24_port, 
                           RFdata_in(23) => WB_data_23_port, RFdata_in(22) => 
                           WB_data_22_port, RFdata_in(21) => WB_data_21_port, 
                           RFdata_in(20) => WB_data_20_port, RFdata_in(19) => 
                           WB_data_19_port, RFdata_in(18) => WB_data_18_port, 
                           RFdata_in(17) => WB_data_17_port, RFdata_in(16) => 
                           WB_data_16_port, RFdata_in(15) => WB_data_15_port, 
                           RFdata_in(14) => WB_data_14_port, RFdata_in(13) => 
                           WB_data_13_port, RFdata_in(12) => WB_data_12_port, 
                           RFdata_in(11) => WB_data_11_port, RFdata_in(10) => 
                           WB_data_10_port, RFdata_in(9) => WB_data_9_port, 
                           RFdata_in(8) => WB_data_8_port, RFdata_in(7) => 
                           WB_data_7_port, RFdata_in(6) => WB_data_6_port, 
                           RFdata_in(5) => WB_data_5_port, RFdata_in(4) => 
                           WB_data_4_port, RFdata_in(3) => WB_data_3_port, 
                           RFdata_in(2) => WB_data_2_port, RFdata_in(1) => 
                           WB_data_1_port, RFdata_in(0) => WB_data_0_port, 
                           RFWA(4) => RD_regwb_4_port, RFWA(3) => 
                           RD_regwb_3_port, RFWA(2) => RD_regwb_2_port, RFWA(1)
                           => RD_regwb_1_port, RFWA(0) => RD_regwb_0_port, 
                           NPC_in(31) => NPC_reg_31_port, NPC_in(30) => 
                           NPC_reg_30_port, NPC_in(29) => NPC_reg_29_port, 
                           NPC_in(28) => NPC_reg_28_port, NPC_in(27) => 
                           NPC_reg_27_port, NPC_in(26) => NPC_reg_26_port, 
                           NPC_in(25) => NPC_reg_25_port, NPC_in(24) => 
                           NPC_reg_24_port, NPC_in(23) => NPC_reg_23_port, 
                           NPC_in(22) => NPC_reg_22_port, NPC_in(21) => 
                           NPC_reg_21_port, NPC_in(20) => NPC_reg_20_port, 
                           NPC_in(19) => NPC_reg_19_port, NPC_in(18) => 
                           NPC_reg_18_port, NPC_in(17) => NPC_reg_17_port, 
                           NPC_in(16) => NPC_reg_16_port, NPC_in(15) => 
                           NPC_reg_15_port, NPC_in(14) => NPC_reg_14_port, 
                           NPC_in(13) => NPC_reg_13_port, NPC_in(12) => 
                           NPC_reg_12_port, NPC_in(11) => NPC_reg_11_port, 
                           NPC_in(10) => NPC_reg_10_port, NPC_in(9) => 
                           NPC_reg_9_port, NPC_in(8) => NPC_reg_8_port, 
                           NPC_in(7) => NPC_reg_7_port, NPC_in(6) => 
                           NPC_reg_6_port, NPC_in(5) => NPC_reg_5_port, 
                           NPC_in(4) => NPC_reg_4_port, NPC_in(3) => 
                           NPC_reg_3_port, NPC_in(2) => NPC_reg_2_port, 
                           NPC_in(1) => NPC_reg_1_port, NPC_in(0) => 
                           NPC_reg_0_port, EXE_RD(4) => RD_regexe_4_port, 
                           EXE_RD(3) => RD_regexe_3_port, EXE_RD(2) => 
                           RD_regexe_2_port, EXE_RD(1) => RD_regexe_1_port, 
                           EXE_RD(0) => RD_regexe_0_port, Ld => Ld, 
                           ALU_regout(31) => ALU_reg_31_port, ALU_regout(30) =>
                           ALU_reg_30_port, ALU_regout(29) => ALU_reg_29_port, 
                           ALU_regout(28) => ALU_reg_28_port, ALU_regout(27) =>
                           ALU_reg_27_port, ALU_regout(26) => ALU_reg_26_port, 
                           ALU_regout(25) => ALU_reg_25_port, ALU_regout(24) =>
                           ALU_reg_24_port, ALU_regout(23) => ALU_reg_23_port, 
                           ALU_regout(22) => ALU_reg_22_port, ALU_regout(21) =>
                           ALU_reg_21_port, ALU_regout(20) => ALU_reg_20_port, 
                           ALU_regout(19) => ALU_reg_19_port, ALU_regout(18) =>
                           ALU_reg_18_port, ALU_regout(17) => ALU_reg_17_port, 
                           ALU_regout(16) => ALU_reg_16_port, ALU_regout(15) =>
                           ALU_reg_15_port, ALU_regout(14) => ALU_reg_14_port, 
                           ALU_regout(13) => ALU_reg_13_port, ALU_regout(12) =>
                           ALU_reg_12_port, ALU_regout(11) => ALU_reg_11_port, 
                           ALU_regout(10) => ALU_reg_10_port, ALU_regout(9) => 
                           ALU_reg_9_port, ALU_regout(8) => ALU_reg_8_port, 
                           ALU_regout(7) => ALU_reg_7_port, ALU_regout(6) => 
                           ALU_reg_6_port, ALU_regout(5) => ALU_reg_5_port, 
                           ALU_regout(4) => ALU_reg_4_port, ALU_regout(3) => 
                           ALU_reg_3_port, ALU_regout(2) => ALU_reg_2_port, 
                           ALU_regout(1) => ALU_reg_1_port, ALU_regout(0) => 
                           ALU_reg_0_port, MEM_RD(4) => RD_regmem_4_port, 
                           MEM_RD(3) => RD_regmem_3_port, MEM_RD(2) => 
                           RD_regmem_2_port, MEM_RD(1) => RD_regmem_1_port, 
                           MEM_RD(0) => RD_regmem_0_port, WB_RD(4) => 
                           RD_regwb_4_port, WB_RD(3) => RD_regwb_3_port, 
                           WB_RD(2) => RD_regwb_2_port, WB_RD(1) => 
                           RD_regwb_1_port, WB_RD(0) => RD_regwb_0_port, 
                           RD_inmul(4) => s_RD_inmul_4_port, RD_inmul(3) => 
                           s_RD_inmul_3_port, RD_inmul(2) => s_RD_inmul_2_port,
                           RD_inmul(1) => s_RD_inmul_1_port, RD_inmul(0) => 
                           s_RD_inmul_0_port, flag_structHzd => 
                           s_flag_structHzd, flag_ismul => s_flag_ismul, RF1 =>
                           RF1, RF2 => RF2, WF1 => WF1, EN1 => EN1, opcode(5) 
                           => opcode(5), opcode(4) => opcode(4), opcode(3) => 
                           opcode(3), opcode(2) => opcode(2), opcode(1) => 
                           opcode(1), opcode(0) => opcode(0), func(10) => 
                           func(10), func(9) => func(9), func(8) => func(8), 
                           func(7) => func(7), func(6) => func(6), func(5) => 
                           func(5), func(4) => func(4), func(3) => func(3), 
                           func(2) => func(2), func(1) => func(1), func(0) => 
                           func(0), IMM(31) => IMM_decout_31_port, IMM(30) => 
                           IMM_decout_30_port, IMM(29) => IMM_decout_29_port, 
                           IMM(28) => IMM_decout_28_port, IMM(27) => 
                           IMM_decout_27_port, IMM(26) => IMM_decout_26_port, 
                           IMM(25) => IMM_decout_25_port, IMM(24) => 
                           IMM_decout_24_port, IMM(23) => IMM_decout_23_port, 
                           IMM(22) => IMM_decout_22_port, IMM(21) => 
                           IMM_decout_21_port, IMM(20) => IMM_decout_20_port, 
                           IMM(19) => IMM_decout_19_port, IMM(18) => 
                           IMM_decout_18_port, IMM(17) => IMM_decout_17_port, 
                           IMM(16) => IMM_decout_16_port, IMM(15) => 
                           IMM_decout_15_port, IMM(14) => IMM_decout_14_port, 
                           IMM(13) => IMM_decout_13_port, IMM(12) => 
                           IMM_decout_12_port, IMM(11) => IMM_decout_11_port, 
                           IMM(10) => IMM_decout_10_port, IMM(9) => 
                           IMM_decout_9_port, IMM(8) => IMM_decout_8_port, 
                           IMM(7) => IMM_decout_7_port, IMM(6) => 
                           IMM_decout_6_port, IMM(5) => IMM_decout_5_port, 
                           IMM(4) => IMM_decout_4_port, IMM(3) => 
                           IMM_decout_3_port, IMM(2) => IMM_decout_2_port, 
                           IMM(1) => IMM_decout_1_port, IMM(0) => 
                           IMM_decout_0_port, RA(31) => RA_decout_31_port, 
                           RA(30) => RA_decout_30_port, RA(29) => 
                           RA_decout_29_port, RA(28) => RA_decout_28_port, 
                           RA(27) => RA_decout_27_port, RA(26) => 
                           RA_decout_26_port, RA(25) => RA_decout_25_port, 
                           RA(24) => RA_decout_24_port, RA(23) => 
                           RA_decout_23_port, RA(22) => RA_decout_22_port, 
                           RA(21) => RA_decout_21_port, RA(20) => 
                           RA_decout_20_port, RA(19) => RA_decout_19_port, 
                           RA(18) => RA_decout_18_port, RA(17) => 
                           RA_decout_17_port, RA(16) => RA_decout_16_port, 
                           RA(15) => RA_decout_15_port, RA(14) => 
                           RA_decout_14_port, RA(13) => RA_decout_13_port, 
                           RA(12) => RA_decout_12_port, RA(11) => 
                           RA_decout_11_port, RA(10) => RA_decout_10_port, 
                           RA(9) => RA_decout_9_port, RA(8) => RA_decout_8_port
                           , RA(7) => RA_decout_7_port, RA(6) => 
                           RA_decout_6_port, RA(5) => RA_decout_5_port, RA(4) 
                           => RA_decout_4_port, RA(3) => RA_decout_3_port, 
                           RA(2) => RA_decout_2_port, RA(1) => RA_decout_1_port
                           , RA(0) => RA_decout_0_port, RB(31) => 
                           RB_decout_31_port, RB(30) => RB_decout_30_port, 
                           RB(29) => RB_decout_29_port, RB(28) => 
                           RB_decout_28_port, RB(27) => RB_decout_27_port, 
                           RB(26) => RB_decout_26_port, RB(25) => 
                           RB_decout_25_port, RB(24) => RB_decout_24_port, 
                           RB(23) => RB_decout_23_port, RB(22) => 
                           RB_decout_22_port, RB(21) => RB_decout_21_port, 
                           RB(20) => RB_decout_20_port, RB(19) => 
                           RB_decout_19_port, RB(18) => RB_decout_18_port, 
                           RB(17) => RB_decout_17_port, RB(16) => 
                           RB_decout_16_port, RB(15) => RB_decout_15_port, 
                           RB(14) => RB_decout_14_port, RB(13) => 
                           RB_decout_13_port, RB(12) => RB_decout_12_port, 
                           RB(11) => RB_decout_11_port, RB(10) => 
                           RB_decout_10_port, RB(9) => RB_decout_9_port, RB(8) 
                           => RB_decout_8_port, RB(7) => RB_decout_7_port, 
                           RB(6) => RB_decout_6_port, RB(5) => RB_decout_5_port
                           , RB(4) => RB_decout_4_port, RB(3) => 
                           RB_decout_3_port, RB(2) => RB_decout_2_port, RB(1) 
                           => RB_decout_1_port, RB(0) => RB_decout_0_port, 
                           RSA(4) => RSA_decout_4_port, RSA(3) => 
                           RSA_decout_3_port, RSA(2) => RSA_decout_2_port, 
                           RSA(1) => RSA_decout_1_port, RSA(0) => 
                           RSA_decout_0_port, RSB(4) => RSB_decout_4_port, 
                           RSB(3) => RSB_decout_3_port, RSB(2) => 
                           RSB_decout_2_port, RSB(1) => RSB_decout_1_port, 
                           RSB(0) => RSB_decout_0_port, RD(4) => 
                           RD_decout_4_port, RD(3) => RD_decout_3_port, RD(2) 
                           => RD_decout_2_port, RD(1) => RD_decout_1_port, 
                           RD(0) => RD_decout_0_port, stall_NPC(31) => 
                           hazard_NPC_31_port, stall_NPC(30) => 
                           hazard_NPC_30_port, stall_NPC(29) => 
                           hazard_NPC_29_port, stall_NPC(28) => 
                           hazard_NPC_28_port, stall_NPC(27) => 
                           hazard_NPC_27_port, stall_NPC(26) => 
                           hazard_NPC_26_port, stall_NPC(25) => 
                           hazard_NPC_25_port, stall_NPC(24) => 
                           hazard_NPC_24_port, stall_NPC(23) => 
                           hazard_NPC_23_port, stall_NPC(22) => 
                           hazard_NPC_22_port, stall_NPC(21) => 
                           hazard_NPC_21_port, stall_NPC(20) => 
                           hazard_NPC_20_port, stall_NPC(19) => 
                           hazard_NPC_19_port, stall_NPC(18) => 
                           hazard_NPC_18_port, stall_NPC(17) => 
                           hazard_NPC_17_port, stall_NPC(16) => 
                           hazard_NPC_16_port, stall_NPC(15) => 
                           hazard_NPC_15_port, stall_NPC(14) => 
                           hazard_NPC_14_port, stall_NPC(13) => 
                           hazard_NPC_13_port, stall_NPC(12) => 
                           hazard_NPC_12_port, stall_NPC(11) => 
                           hazard_NPC_11_port, stall_NPC(10) => 
                           hazard_NPC_10_port, stall_NPC(9) => 
                           hazard_NPC_9_port, stall_NPC(8) => hazard_NPC_8_port
                           , stall_NPC(7) => hazard_NPC_7_port, stall_NPC(6) =>
                           hazard_NPC_6_port, stall_NPC(5) => hazard_NPC_5_port
                           , stall_NPC(4) => hazard_NPC_4_port, stall_NPC(3) =>
                           hazard_NPC_3_port, stall_NPC(2) => hazard_NPC_2_port
                           , stall_NPC(1) => hazard_NPC_1_port, stall_NPC(0) =>
                           hazard_NPC_0_port, PC_sel => hazard_NPC_sel, 
                           dec_flag => flag_signal, NPC_jump(31) => 
                           s_NPC_jump_31_port, NPC_jump(30) => 
                           s_NPC_jump_30_port, NPC_jump(29) => 
                           s_NPC_jump_29_port, NPC_jump(28) => 
                           s_NPC_jump_28_port, NPC_jump(27) => 
                           s_NPC_jump_27_port, NPC_jump(26) => 
                           s_NPC_jump_26_port, NPC_jump(25) => 
                           s_NPC_jump_25_port, NPC_jump(24) => 
                           s_NPC_jump_24_port, NPC_jump(23) => 
                           s_NPC_jump_23_port, NPC_jump(22) => 
                           s_NPC_jump_22_port, NPC_jump(21) => 
                           s_NPC_jump_21_port, NPC_jump(20) => 
                           s_NPC_jump_20_port, NPC_jump(19) => 
                           s_NPC_jump_19_port, NPC_jump(18) => 
                           s_NPC_jump_18_port, NPC_jump(17) => 
                           s_NPC_jump_17_port, NPC_jump(16) => 
                           s_NPC_jump_16_port, NPC_jump(15) => 
                           s_NPC_jump_15_port, NPC_jump(14) => 
                           s_NPC_jump_14_port, NPC_jump(13) => 
                           s_NPC_jump_13_port, NPC_jump(12) => 
                           s_NPC_jump_12_port, NPC_jump(11) => 
                           s_NPC_jump_11_port, NPC_jump(10) => 
                           s_NPC_jump_10_port, NPC_jump(9) => s_NPC_jump_9_port
                           , NPC_jump(8) => s_NPC_jump_8_port, NPC_jump(7) => 
                           s_NPC_jump_7_port, NPC_jump(6) => s_NPC_jump_6_port,
                           NPC_jump(5) => s_NPC_jump_5_port, NPC_jump(4) => 
                           s_NPC_jump_4_port, NPC_jump(3) => s_NPC_jump_3_port,
                           NPC_jump(2) => s_NPC_jump_2_port, NPC_jump(1) => 
                           s_NPC_jump_1_port, NPC_jump(0) => s_NPC_jump_0_port)
                           ;
   exe_stage : EXE port map( CLK => CLK, RST => n4, IMM(31) => Imm_reg_31_port,
                           IMM(30) => Imm_reg_30_port, IMM(29) => 
                           Imm_reg_29_port, IMM(28) => Imm_reg_28_port, IMM(27)
                           => Imm_reg_27_port, IMM(26) => Imm_reg_26_port, 
                           IMM(25) => Imm_reg_25_port, IMM(24) => 
                           Imm_reg_24_port, IMM(23) => Imm_reg_23_port, IMM(22)
                           => Imm_reg_22_port, IMM(21) => Imm_reg_21_port, 
                           IMM(20) => Imm_reg_20_port, IMM(19) => 
                           Imm_reg_19_port, IMM(18) => Imm_reg_18_port, IMM(17)
                           => Imm_reg_17_port, IMM(16) => Imm_reg_16_port, 
                           IMM(15) => Imm_reg_15_port, IMM(14) => 
                           Imm_reg_14_port, IMM(13) => Imm_reg_13_port, IMM(12)
                           => Imm_reg_12_port, IMM(11) => Imm_reg_11_port, 
                           IMM(10) => Imm_reg_10_port, IMM(9) => Imm_reg_9_port
                           , IMM(8) => Imm_reg_8_port, IMM(7) => Imm_reg_7_port
                           , IMM(6) => Imm_reg_6_port, IMM(5) => Imm_reg_5_port
                           , IMM(4) => Imm_reg_4_port, IMM(3) => Imm_reg_3_port
                           , IMM(2) => Imm_reg_2_port, IMM(1) => Imm_reg_1_port
                           , IMM(0) => Imm_reg_0_port, RA(31) => RA_reg_31_port
                           , RA(30) => RA_reg_30_port, RA(29) => RA_reg_29_port
                           , RA(28) => RA_reg_28_port, RA(27) => RA_reg_27_port
                           , RA(26) => RA_reg_26_port, RA(25) => RA_reg_25_port
                           , RA(24) => RA_reg_24_port, RA(23) => RA_reg_23_port
                           , RA(22) => RA_reg_22_port, RA(21) => RA_reg_21_port
                           , RA(20) => RA_reg_20_port, RA(19) => RA_reg_19_port
                           , RA(18) => RA_reg_18_port, RA(17) => RA_reg_17_port
                           , RA(16) => RA_reg_16_port, RA(15) => RA_reg_15_port
                           , RA(14) => RA_reg_14_port, RA(13) => RA_reg_13_port
                           , RA(12) => RA_reg_12_port, RA(11) => RA_reg_11_port
                           , RA(10) => RA_reg_10_port, RA(9) => RA_reg_9_port, 
                           RA(8) => RA_reg_8_port, RA(7) => RA_reg_7_port, 
                           RA(6) => RA_reg_6_port, RA(5) => RA_reg_5_port, 
                           RA(4) => RA_reg_4_port, RA(3) => RA_reg_3_port, 
                           RA(2) => RA_reg_2_port, RA(1) => RA_reg_1_port, 
                           RA(0) => RA_reg_0_port, RB(31) => RB_reg_31_port, 
                           RB(30) => RB_reg_30_port, RB(29) => RB_reg_29_port, 
                           RB(28) => RB_reg_28_port, RB(27) => RB_reg_27_port, 
                           RB(26) => RB_reg_26_port, RB(25) => RB_reg_25_port, 
                           RB(24) => RB_reg_24_port, RB(23) => RB_reg_23_port, 
                           RB(22) => RB_reg_22_port, RB(21) => RB_reg_21_port, 
                           RB(20) => RB_reg_20_port, RB(19) => RB_reg_19_port, 
                           RB(18) => RB_reg_18_port, RB(17) => RB_reg_17_port, 
                           RB(16) => RB_reg_16_port, RB(15) => RB_reg_15_port, 
                           RB(14) => RB_reg_14_port, RB(13) => RB_reg_13_port, 
                           RB(12) => RB_reg_12_port, RB(11) => RB_reg_11_port, 
                           RB(10) => RB_reg_10_port, RB(9) => RB_reg_9_port, 
                           RB(8) => RB_reg_8_port, RB(7) => RB_reg_7_port, 
                           RB(6) => RB_reg_6_port, RB(5) => RB_reg_5_port, 
                           RB(4) => RB_reg_4_port, RB(3) => RB_reg_3_port, 
                           RB(2) => RB_reg_2_port, RB(1) => RB_reg_1_port, 
                           RB(0) => RB_reg_0_port, WA(4) => RD_regexe_4_port, 
                           WA(3) => RD_regexe_3_port, WA(2) => RD_regexe_2_port
                           , WA(1) => RD_regexe_1_port, WA(0) => 
                           RD_regexe_0_port, RSA(4) => RSA_reg_4_port, RSA(3) 
                           => RSA_reg_3_port, RSA(2) => RSA_reg_2_port, RSA(1) 
                           => RSA_reg_1_port, RSA(0) => RSA_reg_0_port, RSB(4) 
                           => RSB_reg_4_port, RSB(3) => RSB_reg_3_port, RSB(2) 
                           => RSB_reg_2_port, RSB(1) => RSB_reg_1_port, RSB(0) 
                           => RSB_reg_0_port, ALU_outmem(31) => ALU_reg_31_port
                           , ALU_outmem(30) => ALU_reg_30_port, ALU_outmem(29) 
                           => ALU_reg_29_port, ALU_outmem(28) => 
                           ALU_reg_28_port, ALU_outmem(27) => ALU_reg_27_port, 
                           ALU_outmem(26) => ALU_reg_26_port, ALU_outmem(25) =>
                           ALU_reg_25_port, ALU_outmem(24) => ALU_reg_24_port, 
                           ALU_outmem(23) => ALU_reg_23_port, ALU_outmem(22) =>
                           ALU_reg_22_port, ALU_outmem(21) => ALU_reg_21_port, 
                           ALU_outmem(20) => ALU_reg_20_port, ALU_outmem(19) =>
                           ALU_reg_19_port, ALU_outmem(18) => ALU_reg_18_port, 
                           ALU_outmem(17) => ALU_reg_17_port, ALU_outmem(16) =>
                           ALU_reg_16_port, ALU_outmem(15) => ALU_reg_15_port, 
                           ALU_outmem(14) => ALU_reg_14_port, ALU_outmem(13) =>
                           ALU_reg_13_port, ALU_outmem(12) => ALU_reg_12_port, 
                           ALU_outmem(11) => ALU_reg_11_port, ALU_outmem(10) =>
                           ALU_reg_10_port, ALU_outmem(9) => ALU_reg_9_port, 
                           ALU_outmem(8) => ALU_reg_8_port, ALU_outmem(7) => 
                           ALU_reg_7_port, ALU_outmem(6) => ALU_reg_6_port, 
                           ALU_outmem(5) => ALU_reg_5_port, ALU_outmem(4) => 
                           ALU_reg_4_port, ALU_outmem(3) => ALU_reg_3_port, 
                           ALU_outmem(2) => ALU_reg_2_port, ALU_outmem(1) => 
                           ALU_reg_1_port, ALU_outmem(0) => ALU_reg_0_port, 
                           WB_out(31) => WB_data_31_port, WB_out(30) => 
                           WB_data_30_port, WB_out(29) => WB_data_29_port, 
                           WB_out(28) => WB_data_28_port, WB_out(27) => 
                           WB_data_27_port, WB_out(26) => WB_data_26_port, 
                           WB_out(25) => WB_data_25_port, WB_out(24) => 
                           WB_data_24_port, WB_out(23) => WB_data_23_port, 
                           WB_out(22) => WB_data_22_port, WB_out(21) => 
                           WB_data_21_port, WB_out(20) => WB_data_20_port, 
                           WB_out(19) => WB_data_19_port, WB_out(18) => 
                           WB_data_18_port, WB_out(17) => WB_data_17_port, 
                           WB_out(16) => WB_data_16_port, WB_out(15) => 
                           WB_data_15_port, WB_out(14) => WB_data_14_port, 
                           WB_out(13) => WB_data_13_port, WB_out(12) => 
                           WB_data_12_port, WB_out(11) => WB_data_11_port, 
                           WB_out(10) => WB_data_10_port, WB_out(9) => 
                           WB_data_9_port, WB_out(8) => WB_data_8_port, 
                           WB_out(7) => WB_data_7_port, WB_out(6) => 
                           WB_data_6_port, WB_out(5) => WB_data_5_port, 
                           WB_out(4) => WB_data_4_port, WB_out(3) => 
                           WB_data_3_port, WB_out(2) => WB_data_2_port, 
                           WB_out(1) => WB_data_1_port, WB_out(0) => 
                           WB_data_0_port, MEM_RD(4) => RD_regmem_4_port, 
                           MEM_RD(3) => RD_regmem_3_port, MEM_RD(2) => 
                           RD_regmem_2_port, MEM_RD(1) => RD_regmem_1_port, 
                           MEM_RD(0) => RD_regmem_0_port, WB_RD(4) => 
                           RD_regwb_4_port, WB_RD(3) => RD_regwb_3_port, 
                           WB_RD(2) => RD_regwb_2_port, WB_RD(1) => 
                           RD_regwb_1_port, WB_RD(0) => RD_regwb_0_port, LD_EN 
                           => EN3, WB_EN => WF1, S1 => S1, S2 => S2, ALU3 => 
                           ALU3, ALU2 => ALU2, ALU1 => ALU1, ALU0 => ALU0, SN 
                           => SN, RD_inmul(4) => s_RD_inmul_4_port, RD_inmul(3)
                           => s_RD_inmul_3_port, RD_inmul(2) => 
                           s_RD_inmul_2_port, RD_inmul(1) => s_RD_inmul_1_port,
                           RD_inmul(0) => s_RD_inmul_0_port, flag_structHzd => 
                           s_flag_structHzd, flag_ismul => s_flag_ismul, OVF =>
                           OVF, output(31) => ALU_exeout_31_port, output(30) =>
                           ALU_exeout_30_port, output(29) => ALU_exeout_29_port
                           , output(28) => ALU_exeout_28_port, output(27) => 
                           ALU_exeout_27_port, output(26) => ALU_exeout_26_port
                           , output(25) => ALU_exeout_25_port, output(24) => 
                           ALU_exeout_24_port, output(23) => ALU_exeout_23_port
                           , output(22) => ALU_exeout_22_port, output(21) => 
                           ALU_exeout_21_port, output(20) => ALU_exeout_20_port
                           , output(19) => ALU_exeout_19_port, output(18) => 
                           ALU_exeout_18_port, output(17) => ALU_exeout_17_port
                           , output(16) => ALU_exeout_16_port, output(15) => 
                           ALU_exeout_15_port, output(14) => ALU_exeout_14_port
                           , output(13) => ALU_exeout_13_port, output(12) => 
                           ALU_exeout_12_port, output(11) => ALU_exeout_11_port
                           , output(10) => ALU_exeout_10_port, output(9) => 
                           ALU_exeout_9_port, output(8) => ALU_exeout_8_port, 
                           output(7) => ALU_exeout_7_port, output(6) => 
                           ALU_exeout_6_port, output(5) => ALU_exeout_5_port, 
                           output(4) => ALU_exeout_4_port, output(3) => 
                           ALU_exeout_3_port, output(2) => ALU_exeout_2_port, 
                           output(1) => ALU_exeout_1_port, output(0) => 
                           ALU_exeout_0_port, ME(31) => ME_exeout_31_port, 
                           ME(30) => ME_exeout_30_port, ME(29) => 
                           ME_exeout_29_port, ME(28) => ME_exeout_28_port, 
                           ME(27) => ME_exeout_27_port, ME(26) => 
                           ME_exeout_26_port, ME(25) => ME_exeout_25_port, 
                           ME(24) => ME_exeout_24_port, ME(23) => 
                           ME_exeout_23_port, ME(22) => ME_exeout_22_port, 
                           ME(21) => ME_exeout_21_port, ME(20) => 
                           ME_exeout_20_port, ME(19) => ME_exeout_19_port, 
                           ME(18) => ME_exeout_18_port, ME(17) => 
                           ME_exeout_17_port, ME(16) => ME_exeout_16_port, 
                           ME(15) => ME_exeout_15_port, ME(14) => 
                           ME_exeout_14_port, ME(13) => ME_exeout_13_port, 
                           ME(12) => ME_exeout_12_port, ME(11) => 
                           ME_exeout_11_port, ME(10) => ME_exeout_10_port, 
                           ME(9) => ME_exeout_9_port, ME(8) => ME_exeout_8_port
                           , ME(7) => ME_exeout_7_port, ME(6) => 
                           ME_exeout_6_port, ME(5) => ME_exeout_5_port, ME(4) 
                           => ME_exeout_4_port, ME(3) => ME_exeout_3_port, 
                           ME(2) => ME_exeout_2_port, ME(1) => ME_exeout_1_port
                           , ME(0) => ME_exeout_0_port, WAout(4) => 
                           RD_exeout_4_port, WAout(3) => RD_exeout_3_port, 
                           WAout(2) => RD_exeout_2_port, WAout(1) => 
                           RD_exeout_1_port, WAout(0) => RD_exeout_0_port);
   mem_stage : MEM_MEMORY_SIZE128 port map( CLK => CLK, RST => n12, ALUout(31) 
                           => ALU_reg_31_port, ALUout(30) => ALU_reg_30_port, 
                           ALUout(29) => ALU_reg_29_port, ALUout(28) => 
                           ALU_reg_28_port, ALUout(27) => ALU_reg_27_port, 
                           ALUout(26) => ALU_reg_26_port, ALUout(25) => 
                           ALU_reg_25_port, ALUout(24) => ALU_reg_24_port, 
                           ALUout(23) => ALU_reg_23_port, ALUout(22) => 
                           ALU_reg_22_port, ALUout(21) => ALU_reg_21_port, 
                           ALUout(20) => ALU_reg_20_port, ALUout(19) => 
                           ALU_reg_19_port, ALUout(18) => ALU_reg_18_port, 
                           ALUout(17) => ALU_reg_17_port, ALUout(16) => 
                           ALU_reg_16_port, ALUout(15) => ALU_reg_15_port, 
                           ALUout(14) => ALU_reg_14_port, ALUout(13) => 
                           ALU_reg_13_port, ALUout(12) => ALU_reg_12_port, 
                           ALUout(11) => ALU_reg_11_port, ALUout(10) => 
                           ALU_reg_10_port, ALUout(9) => ALU_reg_9_port, 
                           ALUout(8) => ALU_reg_8_port, ALUout(7) => 
                           ALU_reg_7_port, ALUout(6) => ALU_reg_6_port, 
                           ALUout(5) => ALU_reg_5_port, ALUout(4) => 
                           ALU_reg_4_port, ALUout(3) => ALU_reg_3_port, 
                           ALUout(2) => ALU_reg_2_port, ALUout(1) => 
                           ALU_reg_1_port, ALUout(0) => ALU_reg_0_port, 
                           MEout(31) => ME_reg_31_port, MEout(30) => 
                           ME_reg_30_port, MEout(29) => ME_reg_29_port, 
                           MEout(28) => ME_reg_28_port, MEout(27) => 
                           ME_reg_27_port, MEout(26) => ME_reg_26_port, 
                           MEout(25) => ME_reg_25_port, MEout(24) => 
                           ME_reg_24_port, MEout(23) => ME_reg_23_port, 
                           MEout(22) => ME_reg_22_port, MEout(21) => 
                           ME_reg_21_port, MEout(20) => ME_reg_20_port, 
                           MEout(19) => ME_reg_19_port, MEout(18) => 
                           ME_reg_18_port, MEout(17) => ME_reg_17_port, 
                           MEout(16) => ME_reg_16_port, MEout(15) => 
                           ME_reg_15_port, MEout(14) => ME_reg_14_port, 
                           MEout(13) => ME_reg_13_port, MEout(12) => 
                           ME_reg_12_port, MEout(11) => ME_reg_11_port, 
                           MEout(10) => ME_reg_10_port, MEout(9) => 
                           ME_reg_9_port, MEout(8) => ME_reg_8_port, MEout(7) 
                           => ME_reg_7_port, MEout(6) => ME_reg_6_port, 
                           MEout(5) => ME_reg_5_port, MEout(4) => ME_reg_4_port
                           , MEout(3) => ME_reg_3_port, MEout(2) => 
                           ME_reg_2_port, MEout(1) => ME_reg_1_port, MEout(0) 
                           => ME_reg_0_port, RDin(4) => RD_regmem_4_port, 
                           RDin(3) => RD_regmem_3_port, RDin(2) => 
                           RD_regmem_2_port, RDin(1) => RD_regmem_1_port, 
                           RDin(0) => RD_regmem_0_port, DRAM_data_out(31) => 
                           DRAM_data_out(31), DRAM_data_out(30) => 
                           DRAM_data_out(30), DRAM_data_out(29) => 
                           DRAM_data_out(29), DRAM_data_out(28) => 
                           DRAM_data_out(28), DRAM_data_out(27) => 
                           DRAM_data_out(27), DRAM_data_out(26) => 
                           DRAM_data_out(26), DRAM_data_out(25) => 
                           DRAM_data_out(25), DRAM_data_out(24) => 
                           DRAM_data_out(24), DRAM_data_out(23) => 
                           DRAM_data_out(23), DRAM_data_out(22) => 
                           DRAM_data_out(22), DRAM_data_out(21) => 
                           DRAM_data_out(21), DRAM_data_out(20) => 
                           DRAM_data_out(20), DRAM_data_out(19) => 
                           DRAM_data_out(19), DRAM_data_out(18) => 
                           DRAM_data_out(18), DRAM_data_out(17) => 
                           DRAM_data_out(17), DRAM_data_out(16) => 
                           DRAM_data_out(16), DRAM_data_out(15) => 
                           DRAM_data_out(15), DRAM_data_out(14) => 
                           DRAM_data_out(14), DRAM_data_out(13) => 
                           DRAM_data_out(13), DRAM_data_out(12) => 
                           DRAM_data_out(12), DRAM_data_out(11) => 
                           DRAM_data_out(11), DRAM_data_out(10) => 
                           DRAM_data_out(10), DRAM_data_out(9) => 
                           DRAM_data_out(9), DRAM_data_out(8) => 
                           DRAM_data_out(8), DRAM_data_out(7) => 
                           DRAM_data_out(7), DRAM_data_out(6) => 
                           DRAM_data_out(6), DRAM_data_out(5) => 
                           DRAM_data_out(5), DRAM_data_out(4) => 
                           DRAM_data_out(4), DRAM_data_out(3) => 
                           DRAM_data_out(3), DRAM_data_out(2) => 
                           DRAM_data_out(2), DRAM_data_out(1) => 
                           DRAM_data_out(1), DRAM_data_out(0) => 
                           DRAM_data_out(0), LnS => LnS, Wrd => Wrd, BHU1 => 
                           BHU1, BHU0 => BHU0, EN3 => EN3, DRAM_addr(8) => 
                           DRAM_addr(8), DRAM_addr(7) => DRAM_addr(7), 
                           DRAM_addr(6) => DRAM_addr(6), DRAM_addr(5) => 
                           DRAM_addr(5), DRAM_addr(4) => DRAM_addr(4), 
                           DRAM_addr(3) => DRAM_addr(3), DRAM_addr(2) => 
                           DRAM_addr(2), DRAM_addr(1) => DRAM_addr(1), 
                           DRAM_addr(0) => DRAM_addr(0), DRAM_data_in(31) => 
                           DRAM_data_in(31), DRAM_data_in(30) => 
                           DRAM_data_in(30), DRAM_data_in(29) => 
                           DRAM_data_in(29), DRAM_data_in(28) => 
                           DRAM_data_in(28), DRAM_data_in(27) => 
                           DRAM_data_in(27), DRAM_data_in(26) => 
                           DRAM_data_in(26), DRAM_data_in(25) => 
                           DRAM_data_in(25), DRAM_data_in(24) => 
                           DRAM_data_in(24), DRAM_data_in(23) => 
                           DRAM_data_in(23), DRAM_data_in(22) => 
                           DRAM_data_in(22), DRAM_data_in(21) => 
                           DRAM_data_in(21), DRAM_data_in(20) => 
                           DRAM_data_in(20), DRAM_data_in(19) => 
                           DRAM_data_in(19), DRAM_data_in(18) => 
                           DRAM_data_in(18), DRAM_data_in(17) => 
                           DRAM_data_in(17), DRAM_data_in(16) => 
                           DRAM_data_in(16), DRAM_data_in(15) => 
                           DRAM_data_in(15), DRAM_data_in(14) => 
                           DRAM_data_in(14), DRAM_data_in(13) => 
                           DRAM_data_in(13), DRAM_data_in(12) => 
                           DRAM_data_in(12), DRAM_data_in(11) => 
                           DRAM_data_in(11), DRAM_data_in(10) => 
                           DRAM_data_in(10), DRAM_data_in(9) => DRAM_data_in(9)
                           , DRAM_data_in(8) => DRAM_data_in(8), 
                           DRAM_data_in(7) => DRAM_data_in(7), DRAM_data_in(6) 
                           => DRAM_data_in(6), DRAM_data_in(5) => 
                           DRAM_data_in(5), DRAM_data_in(4) => DRAM_data_in(4),
                           DRAM_data_in(3) => DRAM_data_in(3), DRAM_data_in(2) 
                           => DRAM_data_in(2), DRAM_data_in(1) => 
                           DRAM_data_in(1), DRAM_data_in(0) => DRAM_data_in(0),
                           MMU_out(1) => MMU_out(1), MMU_out(0) => MMU_out(0), 
                           output(31) => mem_out_31_port, output(30) => 
                           mem_out_30_port, output(29) => mem_out_29_port, 
                           output(28) => mem_out_28_port, output(27) => 
                           mem_out_27_port, output(26) => mem_out_26_port, 
                           output(25) => mem_out_25_port, output(24) => 
                           mem_out_24_port, output(23) => mem_out_23_port, 
                           output(22) => mem_out_22_port, output(21) => 
                           mem_out_21_port, output(20) => mem_out_20_port, 
                           output(19) => mem_out_19_port, output(18) => 
                           mem_out_18_port, output(17) => mem_out_17_port, 
                           output(16) => mem_out_16_port, output(15) => 
                           mem_out_15_port, output(14) => mem_out_14_port, 
                           output(13) => mem_out_13_port, output(12) => 
                           mem_out_12_port, output(11) => mem_out_11_port, 
                           output(10) => mem_out_10_port, output(9) => 
                           mem_out_9_port, output(8) => mem_out_8_port, 
                           output(7) => mem_out_7_port, output(6) => 
                           mem_out_6_port, output(5) => mem_out_5_port, 
                           output(4) => mem_out_4_port, output(3) => 
                           mem_out_3_port, output(2) => mem_out_2_port, 
                           output(1) => mem_out_1_port, output(0) => 
                           mem_out_0_port, alu_out(31) => ALU_memout_31_port, 
                           alu_out(30) => ALU_memout_30_port, alu_out(29) => 
                           ALU_memout_29_port, alu_out(28) => 
                           ALU_memout_28_port, alu_out(27) => 
                           ALU_memout_27_port, alu_out(26) => 
                           ALU_memout_26_port, alu_out(25) => 
                           ALU_memout_25_port, alu_out(24) => 
                           ALU_memout_24_port, alu_out(23) => 
                           ALU_memout_23_port, alu_out(22) => 
                           ALU_memout_22_port, alu_out(21) => 
                           ALU_memout_21_port, alu_out(20) => 
                           ALU_memout_20_port, alu_out(19) => 
                           ALU_memout_19_port, alu_out(18) => 
                           ALU_memout_18_port, alu_out(17) => 
                           ALU_memout_17_port, alu_out(16) => 
                           ALU_memout_16_port, alu_out(15) => 
                           ALU_memout_15_port, alu_out(14) => 
                           ALU_memout_14_port, alu_out(13) => 
                           ALU_memout_13_port, alu_out(12) => 
                           ALU_memout_12_port, alu_out(11) => 
                           ALU_memout_11_port, alu_out(10) => 
                           ALU_memout_10_port, alu_out(9) => ALU_memout_9_port,
                           alu_out(8) => ALU_memout_8_port, alu_out(7) => 
                           ALU_memout_7_port, alu_out(6) => ALU_memout_6_port, 
                           alu_out(5) => ALU_memout_5_port, alu_out(4) => 
                           ALU_memout_4_port, alu_out(3) => ALU_memout_3_port, 
                           alu_out(2) => ALU_memout_2_port, alu_out(1) => 
                           ALU_memout_1_port, alu_out(0) => ALU_memout_0_port, 
                           RDout(4) => RD_memout_4_port, RDout(3) => 
                           RD_memout_3_port, RDout(2) => RD_memout_2_port, 
                           RDout(1) => RD_memout_1_port, RDout(0) => 
                           RD_memout_0_port);
   wb_stage : WB port map( mem_out(31) => LMD_reg_31_port, mem_out(30) => 
                           LMD_reg_30_port, mem_out(29) => LMD_reg_29_port, 
                           mem_out(28) => LMD_reg_28_port, mem_out(27) => 
                           LMD_reg_27_port, mem_out(26) => LMD_reg_26_port, 
                           mem_out(25) => LMD_reg_25_port, mem_out(24) => 
                           LMD_reg_24_port, mem_out(23) => LMD_reg_23_port, 
                           mem_out(22) => LMD_reg_22_port, mem_out(21) => 
                           LMD_reg_21_port, mem_out(20) => LMD_reg_20_port, 
                           mem_out(19) => LMD_reg_19_port, mem_out(18) => 
                           LMD_reg_18_port, mem_out(17) => LMD_reg_17_port, 
                           mem_out(16) => LMD_reg_16_port, mem_out(15) => 
                           LMD_reg_15_port, mem_out(14) => LMD_reg_14_port, 
                           mem_out(13) => LMD_reg_13_port, mem_out(12) => 
                           LMD_reg_12_port, mem_out(11) => LMD_reg_11_port, 
                           mem_out(10) => LMD_reg_10_port, mem_out(9) => 
                           LMD_reg_9_port, mem_out(8) => LMD_reg_8_port, 
                           mem_out(7) => LMD_reg_7_port, mem_out(6) => 
                           LMD_reg_6_port, mem_out(5) => LMD_reg_5_port, 
                           mem_out(4) => LMD_reg_4_port, mem_out(3) => 
                           LMD_reg_3_port, mem_out(2) => LMD_reg_2_port, 
                           mem_out(1) => LMD_reg_1_port, mem_out(0) => 
                           LMD_reg_0_port, alu_out(31) => ALU_regmem_31_port, 
                           alu_out(30) => ALU_regmem_30_port, alu_out(29) => 
                           ALU_regmem_29_port, alu_out(28) => 
                           ALU_regmem_28_port, alu_out(27) => 
                           ALU_regmem_27_port, alu_out(26) => 
                           ALU_regmem_26_port, alu_out(25) => 
                           ALU_regmem_25_port, alu_out(24) => 
                           ALU_regmem_24_port, alu_out(23) => 
                           ALU_regmem_23_port, alu_out(22) => 
                           ALU_regmem_22_port, alu_out(21) => 
                           ALU_regmem_21_port, alu_out(20) => 
                           ALU_regmem_20_port, alu_out(19) => 
                           ALU_regmem_19_port, alu_out(18) => 
                           ALU_regmem_18_port, alu_out(17) => 
                           ALU_regmem_17_port, alu_out(16) => 
                           ALU_regmem_16_port, alu_out(15) => 
                           ALU_regmem_15_port, alu_out(14) => 
                           ALU_regmem_14_port, alu_out(13) => 
                           ALU_regmem_13_port, alu_out(12) => 
                           ALU_regmem_12_port, alu_out(11) => 
                           ALU_regmem_11_port, alu_out(10) => 
                           ALU_regmem_10_port, alu_out(9) => ALU_regmem_9_port,
                           alu_out(8) => ALU_regmem_8_port, alu_out(7) => 
                           ALU_regmem_7_port, alu_out(6) => ALU_regmem_6_port, 
                           alu_out(5) => ALU_regmem_5_port, alu_out(4) => 
                           ALU_regmem_4_port, alu_out(3) => ALU_regmem_3_port, 
                           alu_out(2) => ALU_regmem_2_port, alu_out(1) => 
                           ALU_regmem_1_port, alu_out(0) => ALU_regmem_0_port, 
                           S3 => S3, output(31) => WB_data_31_port, output(30) 
                           => WB_data_30_port, output(29) => WB_data_29_port, 
                           output(28) => WB_data_28_port, output(27) => 
                           WB_data_27_port, output(26) => WB_data_26_port, 
                           output(25) => WB_data_25_port, output(24) => 
                           WB_data_24_port, output(23) => WB_data_23_port, 
                           output(22) => WB_data_22_port, output(21) => 
                           WB_data_21_port, output(20) => WB_data_20_port, 
                           output(19) => WB_data_19_port, output(18) => 
                           WB_data_18_port, output(17) => WB_data_17_port, 
                           output(16) => WB_data_16_port, output(15) => 
                           WB_data_15_port, output(14) => WB_data_14_port, 
                           output(13) => WB_data_13_port, output(12) => 
                           WB_data_12_port, output(11) => WB_data_11_port, 
                           output(10) => WB_data_10_port, output(9) => 
                           WB_data_9_port, output(8) => WB_data_8_port, 
                           output(7) => WB_data_7_port, output(6) => 
                           WB_data_6_port, output(5) => WB_data_5_port, 
                           output(4) => WB_data_4_port, output(3) => 
                           WB_data_3_port, output(2) => WB_data_2_port, 
                           output(1) => WB_data_1_port, output(0) => 
                           WB_data_0_port);
   IR_reg_reg_30_inst : DFFS_X2 port map( D => NOP_MUX_OUT_30_port, CK => CLK, 
                           SN => n12, Q => IR_reg_30_port, QN => n_2321);
   IR_reg_reg_28_inst : DFFS_X1 port map( D => NOP_MUX_OUT_28_port, CK => CLK, 
                           SN => n12, Q => IR_reg_28_port, QN => n_2322);
   U3 : BUF_X2 port map( A => n2, Z => n9);
   U4 : BUF_X2 port map( A => n3, Z => n10);
   U5 : BUF_X2 port map( A => n3, Z => n11);
   U6 : BUF_X2 port map( A => n1, Z => n5);
   U7 : BUF_X2 port map( A => n1, Z => n6);
   U8 : BUF_X2 port map( A => n2, Z => n7);
   U9 : BUF_X2 port map( A => n2, Z => n8);
   U10 : BUF_X2 port map( A => n1, Z => n4);
   U11 : BUF_X1 port map( A => n3, Z => n12);
   U12 : BUF_X1 port map( A => RST, Z => n1);
   U13 : BUF_X1 port map( A => RST, Z => n3);
   U14 : BUF_X1 port map( A => RST, Z => n2);

end SYN_Structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity hardwired_CU is

   port( clk, rst : in std_logic;  opcode : in std_logic_vector (5 downto 0);  
         func : in std_logic_vector (10 downto 0);  RF1, RF2, EN1, S1, S2, ALU3
         , ALU2, ALU1, ALU0, SN, LnS, Wrd, BHU1, BHU0, EN3, S3, WF1, Ld : out 
         std_logic);

end hardwired_CU;

architecture SYN_Behavioral of hardwired_CU is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component SDFFR_X1
      port( D, SI, SE, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Ld_port, cw2_5_port, cw2_4_port, cw2_3_port, cw2_2_port, cw2_1_port, 
      cw2_0_port, cw3_1_port, cw3_0_port, cw21_6_port, cw21_5_port, cw21_4_port
      , cw21_3_port, cw21_2_port, cw21_1_port, cw21_0_port, cw22_6_port, 
      cw22_5_port, cw22_4_port, cw22_3_port, cw22_2_port, cw22_1_port, 
      cw22_0_port, cw23_6_port, cw23_5_port, cw23_4_port, cw23_3_port, 
      cw23_2_port, cw23_1_port, cw23_0_port, exe_type2, exe_type21, exe_type22,
      exe_type23, cw1_13_port, cw1_12_port, cw1_11_port, cw1_10_port, 
      cw1_9_port, cw1_8_port, cw1_7_port, cw1_6_port, cw1_5_port, cw1_4_port, 
      cw1_3_port, cw1_2_port, cw1_1_port, cw1_0_port, N190, n1, n38, n39, n40, 
      n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55
      , n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, 
      n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84
      , n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, 
      n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, 
      n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, 
      n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, 
      n135, n136, n137, n138, n139, n140, n141, n2, n3, n4, n5, n6, n7, n8, n9,
      n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24
      , n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n142, 
      n143, n144, n145, n146, n_2323, n_2324, n_2325, n_2326, n_2327, n_2328, 
      n_2329, n_2330, n_2331, n_2332, n_2333, n_2334, n_2335, n_2336, n_2337, 
      n_2338, n_2339, n_2340, n_2341, n_2342, n_2343, n_2344, n_2345, n_2346, 
      n_2347, n_2348, n_2349, n_2350, n_2351, n_2352, n_2353, n_2354, n_2355, 
      n_2356, n_2357, n_2358, n_2359, n_2360, n_2361, n_2362, n_2363, n_2364, 
      n_2365, n_2366, n_2367, n_2368, n_2369 : std_logic;

begin
   Ld <= Ld_port;
   
   cw2_reg_13_inst : DFFR_X1 port map( D => cw1_13_port, CK => clk, RN => n4, Q
                           => S1, QN => n_2323);
   cw2_reg_12_inst : DFFR_X1 port map( D => cw1_12_port, CK => clk, RN => n2, Q
                           => S2, QN => n_2324);
   cw2_reg_11_inst : DFFR_X1 port map( D => cw1_11_port, CK => clk, RN => n2, Q
                           => ALU3, QN => n_2325);
   cw2_reg_10_inst : DFFR_X1 port map( D => cw1_10_port, CK => clk, RN => n2, Q
                           => ALU2, QN => n_2326);
   cw2_reg_9_inst : DFFR_X1 port map( D => cw1_9_port, CK => clk, RN => n2, Q 
                           => ALU1, QN => n_2327);
   cw2_reg_8_inst : DFFR_X1 port map( D => cw1_8_port, CK => clk, RN => n2, Q 
                           => ALU0, QN => n_2328);
   cw2_reg_7_inst : DFFR_X1 port map( D => cw1_7_port, CK => clk, RN => n2, Q 
                           => SN, QN => n_2329);
   cw2_reg_6_inst : DFFR_X1 port map( D => cw1_6_port, CK => clk, RN => n2, Q 
                           => Ld_port, QN => n_2330);
   cw2_reg_5_inst : DFFR_X1 port map( D => cw1_5_port, CK => clk, RN => n2, Q 
                           => cw2_5_port, QN => n_2331);
   cw2_reg_4_inst : DFFR_X1 port map( D => cw1_4_port, CK => clk, RN => n2, Q 
                           => cw2_4_port, QN => n_2332);
   cw2_reg_3_inst : DFFR_X1 port map( D => cw1_3_port, CK => clk, RN => n2, Q 
                           => cw2_3_port, QN => n_2333);
   cw2_reg_2_inst : DFFR_X1 port map( D => cw1_2_port, CK => clk, RN => n3, Q 
                           => cw2_2_port, QN => n_2334);
   cw2_reg_1_inst : DFFR_X1 port map( D => cw1_1_port, CK => clk, RN => n3, Q 
                           => cw2_1_port, QN => n_2335);
   cw2_reg_0_inst : DFFR_X1 port map( D => cw1_0_port, CK => clk, RN => n3, Q 
                           => cw2_0_port, QN => n_2336);
   cw21_reg_6_inst : DFFR_X1 port map( D => Ld_port, CK => clk, RN => n3, Q => 
                           cw21_6_port, QN => n_2337);
   cw21_reg_5_inst : DFFR_X1 port map( D => cw2_5_port, CK => clk, RN => n3, Q 
                           => cw21_5_port, QN => n_2338);
   cw21_reg_4_inst : DFFR_X1 port map( D => cw2_4_port, CK => clk, RN => n3, Q 
                           => cw21_4_port, QN => n_2339);
   cw21_reg_3_inst : DFFR_X1 port map( D => cw2_3_port, CK => clk, RN => n3, Q 
                           => cw21_3_port, QN => n_2340);
   cw21_reg_2_inst : DFFR_X1 port map( D => cw2_2_port, CK => clk, RN => n3, Q 
                           => cw21_2_port, QN => n_2341);
   cw21_reg_1_inst : DFFR_X1 port map( D => cw2_1_port, CK => clk, RN => n3, Q 
                           => cw21_1_port, QN => n_2342);
   cw21_reg_0_inst : DFFR_X1 port map( D => cw2_0_port, CK => clk, RN => n3, Q 
                           => cw21_0_port, QN => n_2343);
   cw22_reg_6_inst : DFFR_X1 port map( D => cw21_6_port, CK => clk, RN => n3, Q
                           => cw22_6_port, QN => n_2344);
   cw22_reg_5_inst : DFFR_X1 port map( D => cw21_5_port, CK => clk, RN => n4, Q
                           => cw22_5_port, QN => n_2345);
   cw22_reg_4_inst : DFFR_X1 port map( D => cw21_4_port, CK => clk, RN => n4, Q
                           => cw22_4_port, QN => n_2346);
   cw22_reg_3_inst : DFFR_X1 port map( D => cw21_3_port, CK => clk, RN => n4, Q
                           => cw22_3_port, QN => n_2347);
   cw22_reg_2_inst : DFFR_X1 port map( D => cw21_2_port, CK => clk, RN => n4, Q
                           => cw22_2_port, QN => n_2348);
   cw22_reg_1_inst : DFFR_X1 port map( D => cw21_1_port, CK => clk, RN => n4, Q
                           => cw22_1_port, QN => n_2349);
   cw22_reg_0_inst : DFFR_X1 port map( D => cw21_0_port, CK => clk, RN => n4, Q
                           => cw22_0_port, QN => n_2350);
   cw23_reg_6_inst : DFFR_X1 port map( D => cw22_6_port, CK => clk, RN => n4, Q
                           => cw23_6_port, QN => n_2351);
   cw23_reg_5_inst : DFFR_X1 port map( D => cw22_5_port, CK => clk, RN => n4, Q
                           => cw23_5_port, QN => n_2352);
   cw23_reg_4_inst : DFFR_X1 port map( D => cw22_4_port, CK => clk, RN => n4, Q
                           => cw23_4_port, QN => n_2353);
   cw23_reg_3_inst : DFFR_X1 port map( D => cw22_3_port, CK => clk, RN => n4, Q
                           => cw23_3_port, QN => n_2354);
   cw23_reg_2_inst : DFFR_X1 port map( D => cw22_2_port, CK => clk, RN => n5, Q
                           => cw23_2_port, QN => n_2355);
   cw23_reg_1_inst : DFFR_X1 port map( D => cw22_1_port, CK => clk, RN => n5, Q
                           => cw23_1_port, QN => n_2356);
   cw23_reg_0_inst : DFFR_X1 port map( D => cw22_0_port, CK => clk, RN => n5, Q
                           => cw23_0_port, QN => n_2357);
   exe_type2_reg : DFFR_X1 port map( D => N190, CK => clk, RN => n5, Q => 
                           exe_type2, QN => n_2358);
   exe_type21_reg : DFFR_X1 port map( D => exe_type2, CK => clk, RN => n5, Q =>
                           exe_type21, QN => n_2359);
   exe_type22_reg : DFFR_X1 port map( D => exe_type21, CK => clk, RN => n5, Q 
                           => exe_type22, QN => n_2360);
   exe_type23_reg : DFFR_X1 port map( D => exe_type22, CK => clk, RN => n5, Q 
                           => exe_type23, QN => n1);
   cw3_reg_6_inst : SDFFR_X1 port map( D => cw23_6_port, SI => Ld_port, SE => 
                           n1, CK => clk, RN => n5, Q => LnS, QN => n_2361);
   cw3_reg_5_inst : SDFFR_X1 port map( D => cw2_5_port, SI => cw23_5_port, SE 
                           => exe_type23, CK => clk, RN => n5, Q => Wrd, QN => 
                           n_2362);
   cw3_reg_4_inst : SDFFR_X1 port map( D => cw2_4_port, SI => cw23_4_port, SE 
                           => exe_type23, CK => clk, RN => n5, Q => BHU1, QN =>
                           n_2363);
   cw3_reg_3_inst : SDFFR_X1 port map( D => cw2_3_port, SI => cw23_3_port, SE 
                           => exe_type23, CK => clk, RN => n6, Q => BHU0, QN =>
                           n_2364);
   cw3_reg_2_inst : SDFFR_X1 port map( D => cw2_2_port, SI => cw23_2_port, SE 
                           => exe_type23, CK => clk, RN => n6, Q => EN3, QN => 
                           n_2365);
   cw3_reg_1_inst : SDFFR_X1 port map( D => cw2_1_port, SI => cw23_1_port, SE 
                           => exe_type23, CK => clk, RN => n6, Q => cw3_1_port,
                           QN => n_2366);
   cw4_reg_1_inst : DFFR_X1 port map( D => cw3_1_port, CK => clk, RN => n5, Q 
                           => S3, QN => n_2367);
   cw3_reg_0_inst : SDFFR_X1 port map( D => cw2_0_port, SI => cw23_0_port, SE 
                           => exe_type23, CK => clk, RN => n6, Q => cw3_0_port,
                           QN => n_2368);
   cw4_reg_0_inst : DFFR_X1 port map( D => cw3_0_port, CK => clk, RN => n2, Q 
                           => WF1, QN => n_2369);
   U147 : NAND3_X1 port map( A1 => n23, A2 => n19, A3 => opcode(4), ZN => n52);
   U148 : OAI33_X1 port map( A1 => n46, A2 => n77, A3 => n36, B1 => n78, B2 => 
                           n30, B3 => n79, ZN => n76);
   U149 : NAND3_X1 port map( A1 => opcode(5), A2 => opcode(1), A3 => n115, ZN 
                           => n114);
   U150 : NAND3_X1 port map( A1 => n20, A2 => n13, A3 => n24, ZN => n124);
   U151 : NAND3_X1 port map( A1 => func(0), A2 => n36, A3 => func(1), ZN => 
                           n119);
   U152 : NAND3_X1 port map( A1 => n128, A2 => n143, A3 => func(5), ZN => n46);
   U153 : NAND3_X1 port map( A1 => n30, A2 => n36, A3 => func(1), ZN => n98);
   U154 : NAND3_X1 port map( A1 => func(3), A2 => n128, A3 => func(5), ZN => 
                           n118);
   U155 : NAND3_X1 port map( A1 => n30, A2 => n34, A3 => func(2), ZN => n47);
   U156 : NAND3_X1 port map( A1 => n75, A2 => n48, A3 => n94, ZN => n125);
   U157 : NAND3_X1 port map( A1 => n143, A2 => n146, A3 => n128, ZN => n78);
   U158 : NAND3_X1 port map( A1 => opcode(3), A2 => n19, A3 => opcode(1), ZN =>
                           n68);
   U159 : NAND3_X1 port map( A1 => n22, A2 => opcode(5), A3 => n90, ZN => n138)
                           ;
   U160 : NAND3_X1 port map( A1 => n27, A2 => n19, A3 => n8, ZN => n140);
   U3 : NOR2_X1 port map( A1 => n144, A2 => n142, ZN => n45);
   U4 : INV_X1 port map( A => n78, ZN => n37);
   U5 : NAND2_X1 port map( A1 => n37, A2 => n35, ZN => n94);
   U6 : INV_X1 port map( A => n73, ZN => n33);
   U7 : INV_X1 port map( A => n99, ZN => n28);
   U8 : OAI22_X1 port map( A1 => n78, A2 => n47, B1 => n45, B2 => n98, ZN => 
                           n70);
   U9 : NOR3_X1 port map( A1 => n77, A2 => n116, A3 => n36, ZN => n74);
   U10 : AOI21_X1 port map( B1 => n45, B2 => n78, A => n119, ZN => n127);
   U11 : AOI21_X1 port map( B1 => n45, B2 => n46, A => n47, ZN => n42);
   U12 : NOR3_X1 port map( A1 => n102, A2 => n26, A3 => n103, ZN => cw1_4_port)
                           ;
   U13 : NOR2_X1 port map( A1 => n118, A2 => n77, ZN => n73);
   U14 : NAND2_X1 port map( A1 => n80, A2 => n47, ZN => n99);
   U15 : NAND4_X1 port map( A1 => n117, A2 => n33, A3 => n75, A4 => n48, ZN => 
                           n93);
   U16 : OAI21_X1 port map( B1 => n97, B2 => n99, A => n144, ZN => n117);
   U17 : NOR2_X1 port map( A1 => n100, A2 => n101, ZN => cw1_5_port);
   U18 : INV_X1 port map( A => n85, ZN => n24);
   U19 : INV_X1 port map( A => n103, ZN => n8);
   U20 : INV_X1 port map( A => n90, ZN => n14);
   U21 : INV_X1 port map( A => n98, ZN => n29);
   U22 : INV_X1 port map( A => n118, ZN => n144);
   U23 : INV_X1 port map( A => n134, ZN => n21);
   U24 : INV_X1 port map( A => n79, ZN => n35);
   U25 : INV_X1 port map( A => n68, ZN => n16);
   U26 : INV_X1 port map( A => n102, ZN => n17);
   U27 : INV_X1 port map( A => n116, ZN => n142);
   U28 : AND2_X1 port map( A1 => n98, A2 => n119, ZN => n80);
   U29 : OR2_X1 port map( A1 => n8, A2 => n57, ZN => n54);
   U30 : NOR2_X1 port map( A1 => n97, A2 => n29, ZN => n96);
   U31 : INV_X1 port map( A => n48, ZN => n32);
   U32 : NAND2_X1 port map( A1 => n109, A2 => n139, ZN => EN1);
   U33 : OAI21_X1 port map( B1 => n18, B2 => n137, A => n26, ZN => n139);
   U34 : INV_X1 port map( A => n101, ZN => n18);
   U35 : NAND2_X1 port map( A1 => n41, A2 => n135, ZN => RF2);
   U36 : OR3_X1 port map( A1 => n104, A2 => n25, A3 => n100, ZN => n135);
   U37 : NAND2_X1 port map( A1 => n109, A2 => n7, ZN => RF1);
   U38 : NOR2_X1 port map( A1 => n134, A2 => n13, ZN => n141);
   U39 : NOR4_X1 port map( A1 => n145, A2 => n143, A3 => n130, A4 => func(6), 
                           ZN => n129);
   U40 : INV_X1 port map( A => func(4), ZN => n145);
   U41 : INV_X1 port map( A => n67, ZN => n12);
   U42 : NOR3_X1 port map( A1 => func(4), A2 => func(6), A3 => n130, ZN => n128
                           );
   U43 : AOI211_X1 port map( C1 => n13, C2 => n27, A => n19, B => n23, ZN => 
                           n111);
   U44 : OAI211_X1 port map( C1 => n81, C2 => n41, A => n58, B => n82, ZN => 
                           cw1_7_port);
   U45 : NOR3_X1 port map( A1 => n92, A2 => n43, A3 => n93, ZN => n81);
   U46 : OAI22_X1 port map( A1 => n28, A2 => n78, B1 => n96, B2 => n46, ZN => 
                           n92);
   U47 : NAND4_X1 port map( A1 => n17, A2 => n8, A3 => n27, A4 => n26, ZN => 
                           n41);
   U48 : NOR2_X1 port map( A1 => n19, A2 => n53, ZN => n90);
   U49 : NAND4_X1 port map( A1 => n35, A2 => n129, A3 => func(0), A4 => n146, 
                           ZN => n75);
   U50 : INV_X1 port map( A => n110, ZN => n9);
   U51 : OAI211_X1 port map( C1 => n25, C2 => n111, A => n14, B => n101, ZN => 
                           n110);
   U52 : NOR4_X1 port map( A1 => n20, A2 => n27, A3 => n26, A4 => n103, ZN => 
                           cw1_3_port);
   U53 : NAND2_X1 port map( A1 => func(0), A2 => n34, ZN => n77);
   U54 : OAI221_X1 port map( B1 => n13, B2 => n68, C1 => n121, C2 => n41, A => 
                           n122, ZN => cw1_10_port);
   U55 : NOR4_X1 port map( A1 => n125, A2 => n70, A3 => n126, A4 => n127, ZN =>
                           n121);
   U56 : AOI221_X1 port map( B1 => n90, B2 => n22, C1 => n15, C2 => n24, A => 
                           n123, ZN => n122);
   U57 : NOR3_X1 port map( A1 => n46, A2 => func(0), A3 => n79, ZN => n126);
   U58 : OAI221_X1 port map( B1 => n112, B2 => n13, C1 => n113, C2 => n41, A =>
                           n114, ZN => cw1_11_port);
   U59 : AOI211_X1 port map( C1 => n142, C2 => n99, A => n93, B => n74, ZN => 
                           n113);
   U60 : OAI221_X1 port map( B1 => n58, B2 => n27, C1 => n59, C2 => n41, A => 
                           n60, ZN => cw1_8_port);
   U61 : NOR3_X1 port map( A1 => n69, A2 => n44, A3 => n70, ZN => n59);
   U62 : AOI221_X1 port map( B1 => n61, B2 => n26, C1 => n15, C2 => n62, A => 
                           n63, ZN => n60);
   U63 : OAI21_X1 port map( B1 => n80, B2 => n46, A => n33, ZN => n69);
   U64 : NOR2_X1 port map( A1 => n23, A2 => n27, ZN => n57);
   U65 : NAND2_X1 port map( A1 => n19, A2 => n25, ZN => n102);
   U66 : OAI21_X1 port map( B1 => n111, B2 => n25, A => n140, ZN => n137);
   U67 : NAND2_X1 port map( A1 => n13, A2 => n23, ZN => n103);
   U68 : NAND2_X1 port map( A1 => func(1), A2 => func(2), ZN => n79);
   U69 : INV_X1 port map( A => func(2), ZN => n36);
   U70 : NAND2_X1 port map( A1 => n57, A2 => n19, ZN => n101);
   U71 : NAND2_X1 port map( A1 => n85, A2 => n19, ZN => n104);
   U72 : AOI21_X1 port map( B1 => n25, B2 => n65, A => n19, ZN => n120);
   U73 : OAI21_X1 port map( B1 => n8, B2 => n19, A => n53, ZN => n49);
   U74 : INV_X1 port map( A => func(0), ZN => n30);
   U75 : NAND2_X1 port map( A1 => n115, A2 => n23, ZN => n67);
   U76 : INV_X1 port map( A => n66, ZN => n20);
   U77 : INV_X1 port map( A => n136, ZN => n7);
   U78 : NAND2_X1 port map( A1 => func(5), A2 => n129, ZN => n116);
   U79 : OAI21_X1 port map( B1 => n53, B2 => n85, A => n10, ZN => n84);
   U80 : INV_X1 port map( A => n86, ZN => n10);
   U81 : INV_X1 port map( A => n107, ZN => n15);
   U82 : NAND2_X1 port map( A1 => n85, A2 => n66, ZN => n50);
   U83 : INV_X1 port map( A => func(1), ZN => n34);
   U84 : INV_X1 port map( A => func(5), ZN => n146);
   U85 : NAND2_X1 port map( A1 => n71, A2 => n72, ZN => n44);
   U86 : AOI211_X1 port map( C1 => n73, C2 => func(2), A => n74, B => n31, ZN 
                           => n72);
   U87 : AOI21_X1 port map( B1 => n29, B2 => n37, A => n76, ZN => n71);
   U88 : INV_X1 port map( A => n75, ZN => n31);
   U89 : INV_X1 port map( A => n65, ZN => n22);
   U90 : INV_X1 port map( A => func(3), ZN => n143);
   U91 : NAND2_X1 port map( A1 => n94, A2 => n95, ZN => n43);
   U92 : OR3_X1 port map( A1 => n77, A2 => func(2), A3 => n78, ZN => n95);
   U93 : NAND2_X1 port map( A1 => n75, A2 => n138, ZN => N190);
   U94 : NOR3_X1 port map( A1 => func(1), A2 => func(2), A3 => func(0), ZN => 
                           n97);
   U95 : NAND4_X1 port map( A1 => func(3), A2 => n97, A3 => n128, A4 => n146, 
                           ZN => n48);
   U96 : NOR4_X1 port map( A1 => n32, A2 => n42, A3 => n43, A4 => n44, ZN => 
                           n40);
   U97 : AOI221_X1 port map( B1 => n20, B2 => opcode(4), C1 => opcode(2), C2 =>
                           n54, A => n55, ZN => n38);
   U98 : INV_X1 port map( A => n132, ZN => n11);
   U99 : AOI21_X1 port map( B1 => n104, B2 => n105, A => n100, ZN => cw1_2_port
                           );
   U100 : OAI21_X1 port map( B1 => n131, B2 => n26, A => n7, ZN => cw1_0_port);
   U101 : OAI21_X1 port map( B1 => n106, B2 => n107, A => n7, ZN => cw1_1_port)
                           ;
   U102 : OR4_X1 port map( A1 => func(7), A2 => func(10), A3 => func(9), A4 => 
                           func(8), ZN => n130);
   U103 : NAND2_X1 port map( A1 => n52, A2 => n14, ZN => n51);
   U104 : NOR3_X1 port map( A1 => opcode(1), A2 => opcode(5), A3 => n25, ZN => 
                           n89);
   U105 : AOI211_X1 port map( C1 => opcode(1), C2 => n90, A => n12, B => n137, 
                           ZN => n108);
   U106 : NOR3_X1 port map( A1 => opcode(1), A2 => opcode(3), A3 => n115, ZN =>
                           n132);
   U107 : AOI21_X1 port map( B1 => opcode(3), B2 => opcode(1), A => n50, ZN => 
                           n134);
   U108 : NAND2_X1 port map( A1 => opcode(1), A2 => n27, ZN => n85);
   U109 : INV_X1 port map( A => opcode(1), ZN => n23);
   U110 : AOI21_X1 port map( B1 => n23, B2 => n56, A => opcode(3), ZN => n55);
   U111 : AND3_X1 port map( A1 => n64, A2 => opcode(4), A3 => opcode(3), ZN => 
                           n63);
   U112 : OAI21_X1 port map( B1 => opcode(3), B2 => n65, A => n66, ZN => n62);
   U113 : OAI222_X1 port map( A1 => n66, A2 => n65, B1 => opcode(3), B2 => n67,
                           C1 => opcode(4), C2 => n68, ZN => n61);
   U114 : AOI22_X1 port map( A1 => opcode(3), A2 => n88, B1 => n57, B2 => n25, 
                           ZN => n87);
   U115 : NOR3_X1 port map( A1 => n100, A2 => opcode(3), A3 => n64, ZN => 
                           cw1_6_port);
   U116 : NAND2_X1 port map( A1 => opcode(3), A2 => opcode(2), ZN => n66);
   U117 : INV_X1 port map( A => opcode(3), ZN => n25);
   U118 : OAI222_X1 port map( A1 => opcode(5), A2 => n38, B1 => n39, B2 => n26,
                           C1 => n40, C2 => n41, ZN => cw1_9_port);
   U119 : AOI22_X1 port map( A1 => n83, A2 => n26, B1 => opcode(5), B2 => n84, 
                           ZN => n82);
   U120 : NOR2_X1 port map( A1 => n23, A2 => opcode(5), ZN => n91);
   U121 : OAI21_X1 port map( B1 => opcode(5), B2 => n108, A => n109, ZN => 
                           cw1_13_port);
   U122 : OAI21_X1 port map( B1 => opcode(5), B2 => n9, A => n109, ZN => 
                           cw1_12_port);
   U123 : AOI211_X1 port map( C1 => n120, C2 => opcode(5), A => n16, B => n89, 
                           ZN => n112);
   U124 : AOI21_X1 port map( B1 => n14, B2 => n124, A => opcode(5), ZN => n123)
                           ;
   U125 : NAND2_X1 port map( A1 => opcode(5), A2 => opcode(4), ZN => n107);
   U126 : NAND2_X1 port map( A1 => opcode(5), A2 => n13, ZN => n100);
   U127 : AOI21_X1 port map( B1 => n101, B2 => n108, A => opcode(5), ZN => n136
                           );
   U128 : OAI21_X1 port map( B1 => n141, B2 => n86, A => opcode(5), ZN => n109)
                           ;
   U129 : INV_X1 port map( A => opcode(5), ZN => n26);
   U130 : AOI221_X1 port map( B1 => opcode(0), B2 => n49, C1 => n50, C2 => n13,
                           A => n51, ZN => n39);
   U131 : OAI21_X1 port map( B1 => opcode(0), B2 => opcode(4), A => n19, ZN => 
                           n56);
   U132 : NAND2_X1 port map( A1 => opcode(0), A2 => n13, ZN => n88);
   U133 : NAND2_X1 port map( A1 => opcode(0), A2 => n23, ZN => n65);
   U134 : NOR3_X1 port map( A1 => n13, A2 => opcode(0), A3 => n19, ZN => n115);
   U135 : INV_X1 port map( A => opcode(0), ZN => n27);
   U136 : AOI22_X1 port map( A1 => opcode(4), A2 => n89, B1 => n90, B2 => n91, 
                           ZN => n58);
   U137 : AOI211_X1 port map( C1 => opcode(4), C2 => n21, A => n132, B => n133,
                           ZN => n131);
   U138 : NOR3_X1 port map( A1 => n102, A2 => opcode(4), A3 => n27, ZN => n133)
                           ;
   U139 : NAND2_X1 port map( A1 => opcode(4), A2 => n25, ZN => n53);
   U140 : OAI21_X1 port map( B1 => opcode(4), B2 => n104, A => n11, ZN => n86);
   U141 : INV_X1 port map( A => opcode(4), ZN => n13);
   U142 : OAI21_X1 port map( B1 => opcode(2), B2 => n87, A => n67, ZN => n83);
   U143 : NOR2_X1 port map( A1 => n85, A2 => opcode(2), ZN => n64);
   U144 : NAND2_X1 port map( A1 => opcode(2), A2 => n25, ZN => n105);
   U145 : AOI221_X1 port map( B1 => n17, B2 => n23, C1 => n22, C2 => opcode(2),
                           A => n21, ZN => n106);
   U146 : INV_X1 port map( A => opcode(2), ZN => n19);
   U161 : CLKBUF_X1 port map( A => rst, Z => n2);
   U162 : CLKBUF_X1 port map( A => rst, Z => n3);
   U163 : CLKBUF_X1 port map( A => rst, Z => n4);
   U164 : CLKBUF_X1 port map( A => rst, Z => n5);
   U165 : CLKBUF_X1 port map( A => rst, Z => n6);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_MEM_SIZE128_WORD_size32_NREG32.all;

entity DLX_MEM_SIZE128_WORD_size32_NREG32 is

   port( CLK, RST : in std_logic;  from_DRAM_data, IRAM_data : in 
         std_logic_vector (31 downto 0);  DRAM_addr : out std_logic_vector (8 
         downto 0);  IRAM_addr : out std_logic_vector (7 downto 0);  
         to_DRAM_data : out std_logic_vector (31 downto 0);  DRAM_EN, DRAM_LnS 
         : out std_logic;  MMU_out : out std_logic_vector (1 downto 0));

end DLX_MEM_SIZE128_WORD_size32_NREG32;

architecture SYN_Structural of DLX_MEM_SIZE128_WORD_size32_NREG32 is

   component DataPath_MEM_SIZE128_WORD_size32_NREG32
      port( CLK, RST, RF1, RF2, EN1, S1, S2, ALU3, ALU2, ALU1, ALU0, SN, LnS, 
            BHU1, BHU0, Wrd, EN3, S3, WF1, Ld : in std_logic;  instr : in 
            std_logic_vector (31 downto 0);  IRAM_addr : out std_logic_vector 
            (31 downto 0);  DRAM_data_out : in std_logic_vector (31 downto 0); 
            MMU_out : out std_logic_vector (1 downto 0);  DRAM_addr : out 
            std_logic_vector (8 downto 0);  DRAM_data_in : out std_logic_vector
            (31 downto 0);  opcode : out std_logic_vector (5 downto 0);  func :
            out std_logic_vector (10 downto 0);  OVF : out std_logic);
   end component;
   
   component hardwired_CU
      port( clk, rst : in std_logic;  opcode : in std_logic_vector (5 downto 0)
            ;  func : in std_logic_vector (10 downto 0);  RF1, RF2, EN1, S1, S2
            , ALU3, ALU2, ALU1, ALU0, SN, LnS, Wrd, BHU1, BHU0, EN3, S3, WF1, 
            Ld : out std_logic);
   end component;
   
   signal DRAM_EN_port, DRAM_LnS_port, s_opcode_5_port, s_opcode_4_port, 
      s_opcode_3_port, s_opcode_2_port, s_opcode_1_port, s_opcode_0_port, 
      s_func_10_port, s_func_9_port, s_func_8_port, s_func_7_port, 
      s_func_6_port, s_func_5_port, s_func_4_port, s_func_3_port, s_func_2_port
      , s_func_1_port, s_func_0_port, s_RF1, s_RF2, s_EN1, s_S1, s_S2, s_ALU3, 
      s_ALU2, s_ALU1, s_ALU0, s_SN, s_Wrd, s_BHU1, s_BHU0, s_S3, s_WF1, s_Ld, 
      n_2370, n_2371, n_2372, n_2373, n_2374, n_2375, n_2376, n_2377, n_2378, 
      n_2379, n_2380, n_2381, n_2382, n_2383, n_2384, n_2385, n_2386, n_2387, 
      n_2388, n_2389, n_2390, n_2391, n_2392, n_2393, n_2394 : std_logic;

begin
   DRAM_EN <= DRAM_EN_port;
   DRAM_LnS <= DRAM_LnS_port;
   
   control_unit : hardwired_CU port map( clk => CLK, rst => RST, opcode(5) => 
                           s_opcode_5_port, opcode(4) => s_opcode_4_port, 
                           opcode(3) => s_opcode_3_port, opcode(2) => 
                           s_opcode_2_port, opcode(1) => s_opcode_1_port, 
                           opcode(0) => s_opcode_0_port, func(10) => 
                           s_func_10_port, func(9) => s_func_9_port, func(8) =>
                           s_func_8_port, func(7) => s_func_7_port, func(6) => 
                           s_func_6_port, func(5) => s_func_5_port, func(4) => 
                           s_func_4_port, func(3) => s_func_3_port, func(2) => 
                           s_func_2_port, func(1) => s_func_1_port, func(0) => 
                           s_func_0_port, RF1 => s_RF1, RF2 => s_RF2, EN1 => 
                           s_EN1, S1 => s_S1, S2 => s_S2, ALU3 => s_ALU3, ALU2 
                           => s_ALU2, ALU1 => s_ALU1, ALU0 => s_ALU0, SN => 
                           s_SN, LnS => DRAM_LnS_port, Wrd => s_Wrd, BHU1 => 
                           s_BHU1, BHU0 => s_BHU0, EN3 => DRAM_EN_port, S3 => 
                           s_S3, WF1 => s_WF1, Ld => s_Ld);
   data_path : DataPath_MEM_SIZE128_WORD_size32_NREG32 port map( CLK => CLK, 
                           RST => RST, RF1 => s_RF1, RF2 => s_RF2, EN1 => s_EN1
                           , S1 => s_S1, S2 => s_S2, ALU3 => s_ALU3, ALU2 => 
                           s_ALU2, ALU1 => s_ALU1, ALU0 => s_ALU0, SN => s_SN, 
                           LnS => DRAM_LnS_port, BHU1 => s_BHU1, BHU0 => s_BHU0
                           , Wrd => s_Wrd, EN3 => DRAM_EN_port, S3 => s_S3, WF1
                           => s_WF1, Ld => s_Ld, instr(31) => IRAM_data(31), 
                           instr(30) => IRAM_data(30), instr(29) => 
                           IRAM_data(29), instr(28) => IRAM_data(28), instr(27)
                           => IRAM_data(27), instr(26) => IRAM_data(26), 
                           instr(25) => IRAM_data(25), instr(24) => 
                           IRAM_data(24), instr(23) => IRAM_data(23), instr(22)
                           => IRAM_data(22), instr(21) => IRAM_data(21), 
                           instr(20) => IRAM_data(20), instr(19) => 
                           IRAM_data(19), instr(18) => IRAM_data(18), instr(17)
                           => IRAM_data(17), instr(16) => IRAM_data(16), 
                           instr(15) => IRAM_data(15), instr(14) => 
                           IRAM_data(14), instr(13) => IRAM_data(13), instr(12)
                           => IRAM_data(12), instr(11) => IRAM_data(11), 
                           instr(10) => IRAM_data(10), instr(9) => IRAM_data(9)
                           , instr(8) => IRAM_data(8), instr(7) => IRAM_data(7)
                           , instr(6) => IRAM_data(6), instr(5) => IRAM_data(5)
                           , instr(4) => IRAM_data(4), instr(3) => IRAM_data(3)
                           , instr(2) => IRAM_data(2), instr(1) => IRAM_data(1)
                           , instr(0) => IRAM_data(0), IRAM_addr(31) => n_2370,
                           IRAM_addr(30) => n_2371, IRAM_addr(29) => n_2372, 
                           IRAM_addr(28) => n_2373, IRAM_addr(27) => n_2374, 
                           IRAM_addr(26) => n_2375, IRAM_addr(25) => n_2376, 
                           IRAM_addr(24) => n_2377, IRAM_addr(23) => n_2378, 
                           IRAM_addr(22) => n_2379, IRAM_addr(21) => n_2380, 
                           IRAM_addr(20) => n_2381, IRAM_addr(19) => n_2382, 
                           IRAM_addr(18) => n_2383, IRAM_addr(17) => n_2384, 
                           IRAM_addr(16) => n_2385, IRAM_addr(15) => n_2386, 
                           IRAM_addr(14) => n_2387, IRAM_addr(13) => n_2388, 
                           IRAM_addr(12) => n_2389, IRAM_addr(11) => n_2390, 
                           IRAM_addr(10) => n_2391, IRAM_addr(9) => n_2392, 
                           IRAM_addr(8) => n_2393, IRAM_addr(7) => IRAM_addr(7)
                           , IRAM_addr(6) => IRAM_addr(6), IRAM_addr(5) => 
                           IRAM_addr(5), IRAM_addr(4) => IRAM_addr(4), 
                           IRAM_addr(3) => IRAM_addr(3), IRAM_addr(2) => 
                           IRAM_addr(2), IRAM_addr(1) => IRAM_addr(1), 
                           IRAM_addr(0) => IRAM_addr(0), DRAM_data_out(31) => 
                           from_DRAM_data(31), DRAM_data_out(30) => 
                           from_DRAM_data(30), DRAM_data_out(29) => 
                           from_DRAM_data(29), DRAM_data_out(28) => 
                           from_DRAM_data(28), DRAM_data_out(27) => 
                           from_DRAM_data(27), DRAM_data_out(26) => 
                           from_DRAM_data(26), DRAM_data_out(25) => 
                           from_DRAM_data(25), DRAM_data_out(24) => 
                           from_DRAM_data(24), DRAM_data_out(23) => 
                           from_DRAM_data(23), DRAM_data_out(22) => 
                           from_DRAM_data(22), DRAM_data_out(21) => 
                           from_DRAM_data(21), DRAM_data_out(20) => 
                           from_DRAM_data(20), DRAM_data_out(19) => 
                           from_DRAM_data(19), DRAM_data_out(18) => 
                           from_DRAM_data(18), DRAM_data_out(17) => 
                           from_DRAM_data(17), DRAM_data_out(16) => 
                           from_DRAM_data(16), DRAM_data_out(15) => 
                           from_DRAM_data(15), DRAM_data_out(14) => 
                           from_DRAM_data(14), DRAM_data_out(13) => 
                           from_DRAM_data(13), DRAM_data_out(12) => 
                           from_DRAM_data(12), DRAM_data_out(11) => 
                           from_DRAM_data(11), DRAM_data_out(10) => 
                           from_DRAM_data(10), DRAM_data_out(9) => 
                           from_DRAM_data(9), DRAM_data_out(8) => 
                           from_DRAM_data(8), DRAM_data_out(7) => 
                           from_DRAM_data(7), DRAM_data_out(6) => 
                           from_DRAM_data(6), DRAM_data_out(5) => 
                           from_DRAM_data(5), DRAM_data_out(4) => 
                           from_DRAM_data(4), DRAM_data_out(3) => 
                           from_DRAM_data(3), DRAM_data_out(2) => 
                           from_DRAM_data(2), DRAM_data_out(1) => 
                           from_DRAM_data(1), DRAM_data_out(0) => 
                           from_DRAM_data(0), MMU_out(1) => MMU_out(1), 
                           MMU_out(0) => MMU_out(0), DRAM_addr(8) => 
                           DRAM_addr(8), DRAM_addr(7) => DRAM_addr(7), 
                           DRAM_addr(6) => DRAM_addr(6), DRAM_addr(5) => 
                           DRAM_addr(5), DRAM_addr(4) => DRAM_addr(4), 
                           DRAM_addr(3) => DRAM_addr(3), DRAM_addr(2) => 
                           DRAM_addr(2), DRAM_addr(1) => DRAM_addr(1), 
                           DRAM_addr(0) => DRAM_addr(0), DRAM_data_in(31) => 
                           to_DRAM_data(31), DRAM_data_in(30) => 
                           to_DRAM_data(30), DRAM_data_in(29) => 
                           to_DRAM_data(29), DRAM_data_in(28) => 
                           to_DRAM_data(28), DRAM_data_in(27) => 
                           to_DRAM_data(27), DRAM_data_in(26) => 
                           to_DRAM_data(26), DRAM_data_in(25) => 
                           to_DRAM_data(25), DRAM_data_in(24) => 
                           to_DRAM_data(24), DRAM_data_in(23) => 
                           to_DRAM_data(23), DRAM_data_in(22) => 
                           to_DRAM_data(22), DRAM_data_in(21) => 
                           to_DRAM_data(21), DRAM_data_in(20) => 
                           to_DRAM_data(20), DRAM_data_in(19) => 
                           to_DRAM_data(19), DRAM_data_in(18) => 
                           to_DRAM_data(18), DRAM_data_in(17) => 
                           to_DRAM_data(17), DRAM_data_in(16) => 
                           to_DRAM_data(16), DRAM_data_in(15) => 
                           to_DRAM_data(15), DRAM_data_in(14) => 
                           to_DRAM_data(14), DRAM_data_in(13) => 
                           to_DRAM_data(13), DRAM_data_in(12) => 
                           to_DRAM_data(12), DRAM_data_in(11) => 
                           to_DRAM_data(11), DRAM_data_in(10) => 
                           to_DRAM_data(10), DRAM_data_in(9) => to_DRAM_data(9)
                           , DRAM_data_in(8) => to_DRAM_data(8), 
                           DRAM_data_in(7) => to_DRAM_data(7), DRAM_data_in(6) 
                           => to_DRAM_data(6), DRAM_data_in(5) => 
                           to_DRAM_data(5), DRAM_data_in(4) => to_DRAM_data(4),
                           DRAM_data_in(3) => to_DRAM_data(3), DRAM_data_in(2) 
                           => to_DRAM_data(2), DRAM_data_in(1) => 
                           to_DRAM_data(1), DRAM_data_in(0) => to_DRAM_data(0),
                           opcode(5) => s_opcode_5_port, opcode(4) => 
                           s_opcode_4_port, opcode(3) => s_opcode_3_port, 
                           opcode(2) => s_opcode_2_port, opcode(1) => 
                           s_opcode_1_port, opcode(0) => s_opcode_0_port, 
                           func(10) => s_func_10_port, func(9) => s_func_9_port
                           , func(8) => s_func_8_port, func(7) => s_func_7_port
                           , func(6) => s_func_6_port, func(5) => s_func_5_port
                           , func(4) => s_func_4_port, func(3) => s_func_3_port
                           , func(2) => s_func_2_port, func(1) => s_func_1_port
                           , func(0) => s_func_0_port, OVF => n_2394);

end SYN_Structural;
